

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EErsftIDJVF0m0AzARUB1bTNfa1D65PKFzXVCO3IcVnfdNzarCrieLdbzQivIMAadZGQICQFGhS1
QckM881Qig==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oVVLyVCgNzQviLS1eG+3q0tFr/JK9RCUE5+xAA69a5PzCR+NN1kdZCFY3Hih5lupWCZCqlSR2yxj
T/gFuX/P5PwLJG5+6QmvoI5i4SAxY/rHrl8XM8Kicu6z19CTYp1SPiJ9834l0f0lOlXlTmn836kA
Wgmrcs24F99177fCyOw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kW4owDNqb8AMzEcxlafWfz8koQuLn9mxd/TVVOMuiv8YQ3rvx8K/DGu+WboW7BU9KyEVtBG1MjQH
gJKixZB+7AY25kT/0NwJhM5YyjG4KdEl5DSZuDhsBJip1w/5m+kP4N5/vcsnGSfB2gcc5U+hEZN2
tOLv961hH8596MgBAeOrfvnWa5SH9SROtve5GcJIcP2+J4rtDHR6wFKwG2xp/9kU818nQ53uY3x/
7USyyE73h57I6tiR1+FD47Z14CKQGy+J0+yoYnuxOAdrlqmEtQAPiwIuHmV0R7zwgIucScma6/i1
zxERzOQ0UeBZqrcJuNAcQN3PnQ03sEWGfc4Qwg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iAL6wKTA9iQaAsMi/04OqmErqGG219F3T4DtEhjCOkAVV5xns/q62D9v80Yu9LkL7GOPStNaimH0
0fLZZNbLN9aXY+LXsOjLmXKIRD1NJHFD/6y4EmfJhRxv4wTaSxMi35TYjtTPOpBQ9f3kiGqvET6q
oTK12b3zP6bRyeM2ZbhHWjG88vLFxPuV0/g08KIWxnwsizoJce9xWIbPH46yn/atycdYeI6hNlt4
AsWLZjzzPTaNgwoNSmXe6Z/iHwOsFgDluZ4wunNLVxH5Ru3KpxGf9jGPoEfbj76tqe2kxC3Whmb2
TOD3EfgrtAPEX3iiwhkJ68FGwrBXobVCgJLrLQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AYk0GVXSV/oBWSOxjuGlD2oLlqIfBX5t16vozwXg1+siZJZSMUHEbzptzgNoTGyAuDaMihDY3BLO
EtrWbX/36HzF6OYvwf5POdt/VXMiD/WmbkoqBGEm8hBrg/s//Xc8uwTP0aCjxNObZuBko/Q25mgQ
30NgIumW8FqCkhPd5zaKXjVEqWRkZbVy3s9drUMCg7SmsRWiURkSk2U7gJHgxqNeqEvn/U3HMsD5
przVbreKAnJv/RzsnAueSJ7se+zz3ea7TcdOm8FG4lJPtFHb6jvhIcFQ6qftny2xQ/73EGrSBx8k
emkzKeZp3UgSKQV+dZEMJkjg6+hPhExCSG3ddw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z2aYnMPHx9JY2YhtHwU80KMSOWZwPC6TzLQf1GQQ4Vnr361DuLoPMu0MbOnkBR90QGDH/qF7P5Cr
Ly2yiYO0/eJzmgzCpSyJ27rzee68zFBRRDPmlOAN8FHZvnbWm8t3N4kjdk2vzG0NcvKGeDmWVBg8
WX1YKAu49GjIv50pk7s=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZhLzhPI8pgMrQMSYddC1+njODiKwQHec1wBB4U5W8/l4gRoB3jhisEMfFb5EoL+ePeazVA8YvpBO
fy15vYUdxOsCKx+vVBouvB0iJLQJ7MJ2yB0Atezf8W/dnulTtecMT4xYThtmLmUoLpjc/XY+sv5+
kYuBtkUrJcr6xJNsQtV8JIkAU/9rh0McphkltAYVfKvFQQ4iPL6Vn52nStdWLo/EzZRGxkA2w3hx
RxGGI0fCa662AzFgfo3+9jW4FVA/MfRfrEnMa/qSzvX29NQHmhsMx87TbESpFUhf8rcOf4pNxnvZ
Kz+Rm+SekS5sOFDAnkaGJ2fOU9v6YhYC3w3/eA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
ZiaIorTEQaAfy2fHmnjgXagXExWTMsa2qSIOX4q6xKeTyHrEAfLMwVyAyU6dEnoWQmAvy9n4o8+A
rfFfKIVCPow3aGuspd5Fo6xTxdwqLZjX8zfOVBeb9vgrbGZHE9iKq/MSQcdUYL9I34eqI/Ixle3a
kW5B5C/jfb08ZIj1O83aytZvHnYF2qwC+y7tX3BYrZP6ScXQe7Hyw1oquhiO/rPCUS53gsZeTSRb
Gvv/9eHAhCqtqXj3VnG/o6nQ5maYsHZ99knjsPkrcYalwK9zZNfwZC2+VH8ybpTkOs/fUrBoWzp/
El95XZ4pIC5UkIYA7ajmLuDgZ7HgqYwNFK2BumrNxdpXAb7FPZL7nNrgLMseUz3gOl0woHwXCQj0
XVKviKz+n50hg4+rWOSJr5jUKJoGTzoXA0E2kwUzlbNFb0VwWhATUXMqBPpE6L5lSjcRvhgnTYU0
vzOKlJC/qqsAqi79i8l6AmnCa6FJpVsskCofpi+KifynALL9osNISuawmn0OCuzC4Dldm4nC8aUP
orshik7f3/LAgBVq5/vJCG/HK9LJGZLrVIgmgAVtx/dKIG5kIIVPS8/x1zE6PgWX9W0fm4a3NSJA
FtrCbeh9SH3RRu7DkKP6DCNEZJjkFJK6YQ1ieYi11nSa8tw3Y30dVT1hsuOJjxaJ27n6kgPKI6Mi
pAEfnPblEIyFEvAqez9hkJGVbHVzmPbYdWfujBWYfllgYIEQnkI0p1/coD8DSwbZhK+mVinkWEeC
4MqtfPKd/RP73A0DPXgknOOpJwAzJZgoqz/NCB2hsyL9ijRI+6Ql+3fqM6QyXmtZFqQuF4ovfyc+
izYEd7uJ3lFs9pnwfzcu18ICnkbwhUJ44MRXi/SxFYm9cHRsGT4+TMwiZ1x99IvRu4PbVP4rcgmC
+glEdmMmvr9/dzVFBxZuamGaOL9raB3zWaBUpnLTtcpX/Qr2m9pbnemzv3cNYfCPPfRcxafY6m8c
LJLX5+lChrJselNRN91ZZezBXV5DvuR5y4c8fZLqrILcw+2ox4HKI1utUPEOoM4Z+K6uX1e3nt4e
pHR55+s4hAgmqxTqwo6TVbHfOTk2EpDEOyUbOecBpLTskzDH1CP+I7r7di4S3r3sBOBKUC9cib92
OwzKiudiM3f61uPVVNCwtrBy7/Z+sacagJVmGi9pz6xRT8PtbIBK3erNVxFSrXYTPuHUIlHZVbwd
uKeZK/TIbZac2gkCs4qBq7SXzgSvgfc9NwnZwJwgT3bHPAtnwY/xL84xPrsk2q/UEWKRIMUClIsb
xbJu+cC6OPw3ywMjHAyqDHGKP4z27ctyHfOkBSbmfiTTcrskwpw7ek0kpNPueQUmrtJ+Uznzs0jJ
jn+to2w9Pu+LzX1EKZ+YQjsAW5YLlksnyorI14Kt8kCDuwsqRKQIa4NbRtKNJ6ohVCqsPJFA3pYL
XPx2oDETODPAjmah8i9mtvh25eTJmvJ4aZklchwFYgNWVYEv5rhrkx6fxWiRDMIOkk1iVRdG/BWV
fY6jYuByA5qrqXQUJ26DrWV34JgvI3zbtCBKAm9XkkM0vKkHPbSL3W1CrZOu8jhWaYAm6BdIYqwL
CPOn+RnDrIT0DVt3kog6Panyff2fYWhy2bNIi06tcRtpFP6wtjCFqnHnVBlpDTJpWOuWxMiBNOyF
pi7ZTIuFgS+d3Lkh2dTNZSQiQc/7UAgMZGSV+LAIVR+xt1giCM0vZXNolD1eZ5eLoQlPYe/YDo6L
wmhjkHRn0J0NjVwusUCEUQbGmJqFbWA4aQB3a2BF5hH638gUfqO9lsPA8HBn/v4bItlrrf/AsKcj
A7/nION2x/PnvORxewTlEKZLGJqEmAbOMhN+pcsphkqzC5q4fk782Kesr/VgWtEPeho30GQ9UQyA
WzaKzNl7UW5Uxb62o7A0xD2ebgKhjxamVX30LtkoatNKH+dWljl/fywiiOxF+7NMdr+1n0dYD1Wd
+AOknIOoXtYaE1J9hm+Vq+ErTYFuWIC4ZhXPRLnHHAcVMpLf+Ak351KQlzdVOQKD7Yd/L6Z/wnJ8
NGsdvhMJCOkDfwt8PQn2pFJAjdmCh7HfQVPokE81fq84lJe5JTpku5EVXqSdBznwTRfUqB087DoI
SN4+S3yB1xULXuIeNLLoa9hiuoYccruOONn4V6s8qGFy2coox20drml4HBFkqvzNMI2nWu1G51H7
61d5TfDO05+hV1mID9QpZpNaA4pD7CS5i1sYXqsfibQaZW16ixo2cRhpj8Wx2E275JQHV/uHmggl
OfF7RLpaLSo4y0H+jXSgvrW3o9UaQkGqrFCdCveNcd+bYXtMRG/y5PA7HZOOXbtxM5Lhho+zCaxk
Ioc9Ahr7aU4Cfzy/zUjvd6/8OD82m4iibyJEiZagDd5sdAvRayD/URfhQRmY/WGcFPmKLPqG1jJ5
Fjzt4tA3R+uimdsJi8Fxgli8xWMSKmQmKdlgUWNXTC2eVvkYjjsR9mNZGxiufeKWLWFv7XBlsBf1
U8HFEHfMeUUHCGNn66LlR0o5GwmWeArdNCB67wQGmzYKGnqS4NaV4QntvQYTObf/ry4MGK0kI2ti
ymNr0clULNXyoE5ECeSxNnt6mp/gO+QHsxOZCqTyS5eBs3o8Q4Ocw3a6b4tLUWWp7KmwSorvbn8D
AL2kyUwCO0hRERwOcCMAf3Jwkhq36e69tMWQvvSiLzo3NLHfGnKt0xlxRssIF9wywrE6sX7fzJf+
LvUQ2hcJH9wlYDzPrMW+oDOgzYT1y+M68AA1DmKN/nmkpj9Y+41CS59GNJwog6w6G/WUHOnlKluB
rR1Cq9Y5OjRrNc8ZrY/6T+PsSgQZUm6tKoUGaOq7OX63CMpUGHjmvTYt13prxHi9Kxn/Tqtr7oIy
5YgPe2chH/WZ7tpmkZ+13k8Du/8V0bCdTx8WyeJOWXaSAdNdlSmHAJNCzUnrDMoFP8y7sNz/4KFv
RErZha62OlxnZkow/W1C9mGu8lbhnwvKbIPSRy73tIB9HNhlXcQ5XJO7J8RR5tlaMEg/0/2J7Dsc
SyQ/BTL6456Y1+W63NVvY09F5BYGMhFAyRXKlhLh3LdNVv4iUO0KwiGpufvKyjm0cvsXK5rtO0wv
XAPjypwHl97BLN2fleMryPN0R3m7NtIlTZS6M3FMAjEbxyL6f3QfDrCVkRb0fuPP7ZCc57kbO1xb
qd41ovKUqvhPa5+FmwqMJ0zkXxRhNNNWCOwbfzsV7gGHIAnbe9uwXfw6OuhcfWNOp7NPb3viL4xf
JQXZupBwgthOVa2bzrCR8s63SZbn5i+/XpHHc3esLB7ve7mCMoU2fgSQWB2H+eqHE6vYc+21Sj2S
AP7IzOqtOB0DMMNMLfiaP2tYvVlrnAmTVTRERsAysnFv0OJdiNGC6EnTfsXTrdPhvWBBn37BuBVh
UNTc2Ba7Tkfu4RuDIToltCwndAn4qz3xZUFiZFN0Y7tzOelZcPKwyA+gL6rrVIyJ0j7ojcxpuGcC
Gaq4gACH0VjESafQtAuWkKKSt8lW0srNBY8OjbmP/ujWoSPLee/URTudMujWIoZ6IQ4PblZA88kT
NObu6+KxVkO47tH2U6rYisYs1M9SugiodIPAGcpErb3ZxXGrE++wwMOFpUJ1Pu2TXKrTYNoY8Rx+
vgLT0LIDYm7i5H6WdzPhsT7VEXZWuL1IgbDEbkcNwvxpD6SUswfUeriIfZYZ7VDayQoYEtoeyqyy
e1Iy+jJTcOP1ToWJ8/xzSWXUYZ8MWoa9CZ+JiBtUKdiAWg4ey8577ehNM5d1qw0tKjS2q9wBjPKr
ny05TpZNF79g7taMuu7pUfqH/FCkODpn9LsSPhKx+kF6fIqfgSPxlOnauOZZ5ZVOh0BcBjBh5mXr
vdNouoRonwrpjHQkM8PU20eqxFdE/byLsyVUD+CL3Ble1kGxsE1mAbkANdztQ13WJpj2k8EJrGlo
+f5FGvu5H8uC96NjAdnQRp2yTt47LBSZisH4YGVWCcj/u0AATQVIaqnIlgtZho95bfb2/lwboYdA
2HFZlNf+t5xSTaxiRmb1We3u0byv8XTNYtk09FrkS9iDeggsG1uAarbfp2glCr6LLI5gzj6J7/XE
bwm5VV+6dPG/KRfjUtp2bDIpD31zvoJKR3+s/y7T5+fIfgPM3B/Lg8ZbfN0x+0CS8wW4rRPvcIAy
IFe0stiGEkCaGocZSRxE84+r1+EsWx2rYeFGLO5WNEH6Eq7l2aW7eok1zNawDpZm/CiPJIbuKJbA
vCJyNTflkIopcovNcI3O/U7BW5wXYAKc5lryUFqHZHJUVGcmSXzNqB5VkDHnNLKtpMa8dD4SJFNU
CBbRKYt6PdJkE0o0uXyUYFxd02SVXbYDbQSdo++G1gwB7cX1tYTbuJA3lFzxqmnzjuQQ4vQgqTok
XbnZVR8q83BJuuN+x6hj/uNpsBSKBDoGrZFppjfM86rMvMax1yqUHTXdC+sRbu0RJyd+BfWxTMUF
tAwP1YcbmvxzuavHuqKcBwwtVjQ0bcuwIXNJMBCn1bGkHNDuSeWCujUhLgTzeNnE5z4boseYWfOE
hokxiAuNiRwbrVJQRYyoEhEkDUn0K3LYHuCVDeTIhhuQsSLI8WLs0WRN2Ocpc1vUw37ZYfAJn+b5
z4IBsJUF5bqYKEiMIkakeR8ywRzw9pHexbypM2dlm4ROGK5qFppfXj7RD1b4/dmibgPFq5S3qHZv
xTA79uSAM2Sp9nhCH7ShTtYyBZLtaqmNQ2/GdcZQ/U9B0HnxBOeRHoIvrThEWYLN/O6icSt3ktni
fq7y9ZNtt/pxHIBNx2HYOUJSVJs3F++wwnWlxQUYPkW7DmH3q3bMSa7IiU3QeGxRr9OSClh3ekrk
Nzrpu0CbADwUUi9NDTnv6ob/52BJ2lQwYKNAhfGUV0PEr33WgIweIGOizDtLPeuI5x0XOFW2Z4DY
9m5uxzdJsdI/Ge9lBOVYj4Odmmhxt8uHw2OrPIGONrFRA6sVlw4XTgcdFls0vrMLcwireropESzz
8i1qMWutNAswE4GKTeWycQSeHZjb7FAMUGGqRdMJotIZcsC0iafvon0QHoWNfxfMCGkYGmr0YA3K
eaJHDlrRgof+D+Dlj9Xb/AIzVBFYOYFIDbmTnBIUy5VfQtqGp9TIa4oA02xC6frg5/qKzPC0Q1Qp
onLeGHtkDjJyDlXq6/3DvS/6pHjNMoYupqnk0DuNKsDwA7MpS85mykqQnn5S0ayFPfIZ0QJ2oc/g
b60c9+hRr0s8WllBo0qaYALOQXDVWWaiD3wL4cyQBDdNX0o0wehg9xhHtBnddZ7lv93iDVE3Vij7
jkaDpyWyMuj19JgpAwtwZl2140FkWV2rBDXDg8oYEm0u8G0H4quIIdV3WjAlwq1mYg/buuhSWwzk
ngxyPenrOBHjUvqYOo0AwqJDDCd67GMpL0jgkDb6z6MCSAoFDzWi9EwgUlAY6xtr7D7VVOcwNVOd
rZwwUqwnBSNa8M0+yx7IlVhNPR2O4EITTXg9YZJRklxXdHMuZsSWX7TLluVGHvE48fcX4IeVl1x4
WjFhvhQU78qUrJM8x8v9/Heum/1s8D6/y9GmnQwnvkR1e+vVwYVVfptj7AD3S9TdCavfI1va2OSt
QN/WDH6/Rl5TE5FS1vQIlWgBKODuBZqlVxxuw6JWuW9FysIS1BR+Xd9XiBWlWiWNze2P+Mq5ozNV
gRRUPY9osI7Dpcy2mGMlfSbxfKZ9jBdHQUxyw3Wx7v9PLSHLE7NxIXk5SbXWqdrrGNb0WTQIU1QU
F5AdBL4Z/4uVQQqTPHI1k32Y3AXA5lG8XpRr3TWigTDMs3LqQ/Kt8fBPWaur6/ARFDnU5VeSOh5c
4VrUeI3DgTZrJirwcw1/pLjaWaGCzcbW6RDy3vxoUfsytaoHDLZoW66WT84eMZp8OklwgTQCeyqu
u2EJMddJip+XIMoleppg1P0zEXxdWpWAAszV7wUaw53h7YNbj6Aw8vJnml92Ks8al0lsUG6ayk8e
EzCYdZfvUkII3sN7DeQNreXlzoSwTCULpa04z3UcuY6Pyd0NfXaJYQJlUBCBgn6+McozrAthPEuy
wOyNmOSfBM9uMJQtmJQu4Nz0qPcowWArtuiyod296AR/EMzam0vEFTPUg8eiyGuKlKYSWBOPZmuR
510s4ReMwq5N472kGuzwu64t2mSMTbPajcdKmV5V6iIMz9LMCBkVD298ChiWyW82zGGIclOvXC9J
TDP8mNdosELgJUQ8i6XkBbuduZR/TeZQP3L4V/Nqjf33ZoPQ9E1c4Vrrpy2al0J0+c2+hL+QUELM
sJzphFLZLsUPL55vhb2tYVnz8r94q00RWsWpdgr21gTp4Ihf9QsAeeYrQN6dk1oeaal3S1AqVgVX
a2Djkm/xZrhn8Ot+ksoTWBvz0tNaqL4NQmhJCsvyR7/mUNtItKXpMUJIqxlW5BJco/ZQN3QxbwfP
b8a5EBl6qV/1kG2MTAxinmsrzOhZbooMcsTCxhJ7jzQ+dPksHrqaaYMMLl/9vpHoCYvERYdzo+1O
KutVtMFp7BiQBzeDJvBe9OxzMpZyxSkZ7TIXadqIkZ5JGsiBBdS6ZWZmlLDvGaoZwkp9svCwXmwp
LCxORw746s0omLiC+nlMWC/rAk9vPJ4z6haujshFZ60nDW0asBbUoxR43RhikPrBsASMglBJFN0Y
LXSfc6CPpSgEjBlkZfz721jPgx++uwnXoWZ6Bndiq2RZB2MdQ2HPJFStq2bHtiktKKqcWK9YVGXm
bk2nGgFkTJqq8tFzlXWCE9VTClk6zjenRW9lcbMlG9VN+k+b6vyjaB2FOLhBlk7Qu6jjku4kWxDh
JgN3jSAYuvm00kNqJ+holMvCiNG6srPEm0WiZDWDE6ltr12YoTbv6HVr/mykGnTlssLXv3Bi57z8
Pm92GrSNDczdShoccUXXOvefFalbXzHi9L7bNZR+hcBcc7QHnMMmpV4FTrATcub0p/NPT43dSP+E
rn2zJzcfWoigNjU0fic/sQX/OqDXFv4i8cXRt1rPsZ/98BMmVCmDtFBd6L/ltdwhHaOAzcmbwqm4
jz0YU7IfLd8+JzKM/yGXiI+6Vmtn1BzZbRHYwtU95QEC9MGWSNj9hRxnOftNisy8mwHENz8PzlTr
YKCDxy4OGmFLrxq2m2JY+984XZyltYD0S0UaD1PuqWYi5dwzGF1WQ+2FmcxM0dVkbhP+YnvrkDI6
sqI3sK9MGLi/7XLheoPDBezHo3HY9W+7jJCUS1xDjT0sjzzZD3LErGVOU2vH+tTrnFltbTyIjQBo
uulcdCYL33R9KCXMiAEAUg4qTxeD1oz6yHpvZpQB95tqnToPlm3vEjAaxnGHcLmWbCu6fUkz5WhL
dHZUDk8woEp9OP0rxGCU/2d90q8qDaQUcrXbeaaVhfS3qCPsfa/QcMq4YNHQ758kfCm1TyFIlhul
wB7M7/+YEmUQJGftLc8qzB7mszuGu6XT+fXwetWDk8uiQGY21XP8uT6nn1Mj4cjWMI4fiesuHaZ1
HsEaRFKaAC7ntyNakCcAmP29XlXXRg1mMeNgLBiqZwzjbp16Hu8WYDZZV88t1UT1ZFFSsWaoIL3D
87MfM761e7a8d8w/sBHcVRohyVbeVYor2ueZRqiEtX4tmZKiRmW1/0YW4h+y6FacNw8k2b2VrcXV
JEMD/VZqr4hVtiwwUAXRJxzXbq7s3ZP+gTDKo0IYgNAdU+fJG25Io8OskU6FOz7Bdoo3N6G5aXJC
1sfMjUt7CgORvyp5ZSluiuaVmP0ljtK471c/6R4lmsDHA1j0GrMQOrXeRNgATwY/7KJw2Ns8GqVf
GHvHgXBAN8gD6t3wfzfDkzB5vWOyIm+bphFnDhWdNOGTk5nhQlfbQivWXWQ8Nf1P9jp4ye7X7A9c
04i4xquS5WWT2RVTGzhLrA7BB1oru7cG5fgWqrYJLEX2zpdsWuYOVFb2KO78miQp42tXSOiTjRNA
wza4GwuIjfaQmA/zezrsXQ469y5/XnqwtFCzp0CDetYq1wccCeD+sdvySGbBb5CRbL0oqvf/ccTg
GU8NZnpJ3gVeRN3khKz8OD9NlJ7j5yZhOryYpHdNU7i4lOkKR93p0kinH6NzspwdG/+IMoHAuXMu
TV0gziCBgNdIw5VEtYieyZsNIeBYKKICTR8Oa8sIEkxn/pX9AQ5YGYZNaYeXVXfB8s+4Zhweb0yJ
L9yoR2l9HbnwsikYeMFETFY3nmIWakjuE113v1N+MGiG3QwM3tbF+hBc82bQ7yqhNXWAfSeMiHd1
pc8vcEWijzeqY/btHqsE0pWLcVVe1aCt0pi3WcHv6/0W16ansS65Sb/slxqkw/4n00u/GqoRZ1hk
NAur4PG9sWnNnUmnywgeCSSmteE+6ilImeAIJmgm89rTQY9tGyRrH6FKYo2SC0jpESRNR2L0qtfN
KcRl8KP33ODyGEPjjXu/matC3BFIl7Y6LMzbWaXSuqs7X7UXyIUitHIBOxY5K1FM8AVkKSFJCINE
8f78tS7zwywAcWTFQRQXWk0T/V69Z2OhIwuKn05HLzJ7JXhB+cIlFcKplhzn2kO2q4YgucQv7MMe
rst1AJmBsWxQUa2rotoL4urvlVUf91p3ysOz525ewPpwZDlJWrDgnh7CDfaoWveUBfmATHLdwQ5W
wjXTtEcbPeSJA4YZqJ8dSntIGL+m/ipyoER0PTsU/y/yyUkC0uY6IzteikicjzaAts2YY5m8ARhA
dIgo9aVN+IyC5/c37GikmJmHkZV77T74de9sQNwKHuRJqKWa6iTmvJJ7+TQYdr68ezA2Lmsy1Son
2xJnze2QEru1nE2g2Q64yUMCqG9+slh084OP5fdcMrbH2bIdzq6YeAFKBGS/mnmh/jCxnxdc2PCY
xn6FQd4l6ko7XZAqOsjOP1EUJfrlsCr5qF08bpNrxvXUGyWEgLBQMOxAUhr1m/CViWNkbveQ/00j
ptRrJUcV/tF3D4o5Us5j9mkhTl+iFwyiDGRvw6qV30vwHzJVshcZD8Rp4NZvIDwgQ3DDcP3kk8+H
Db9vU0QmjjaXe7TJNJDMBk4NKdQyHoy3V6ZUuA5zZwC8tKzCA/xeDv/qK0U8Ouk+rSW0znE2fBgg
B1qL5brv7eLEAujVcIRrID7uNzKIFQ3gOte5ILnFgw9WqWNhIHAz1sqfjk7SPVfKFlkieAX6jMQO
V+A8bRg6elcZyIXn6CXM49ewFzOyrytBZ6Cjw9naqvDjYWhI+/F8YJfSkYN0veFyzNqwqHiqiz02
rLO4TcqB0oAZWCNZuuplhx7X54Qp+PYjr/Lmxbe1Kz7Qjax630GfAb8Mx8n+h8n5fPcJ456BA6NU
M++jSym9t4a/f1Sa5YX7Ciaxr4MFLhgxmbqi1AFXJXWfiUGrRF9RCrGbc8x75ZJ9Dg+WV9Rj+CvI
ebvYbn05Aw3WaQuDtceeCxsL79+WO0Wr9g1PajJ/383lmt7ljUIJsSrO7CaZ/o11uRy3+upuP3aO
8AG19xCC/c/lc6YdhtwCJBI4G3GtZ2wl5KaWIJDDX5M0K15eEbmu+CWGwyHcbHmIh912FysB32sq
a7Qu4PDEYkxb8zmEh8a0uwwo+EMYu3Os/A4k59LGAaf9u54zIoQ3iee2+YjlBKsV1ZnW3lUBuPId
1s8cV3/nK+emDq6wjo5YFV2V/8aDuckuSVU0zqirTzDqpiNwaiVNfmXbteDq/eqOW4KLt7xe7BrE
AoTwyhvEYQ1jOck+aHzXx5zT41sTNhqGvUpZekL9RGo5jy96fCmFkQWpgCc95NoCZCZLVvITkcek
HzdhR0UO+K/iZxgeU+6ff65pjb/aH1Q30Pa/ZEzrHQrcLFyQoMfQ1k58PHcrfYrhbBe9t9IVw7//
f6QqT+HG2CS9YCPUjFVGmF+vZLiVJA8B58KzkiUfJqzYmz8caot55swzfCmQrvS2Kbz3e81PCCGe
VdWpvxVEJxlhQQBANh4dHxkFaNeIKxn/cRzFex3ANSt3OOEOinQJmL3L29ahp0rLysSBG+5ELmO8
NkrMNOsIcQozN/+0TCtvSshz/cTN4GIice4SSgai9hsYd4qZmgQFP3zvfV5lxfc2f7mNLDO+C9nP
2Ygpycsn7UFIVISVI0SeRseYwGt5tuXu+5tPdWjDea5aPoGXD/ZVw3tz4OFDRi67PLfwWwjvJ+YI
BvcP+pyg/+Oq+I0tS23bgqMn+V47xVBJVt4chVq8rKJ+ZYR97BJ6VrsihVmRzED+bqjJvjgXFFnb
2Jj4An+8fOeNdqvImVDZGacFt88qPGsedbx0QujwAR50FE25ki5ITb1Zqgts4ppy5ZJsVHrfMXGk
HWr8sUWVl0ciDLOFUCM186S2/x/qTZxl5Bl4Sp6HP4vGxp68t1GB22DG7nq0+8X45oLYNzgFUJT4
P7JRVrNfGdUMIoWQizUSDW/0F3CPtWiVhWZavGHZCt19kWyjMSV2fHlPiT32vtpq8ch8oC6CV0mz
QBiJM/wptb/sZl5UX6MjMYDW2ve7RvVhnENLzEIepewLiqnQqWeKz1y/i+K2Riifm96uCXP5cmEa
1JPbGVItZIBVp6NNny0wL4EeoqH8q4eRputUnZLmkU8qVuzzc/Qhj1AhO5R4Pb7Jzr6vv54C0C/A
kvgFjCRXRcdVGiw+e649ftrSIkTNrIdVoE6R6mr0DmwckwXYVDS2O+OfDfMxQdrkKaBkeuiWF0D/
c31yEk4fyxl96xu24qT3y/c3aFTg74p/+4ZT2zpQiWxdfzsSqpRM0fPX9JnVtYa0dOeFWQC89aC2
oHxXNEJGgcpGDM39Jx6uIIDN1IWVbhrreI4qJOcNxeK7SpCyviLEbPA5uGUxviYr8wxQl77eDZH9
0gOO/ntks6tpm9ZAUVCBM90gdjvvP5LGBazhu9OBe/TjlHgbwH2YU0FCLisDjOmxnajSaX9TzjNF
jM7XUdH+HL7Kqsc9wTrFuTWdh65ERbHpLkluzylSJJ+6d50//r+I670ljLE7TdnltUrRVifodVI3
9O5ws4L5HyB3dKDaVR19qPomCuW8xrM9VzGZ/nmPWqvtFwJprSgVVU6VZS0hGXSeXfAjHuzX2EHz
h+oUlIbqS9ma4H0Iu9eEZjBxdUMLnrlk7SCH9+p7mF5pJVoS7yu7O5h1FKtSkLBYx4AIK6DtWWq1
npifH1Jo3kCHXbOOQgOTdGrnUSrTPrX9gnfwRtgL65R+UGtsVfuaM7lInrF+o+vjMf18Rl1Tbpow
owHCDvBIcZJklXUHW2ymAzL866MMdN8e6TR+bC5dr0CdYBR8+oKGgWObjePxNwOz0Kob/PNV5sNT
nhDgxGnjO8OxJCRk4pgaQp4GaozoYUGSRXohCYXho1jE43HM3jxhxrC8yZkBGNo1XvsCs0cVHWSt
OC71AobVAtOMvXQVGQCkr/UZFCoFMww/mGv4GZLg/UZ5IxKwsiwofbju//tfsdtHPZfzbSTFBr/4
Ke7K1xmGxV1dcm5tV9k85wUdqtjN51aiLZNPNma65ZwYtNSAIAxSPGv5SU4cSSXORemus9nyTj8R
hJwr1dNhTUnSE0jI6faJFD/+HKLrEzEcL9aDvhdVTXGalbLdspO3Sw7kWz1KLfnY3jFPbkNX70sy
1raAdrNFFNqMoxxEyhJ6fTBgy1dczpNngWmiRC5/d0iV02XoHnXVGOf2gF41bvDzkvSSwV1kj07H
RGAuzbI31p3uExnQGkoo1q1RgfTnjo6B+o37/OyuJ3k6faJIVFGICbt1nl9VCLTkM4w7b2l2RXB8
5BM49DLhZiUu6l5wYNnHivMKzMkpmT2l9BWclOtdr/dXEAW73W7aQCGxnGGxjnunbb94Dj12MUz+
k5lSm93XeP4fVEeUnr0sniht7xAig1XxLmR9fLfzsiT80QIYeoGgmD1oiETto2AEd/7F7SRMSDjc
rdvc63YYgeCve8A2StY91LmF39vGLEKc1bdGGsoIiPUGdahKwf9H032rl+VSzB688x+UmC4fajM4
/FQoDroONyA+r05OpdXfD0ajerMGeVxe9/eoHC/QtP2/9YspXjCTOR5WGEuSPF1fhqZm7c17Zu8L
r/4O2kkPTSal2aahMXHFNKyD8uigcbXrs364GT82H1kPLaTNNTGfynlCIfWqVnAC8c9jTau7Idzl
0WOWl3c/cq3hKcwV8ciDok2NqFhzcjEgmpdDKTnEubxD5RKy323ZAC1lJ5t0UZhjbsWilYo2sN90
DYIwP/rZ4Aeemyj7u3vh2ghfR/+/a11S8zGRiVLQI2FVlwHiX8AReKfjI/6Puw4eIeAt/zmYM1Dx
UHWC7Y5XOd6NcfBzF86uWxwp91N/DzfRMU1Qh3uhwbSaqshjO3qfF5b3EQ6J1rK72wjxTNhCbMZH
UiyFoqAD48zh8G0cMpCcJ/CDlMxpfSwReFg4VhKI24rwkcrnG3NwZLnmqwSoFTJ0k58qiFABKzBS
q/PAHuIGU5Wjv6J0oiaUXEhsegouEaI3XAg6pJAPUXISHv2ES1CrbzmfoJ+hnHfPCJvJsDjmDo0H
2W55WYJ8Aq+7IjbtxNS4rE2BmFokEEt7LOfsYgI4TkvwblrSQgRvcKbBBIshIttfC2yGxXCq6LnW
+Em7D6i9VwfrXqmV/X09VTCphvSGIwZVfSYGWa5sOPCNI3nhM6SPR2+kTJdspQD9v8FBap34Gtp9
qUl5Rxp9XhV55UrDMOVrqJzQO+EYzPwcHUHjqroSfBN217sYD2GrNQVzJ8NCI2Z9eeUnUodtGjoM
3BH6RTACrbr7AaC+g0YiZOat51QYkeRiQPvBc8eGBREmYwRuHwnWM1nWY4qvoVU6oRNGZjSOPRBV
Y5s5xK370BDchCjt/T7gpiYrq89Jb7hlOgU3hfww7fXFCgfDJJ6ZpUGoZ0BCz/PmE41e2HQ/bz5t
4L/vdpW83iFcz9BaJMpiIk+57xyjBPXedNx+MTO0xUqKhRt9GpkvkQdkcSVtbFyPgdsFDHfhFI7b
XMTBhDHU7ecoDwYfjrmj8I3WP0orv5mNXMNaHlmL+XR2L4BmZnlaHqi11FVPDdo8H+oHdTqDhW+B
pmx7J7C9PwQkQqsMwrValENJ9Ft//82qinNITOXTsNxQ7LDB2CmyQchuZgTWs4JubWQaRdqKGa48
TblR2BxNdiElxVVi7H7D+lXHPGpzZ/FajMdHeNTk2d/cyGInwK7Vcthk94DgPzdtsXy4FaYCsvxl
1S3jZijpFQ6sRyrxim9mc0laoKlYJ+xwHLBg5eSk9xA3eAb+nwUpcrAn4f5VWL17ptE59WO+LvO+
o48HfXSC9D+N5rUYjWPhuEgG5RxUyDuUkrh/776UwcP06SGgHBuWAyQiaXOKlUQCaCeG8Np2WGNp
VMEO72eB3Irkf/p8XO9L2OgJh6qeMmZ4c44Qu+EhprfO9hBQtaBLAECIFzJCK1nL9Sm4Ofq3ERAA
k8hvlcdIz0jqPC8xQiOoqBz5NOFrjDLuP0twE4xD6JGV1Qe+Psls6+n6MbJBuwlsWLlstgdaxlkH
zB386kxZc1AUT6jSx6kR7NBy7jtQZiQ9jtafVP+w2zxDXwQf/0vLqv1XY2qWr8G5jpPre2kzBHHA
qSHoh6D2tvckNCgPEVCP/oekVfsc722PJDh7uDuD6t9E9v1I26kBMRCetIb1ux3I6st588etIDxy
e6lx4Ki11wzUSV9sdyZwgZEchIFZNDjoojVSUB31GtEtxXOT2/dVhyfVfiC8QzDu+bOpzUTHOoM/
LDP2qGnwaCRrG6dcDqjaN7bAOUR9tuhYnPIb1oAmplecCAqN6vuhU1X1P4oVG/QoqQXoIipcKfWE
Mza4FzPJhTVPIeNOQFlu25qg5vgG7Bl6JjkDBq0FIyTF+qDAYb2xaLgRNUGzsO7xWA/N8wV39vDq
wvpx44ymIJHc+IVswaM+t8MLJxOV6AolkhgM5betG9IDLf8ZB7JEvhQ2WBto06HH+7+XwKdXJVxE
DbE6UH+VH0Md5zhY0iUBflhG6fPxIf2WCZBOKY+NrlqbzH452UsOtw7Va0hMCd8Q7vwSfZYRFbgc
SE4Duz6tH17g+V6OAMX5eKZHE3DAu/wF8C1eaTPLskVESlUFaf3ZvYSjEqG8Kyf3NroiQ4qasfgc
5zLZJoF4F6R8gTctcCJgk2Bcr9ClZ8uSRKG1U8oIICLOeT5Psawl6IlnZyvsYiM5kzm9hwZwtbCd
L61480RFOG4AJzuqsad+OAP5ALf4nMgrhCIGN/93GLMJIhwtwes5biXkQ4e7MCIU9U6Z2tke9+LT
25g4CezAp7kJxrcRJBMohNakkfTA4WvYvn+P2WmDMa+jNAUOq5Fzn07tqqbK3sCkbf7gg62WmvoI
l+ERL8JucaAO0jtXRYWaxBnP1YxRhb9we8Z3cDvVrJVIXC3c4iu6wp/tH59/JAKfHU2VmRwEOpi8
yXjv5VwdtzfWx/m9cvCk5bdUm1d/3vK7qITqBvuxYwg6HeGBWcHeXwLXoxbpzuKVuU+VVlE+Mhxt
3AlRlffQSl7f/1KpPBCEkasR+ygjif3GiosMojXuL0pL2vrSrR2w2jnkoeD4QXgUcE+A2r/xNx3T
j1o3xS4c92sGFb8T8JBeN49gCFcuK4Xw4RFPOlkwpSf0jvxlLKfLsIdgscIX5yqf85hiXTv5S5Ce
lYGbNPBtOsST4sgaxhI/eezO3aU/Uvx8ECWGqLSSxea/3Ap0yVCgQEYzaMVbhblZUJEC+ElVtuil
NCT832L2NEupi4dVYB4qnmQKdYuLNMiJ/WCGurN3rmcqRyaGDXObV1A4RhkxYSC93CET0sXon2Ne
DKyqGeIBHWhlGDvuMDmcMaS+5dc3pN6pKFif/IDr4D5eU6UMdiNQ1m8HzRZ9Pg+3gm/Rbly5euIi
+dbYCYhgcFghLv/9wDn3ElSGjK5tY5oL9ZJBIrjgtm21uL1gbNSzcS3GeUaSSZwuOS0CeeId9IiY
dV2RYoMrdIxYbZxX+ZotgZDTBijQpGNvgMdorGXWd/fN2Cl7HuP9djKm24EleJFn5ompqtXnZ7H+
EF91BsaXIbRTsUFJ/yaMDVELnS7XSqsX6bCsTvr+Gjjc3fxqkzbIc1GvAn/44LT/1mM86hLEJjZB
4D4xaujFzky3tuyq0VuDHqyj36fzH/js5VZ2FEc7aVeErVEwebbHirYiZNwoC/bsAkH585zZdTb3
URaShwBI0IFCZ3woQenR5uMjZ7vUZNzby0zbmCZTwaszxKpzwTV6Vm4rKqOxwoiu6ZKvF09LkVp8
I0O4MzCtpJ4B/pvTl/GvBlDK5UW2bleeXePNIPWDGR/DRV2QSvDHw3MSkPEKbcatakFhGIqQSCdq
OYA7XgBEKtvDQYMxl57KipP0BNETNvm0yQmf9XJKYkPvEkSYuBPRgLoAf/VGwA5d1Hjg91YYiYsI
R4wS57xhm4yvUtUfrSYUC7a4cEYcHZQF5IDg/ble8zz2Xpda6d2Nvyaom/KRhbLBejKbe5uhsTHb
ktrrhAxyQ0zOd193CFRA6988SYQwwNlQHI1T6kzNh+ICvQhiBTtB1ZVyXlEi7INuXde9l2mU5Ob3
mxWo4CVloHbZHFlE6Jxi5PEvFaNRysoP5ZZUspXBo8nqev90LzMGpq2BhLzYIAY+1jCcjmpzl9SB
2z6RG8MCGYrsM9x3Bnfgu/zi1BlUnnIe6aLLTkD2FQc5TIWpxn4tv3w9rEcUkAE3Kk80ZemMI4lP
pVFaXvni+l1H/5GvsVu0NgSZgeScUK8fOv74fTtu/k/YC/48qJestjHz5P28g40AY5PgG3GEn+4U
GdaSp3Ina2EqUqWFMFi7Q1q/qs6GndCwfNC7fdihD99V+U577HjA3FGCqP2JO/9RHefOX7uL2s5g
plLG0vxvafZlaeqbrt38NdWK+1A5r333YKr4+sVONQAzF1Jb72YCr5LpltK0ZjwYgS7sxZGPnqZ3
Por/N6wOnxYl2JBv8KGKBu/MS3P8ItfU7GO0pOHgGQFmaPX2SdiGEtNKeXwgpRHsB6KrbWVJiDWb
O7/Lhi/1RN01xl2Lh5KnqWTj1yRb4zjInG6TabsQad5kJ4HnB2prCJC+9al10pCrGf+nxndUb6oo
i3ZQoh7GKG0aWrPhyujt+3j2gOsa9cvbHlqAhKao/+z5xAB8SdXjpipVQYiAPRko5uEHD6vE8ZSh
yzTvsqaffbyA3WXSjaRDzKk/TE/kFydvhbiLAh0/4Qd9ucCMNVm6RXcE59efYZxsDpGkPhmu0nPC
xj9FqHDx+sYRjBPCgTJTnw0wXI+ZC2LBxDPBxZu2tEtu8+CMUmClaXq/LW9GbZKaAxRbrKLo9gLp
uStu54Wqa+x45QPmw5dgfq7TACPwgEKY9gkOf4vqYPwSSjrscZ6xXmZXhxrylt65l1Lz5rFKdMt8
iFEnbNLKecfUe/yp11NBRY24cwGAomJg0XmOEpnFW+O7ZpLi4KDrBOLt41W8ndXWyKjX6P4BPVUG
aqnivymZq2Dxy+TNjbmMvxbCf3uA5QB9rdJEYu88UwP+ez+cot7x4if77qiWEcz4m8yxgoQaOptj
LYtiFJ578hEwsTyJVyaYtJF/Ccbn2aIFvqbXFebrKmNzvQaC5ADHKbAG8MEnVBxHU+CamdTvdlR2
ngYOR5d24TGMLZuIPrkri+K7HIdXlXYjveYGx1ok+ln8b/smINiDa3pLvzq6Ueq9FDaLVPRmhrDi
HPFTmMl+8yzP4o7sxA6NaE9G47O6vIsSw7bk01d7h2SBIql4aVphL41ILURIFChaYndibCQHiuJ4
pKBiFpAUnhk2qE52+eICQS/eIyMCapoq7tHJVoKFXH/eRgHQhm6mKno2kGFLUuvPi86Cw71CSORJ
eaYxtEucz/ZQL0mUY9x70Cg5FRP8fAoNXoyMb3KQOPzEh0XRInfqKD68LYbMWT0tjeTjsxAY/j1k
uix0hy5J3RKurJDPhj3ZNA8wibCQ0QKX4naeaw3vRNOiL7jH4n47tQh4xtzaFoPhvEz1MKrCWMHj
IdnNht4tMh8lvLOT1o4/O+JtsyBhTb07WaySWWwavLAjWkDp48MHQf3fjhhv295jOjwo81y/CgHr
p4LDQxUcBcQaLwkdbFnwP7SnjQbC05dN8cb6RCrXcjtMbfZMnTnaA4bImK2L6d5q0YKXsaYXQwub
2X8Uz4UlPwLU4ydy2HOh7YQBekCD7ZMnA8Wk3z+XeYy6Pvn2cmLAJyLomBxENvSSZOA8h95HiwXA
YDtQtimOrJfOu0tDUak79j6z9P1bAFA/dY9+8V0K1BkrzvCnHHWzTcTKjjwiQerhwikwQQAnN7Jc
5U4+KYv/ea3fxHPVY/jrboLFY66RXgXLgPYeuc0dgYbR2VSMaLOQQK7jJWu+DVmPSwJID8f0/68G
LPmdMWOd6QPam+JemBdwKDd40IspNMTfLFgB2PJznSUdY671E9Re2mDI5u+hpjufHsH/gaee0DtN
hlsi5Ifv7vTtiQj2lOq+C3VD08Vg5F2hPFJzMPHBKxex4VHwjKu7DPf6A0AgW2UveumbbvUUfzhO
NWGKdP5l1MYuf0OrJdPMKgtU5VS/LzV/TgjwbmboV2j7SYpCQDBlslaLo6tiwt0efq3crjPZsi1b
oGbnOrwRcjOMKQj0Oi/07uOX7tg+kACuTC+a4brppah8bClB+uvXoL+cdmybcSucfxNncT8nHkth
ERov7b/jctTQ2NEDvBWpJvLovDDpE/eB+PA6E3/NRye/T4eD8sPXkPteR2oc/RuyUDNXSLWv1xGH
z3XtqtDjrGDonOQrJzZNRzAn9F+v3a701xsaAkIU/IJ1B7MrFeTWAMlIdpFDoGjSqYdtxquBOGsA
VLXs389C6bQW+f/HIC22M9GcluPpBxPBJAzJMpaasTkHMMzzdR5xuup+NUDsfMzggexQ2poluQtD
OnfW0zPrwiGnXSAT4mXFM3tdO2Epg5SDMYNr6Q5ndHDEm505qyILzLUfbnDEi9jRUwC9uQmhkUTg
nnJlblsPL587PR3Q9+N23RIJmCvCZ046xxpwZiKw74Orcvn5022OTVdK1beB42LrZwX4WwLpppac
VbrJdHVGqDcbG8r9bEYhhfzmIvDQwBZ46f2zO1W5onUJpaF3tA+HXNons9MDxR+v7tAGaWYs/xXa
fg5H9opuq3YgGdqKlzNMKZyhTQK2ng6Pn7xzlfE8zpIaDhk62maEu7a0Eb8f6yUJglB3UPWstuLF
55LNjMQaVIt8+Cy5kTofv/CPLbyMNajCS87BXC+UvKxrLtKyTr1xel8xWEQcwRbeGOPHBdPeLh62
C+c4M7bl4J0Ag/SqBHgXlwQA0mZ8EvdGjg44fbWxmxOdBjDwmG0niOTutg+y7gEJjztFiGukHTmf
/OqSvQkBvL7spMHqI/LCfzCdPy8wt7tIK8qTeQbO2STrMNzI43ftzJhfQMwLKU/LXlpqvauC+GEH
l8OdKe0bYyVG8DTAeAJKiH8fzQ/UkE4NsAmuqyRTmuqpmdqgoJSp1w5TKPut+IFGhaIyCxIoIXS0
IBmllCJ0+vvyaTJGZx8mBYRsUsppzIYFiiCllv+CRi4JSolBNVaHXAdQbkafqkD6pVmpd3eGzLRJ
yG31XtmRL0AiKoCDswXmfbdaGT4p7/QWkrQzxLrjK6+JywtXziyPl1/4PFx6X/hr08NwnJ+pWPdR
3FHOnpqe4w7u5FgFNCzavGY7aBRTmUBm/i8TtAT/hGudX5nP57ZHxQSG5yJ774WVL1prrrEJlch8
pX3iKj7hBpyfEKSHuI/tZVkQMsfVyBgrMT/Udib7QBhyAyKyjMJme6cVXaWDbEqZ6BhAipvNF31/
9NNcvLcpROxFSG0lx+VqtlwPaC+SR6vmlY9t6YNMIzUUlhdU3+ffGhM+jt7QQDpehaEZV0r0iEYw
ONwIIq0L1m6919/tJlykO3AjfvWfRq3CcxjeNgqA7F6zj92ysIcjXxGJCyspuNqMCBLdDt0rNaYQ
/3rDop/+TWHquN7YMpTy/HC5Fnoz9UIZWSXBDl0A0kpPNHA9T70wnRg5BTRYjpgi2zpMN3QinQzR
7G4Cx80mx2HreNN49IBYQFZdn8eQehF3f/DFS50R+QWDJJZs9vy26ZjOA51BgHAB6GrVRNfMkbud
YfUoED45lMRdEPEIGUf1w2Uo5jnbYGq3+yQa9c1qX65oD3e3W8u+URQavS03s4jzBhjv4+td9giR
uzda/j887FjoavjQkrLWYwX8SVhWiAj+lM1+DAg+Z712gK31j7JA6SjYhrzmBVnqGH4A9EIN6U+I
A1kwdK/HQDbFQzinrIPUJRanKi6Dz4mDPvviZL252oUUrA4r5jZBkxCkemHk5O0DvHU5yRs4IZAn
/cbhxzsapCCyw4FqgG/VkkbL7TnWBmGhdvqMw2yd5v+LM+EdFIG9dxkKL6GfJoAu3v4rCWoK55SD
OrQf//iQQnGrVz+5glbHkJ/76dAwAOil8KJ7/r4TMF/df11OOgNk0x+TIKryzb1jW9yfykxw+IV9
fK0cnEFJiJ+F52icttiXXU1ayuT/JqPzhtxl5RcVJQUvI33I6Jf+F0EdIpL+x2chlBMsmfFqih9q
4ofHTBl9n3a4d+/NLIr/zpe239ElFldxtGt+9EwYGZnmwAU2EZbm7FzT64Sgz2qj5j3tsHKrzu05
HOYMVSrDV7KmnIiHIXdX2Z8DhaULtDdIgH2D4dkHUKhRIW86JCWZibVhUn+Wv9NJoNb9dDV289b1
X8Pcg8geWL2vcBYGdhjxJI40xcZ70f1nSe02NpGWS/RCHmunT2SoRlcdMoQ0Wd/Sm1SB8eoqSRnG
fcpK4XmN1FUn/xqBl19J1TsTJOIETIdIEjt3qdC+bN7XtbjnvfcbfSBUBo5NT9cyNNalInajQpyi
aaZwP5QwgLPVPPsU1iTBUQatsyHlSu/3jIJMvF7223e5oT6XxScq3sLmHLjtemRwRvANW6FfK7Sy
S9LhTFclz9BqdXQAjYs6YM6YyGr953ro/+VKk90/m3EXjfGMJlTUppyfL/j7ZksMyHNbWLmbVjNY
ktgzNHDGwsLvdQtoomn05kmLCHASnLlKljSAmJiIi3rsDclAvSauMsZI1Ck4ZmBYpQ6H768fbPSb
YOkuoAsvvk4ZqPYtrcOMgi3KTkbGJWCkOxSXQqX0OH7yK+XKiGa5399qyaMu7P1eKZejnbvslF3a
wUCXNHSM6ImPFV5qUkfAZkbUKA5hvxTW3nazWLpQEqlvI0m8JFlkhOJX5n8DH9oHCXIhdHp7A2ha
ZFADBodDTz4hE0JMpP7x3s0yf5JROPPEJ9mYHxrjqEw2u7CelGWaZCTFigDeGal+1VKYGriI85Tx
blxiAWKqNhj1E0uN5YPB6YlBsj8JLmIXzGMc53jrTy9byN1K0d33ts9IThnEgpDw6ykxIeRJcZPn
IEZrosPbqZCtnkxK7ZpIrBPhYtuIWvhkHI0G1VyMspmKWvLu3lXnTUxowPNfGDdAtUmIIUF9WOk1
TjHMjU6HOyNHQmvCLAkxdnqKfI9+MouLQmMWgslCLObomwFU2liK3dCnhdlgrnoz5wLogi5rbJBg
MikA9WkJsJ4fX3trqiDvyU9gTIVJfahYVHhfmNe/ZJy6vee9BJ1EtKRkw0sb9k85WaRyv8nlmGmG
Fe8b72J0Pxv4ElNy1VWpidNzEzzz1b4rFPO+r1Tyk32YJ9VIayCDfZiquA6/utYXzoxzUzSdH9Kf
4D4fnD2Om9kSUvVaxU+xU17mAVfjl6BUp16tqvajU5UtLmYW1M2OfpQe/1vYW6pHivzQx9Mv+qok
vgdSkKxuEQAsU76vb6Tmp2Zah6gzy3/ObNsHf1aQu8eU2B7+5goYH3k6M9FBXP/AQ4iHnf36X2m8
DbSbEuzNJoKsZxXpeFAQLw72TG5WUsbV7LJboH9+ORPlcSfPkCT26ozMKVJFUvqUGwLYJr9w/kBU
unwIZAmLThicqrUF2J+FrD1P2zR+pY0194WNYqoH08bQ2HKe/u29PnU0E9oXHIbvDf8jROiALKu/
G2ksinrly/jTvf/fGJx0srTI8BRjaYgXaRICHPDQhf92XRsdibKGReL3eqW6W8KlCN500vXOCzR6
amv1W7YBxyD8dXu+D3pHNBcW/dra2Lh4IUxvAPytTeA86wBdbO1Q3K1wsS+EOvKW15ZtTjwWFNFq
RYrD+e0OKHqqVQU+ejILHjDQWrzSn4egH6hCVjedqVWLshVLVF7eXdEiU+s0oLriCCx/4sCLelN/
bLbdYEH4cX8JOyUwyeqiGrtLLM2eHrg26EZfOjgg8wOsZCy154CfLtqUp7d1vT586vhZuRahvQ4w
EF3EB2Yesegh8qUqkkCf/3cmDPJUtPOWPX1upJpOeexQra0m0tMZ2eGIkfwHrJ5X/Nt541tcAo7a
rON2/iU3ue+gC4+kegIim7U8tTHm1TLgJmxD7Y0sW+pu0gwd8SrZUN9eBJmpPRObP7fc7xb1B7qy
fE1qahq5ULnjAsKW5ML4hVcH5SZa/XT11pINdYft5UrNTpRlJInmK81o20jZsKaG0CkGTtN1uqCz
r5/Letv40PInv7JIvA5hh+WvujiTX8SWrrc6E7mmAw5fkV3elumG/HCzSMMiqRt02bbFUB0wF0Nx
BQst/dfbtdbquReRK+rE28orqIcY4y/tRpHeAlm6TgspJ7En8sUbKLF2+gukU//0vh4Q4hckbqED
WamhSj2InLNa8mgT+MR2lawDIiBSGLJPuIAUllGkV0KVxsEXy+FV8j+AZ81//xZfnGxW76MXPHuz
TvnwZnAZll8Z5JdpcIOF4xknuUyf57FRSWmXyxgOeRbTO7Ob815vwFYueXmGvq6eWs3N7iKfVqVS
SgDvOWC+ZxlBu0qdbYvSU+JYVcPrphydfUm9VzAO7bEDoSI8kzzMxNVfvtKEllLkygYO2C/5XEuZ
wa5T0WRdEAqs2T14JojuX+29H4bRzDU2oU2K+ADsQusMfflPFWBZBPimp792uqQINH6GsIYKmL8y
wxHM5vsoLyCNUDn4MncmRXQm+iT1JcJUg4iyRQJkg7OIV9aMu5IU7HLgKrxrPE9Owcn40CqAdg29
EzHWMsUsXQ4vGHAyb0dWCE3sJnUUwMyiMSTA6U4FPWxHlZPvpK9OoeDyLYpm8L9Je3Ft8XFDi67i
FkK0XA2353KBZy4pXFCqDUZBdYhErdsTdnoqt9sM6akBznGbKOKFT+uSHYeS/cF2bDCknCQiFmgf
h31P6F711lwknkN4Ub7oKXDY5+kATZacwWKXL+vtyeKl23LXi2a7cNh+KFTZrIxBRJQ8E6+ByAED
+dbhMpD5WS/jPw3/qWaDABUl1kgl5ncq0AUBbgSiLnK0WKaia81NnpMN2Jul5vIptwD49GrNz+qD
XEsyh/KmfidfLZShU2twvML4TaZy3LTj2xtsO29nmD1AKIK2W8qzN6DR+UFqCNUdegIaJiSOvmSW
Xms/6T8jW3H7Rr3GdmyowT+dJEBaoQWpSM2JqRSSA8AEFODsxFBCPLqvO0dxEZ4kGvGHE/qrybYG
aJ/8s7KAlg1NlOZZc0E9nvohKpDAolV1Zqqc7iaWhz/JyMvBI+2PqG6SwUc1MNZI5Ruim3KIrizD
JWHOMdhxPmdIhjR9YIHfjTFBvPaSktwa9c3K7m0xFt7rJOxsyR2c1+kz8m4OGbwAevp5Fx0kqkk3
Q0rE7ue1bJU3HtnOS541Ocdr2+GW1ykqxNY4KeCrfC9qvHfejXNhocny+D/YnG1c2GB/2VA3PG8n
AZWTmy9w3PGUAcunLscBIxTWYPHAG1G068g767ArAYeB5Vx+jHLhcAF0UF0FzXzM1S35ub4b1dzQ
40HpCsUYVKbd08gcawWSvBr1BaUTtrY2qD1BsLxFgJSlnlkGQlN78abnZ2CmuB9sy0amMh9ijKH4
SspkoV2ObufrM3mbVlDOy9QZibUy6ii44bmqYGUg8baiD3IlO5GYPQWEfMOMC/jmDo5KZvelrxRu
/Uh2tJhp0rQcYOhlfhWOonrMWpHOGwq7XJHjFw9FXij+VrG7RZadGOiYBtJXFVbYM57vmpM0Ou2Y
AulipgQbYcQ1NdN5lOEV9yfXvGo1EDhnvqn45x/5zAWLBbx0o9eJLCTXeJL3PY/D4nn8YOq/psJ5
Dy6lmZio4xk9Sg+J/I09oxOeyY9e/ZLwAeLMPA7wYyDg9mYEJiaUtvRQSkzfqCcAdvJR/0mXeQnx
bikQ0G0eS2cYpfV8KUzf+1AU8dLxyEG5E11hGLACD+zWaka6qv1yO2MvU2Dk0Wbfxs7u5S8Pp+pq
jM2vS9EXKRWnt1jOYByDkL1fSIczmkjmeE0uKUPxxyQhDqOig9wHKTdNHi567J8+wbdWByKpPZYb
CMhET801lmi0ljDeV+XJiwXZ8+/LlgkJ3zE3LF96WUi3i0pDj0ebt55vcmW1Hq7+HffU68D475eZ
V1OrBL2dvp1xH+QxExk+pWwQ6KE5pKZUr+L48pXNn2Eb9HsjLJW+YafhHgE8q012T8Lpo0mjVa6w
JYALL/lgxRjHlLREnlOa4mndSApnU1rJIJrq9nzFQ92A8S5cEBF7dN58Ug2hsDGCJY8ICgJUFcew
wOJhWHX/a3vCwOzEK8zgS0yVDt5qAxeZvygDKkHBS9TTAs2mwD1NRk/c0o5YZZHnlAUSvuNj2tU4
w6prFaI0gx+t3xOPC6zj/FmpjIy4sp+BNaGhFCj3jBkeJiYVBGoloWGRh6BGsM9oO0c6p5Y0Brx+
xRiIJFco62ntQGZrxxDHT0U6jlkQULSGVLv6AYhL93/FFIFuh7vmdVUt4RLr7YMegaYdabp6r+o8
WVdimT+Joecl+0IL1rORFfw1XfWe9Kazjx/0Awz7I8FSiNMuaasW8XhtmeZ1c4y4NrOi5mFoBXZO
NRqTFcbZKN31iUVBBwAaYQl94fARrts7ItQE0I4/44LdVgo/M0UvyivayxJYPKqNshjF+ISNFmNN
nYLK0a5VqVaqH4uQLcxDsVa2Hm0wvXqFC7y4J7D1akv8AGOAJ1yEmbDbBg1oVf112DN5jvzhJuys
GODck/k3OKua22XnsqQGBX1Ngstk99zTR2AEfrnoJRvov/tf0I4V6iOK0Ry77PMI7hh2tN0XKuD6
0Sok8ZGjkrn8wOCBkMrnxq8eRBYToP9BbjoJxiPyIBMjReoKSXKWCL5Prls+cFyUj8Tw5bHZDiZy
NWUM7kI3aMX3Orcf8wD7lrDt55trrEeQAkydsMZYybTsKI3J5w51JTqk6caz/ez4P/lIYPgoptXG
TNGn15sNkXeqdjlE/eVBEW+S00nOcT9YfeHyUCyDv6Sa3xyCRPXvnuoNaXbJy+jY7ygMYc5QoLyD
cGl6i4fTt8NGZBqarBV9HTp1K/Tsyeyy6q1PBOdzp8ljcBZto/y9bHqL2M9mXxb0sdR8qCczEbeW
wP/J5OLX/3vTKMYUCuF4k299lHBiuvHQM9qJteR3bDpb0bf6O+cmN6075xaia/d4ud0PTmE2dzXL
wCDgmt7FbvoGniWHYKDFB5vmKR63DWCkPLWQwUuRfDBHW6HV5bojGLTW5romplIRfBEueCSAU0rw
PHCanmcfzfX4X3a5izeKJPUwlUqldOCXzzZH03uSPGQK2VKecnD7D/xux2sB2e/SnznVeHddh3J1
Br6zNqAbL2IjMVpqBbZigBOBjUIGpB0VqtQ/oWH+XhZDXWQ6zlJk6uMlI3SE50gui9v+blaP2Y7f
W8DkTQ5OLckUd/VA8k8euDt2H8TuHmeXLYuiZYmYtX4TEFNDOzSCDIfjG1GI93O6+EwTlZv8+PGn
wwELf/jKFMoCE9mSLyy1OR85tJaxcWcMY1w737bC+SJhZ6pzkVtWgV3NMPTCH2C6aHDRS9t8p9bY
qoVlPwFkms/70SmIGTT97cmK8fKCW0Z9cF3kXEs9csSyPepw1nkP/X8K1LJFdOjowXJV1dzIwnn1
wwyRV0aPvvpZP00J5iLsZcCVby3O9q0ptxlMc+PJTfoNvqaIClaN1Ta3Ww6888mO5LZSTq7cehO8
8j1BEYvC3q0V8WEmoRc2qdFeUML0tHbqS5JPONIx3RB66ur3sDUFRNP8I5DOZwFnabUOJ+iHJMaa
WVyeYODSZMInr4GzcueAgp8+xFLiWPmyHmJ0286aVOCgP5hO/2RqFws0ABW1i0civalUJ64WBXr8
R0fEpL9LSgGyLpSV9rhf0MdPmqdIpN9uLb+pTNMOb/JMWiOPC9pxQAYsuychPVtKApmB7361/mTi
x5OkTPsypjFwzKE60JnD0k9V+LzlaSujfnuJ8xBrCrHJKpE0H65M9kemKDEcr4G5NJ56Js8SJRIO
UFxFg8pxOWMAZ3T+WK1isJ9uV0Q3r1GxFAt/sdTm01wm9jlLKLkLDTpV/lkXvYGgvLx+JHcv98kw
/Q0ER9a4IH+7oyDe1mcc+iLZgA9QxfcfgmGmBsLC5IGxpc6vm6OD+Sz6Jgr/sgFM7tCsIn+0IFft
Hpyl2TpkaG0q2K6bYsWPIIuAe495nBGe5zTHV4WLo0/DMw6iB1UQDQN7yfeuFf0JopqAcK00YtGT
yNxR4tsStqLlm6NXe6RD+N6OaYePprqPyI3Pw7iR34Kbz2ct/eI13QHw+gVZ2tfY7+4T3ZZnHtJy
tFEVyD/Qsvol8jbZGooypLelS9Fw6L9eS0Bub5c8rQCh9DV3jbiad0OuWU91dVRdfBf9MUAa2B+8
X2uLA81NjfPPspQ+4YU/kP9F2RT27DN0EFH0SCBw5nzMG/30TTyT/lhFldwpJHBP3Y1jnaihryNe
HmfnK8K9jGYBJQH1hHVFRo2QBItkoftUNAQPfRB3XIVs8E7YdwcqxUrRiJe0y8jyzJ9WxdBm5BrS
s041dxfvBp2qT1mvOB2r4grN9ejYxMU7usEjIouFMsktLUwt8QdE2Ep8fQ8QxIrnvR8wVYOoPHca
7vsI4ZYDwTntCTQ8qwacXahF8yFALwoVpqM15azZvT8RR+j/DRryIKFDOx7oAbkph+XfcTe+0nsZ
NRtAk0RjhaYCEJ0KazuicW2ZXlhB/hqKUX1rcWuqc6CTkiVirbD2bNIU9VAbkJQGl3Q8wwqxD897
Wof16NRilCtqJl1EAMouOyZXPbAVjkGw66YyDFamZIBq5hEhXpwD2lyNWCPsB0Oc+UBPLwnieZiY
43AUgMcndy2CdY4rzreqFGtBYR3zEzBiWdhwak+Zg3xi+BBzDT6J9JEE20V1ZvDODT2DYKN2176o
Wobvol92U2oy/Q9/07VgtBSEDBlxbd6eyVMLpHeDmbpULLbakmIIqsetpcun0FvgcTftzRxnVKIt
pr7/wX1vARvq3HzKPkWVYxDihmjDs6P3IpQrCQcWGP6UBBcTExanzClpkdvYpGUHUu6FqKFcko2J
iQ3r2+6j0gGhN9BBjZ0OXrug8q3pZEMoDlDGgwwsOYZksm5JJRrmQQ6D3q7BVKkr1vEi2etLHreW
ClEZc1a5us72qZbGlfJz/6jq+CCnTuuRwOXjGUWX90sF+n/bNC5tIbil5PgbZEn6CVyz0MIRPQ1k
wQIFWb70gBFJ2/aeSdlyyMepdTZ77a5XYo7JZHGEtv9hI+PD468PRSYc7dBHVZUb1l5nEWKhD1tg
t3V7XQkISEbqaxvCexqZbIAOpxJ47kfApBi/MyhUZ/UsU75AGitI1tqyq3M8UIwESHLL0k6OYhrz
bNdtDg94BDCbUo7UQ7B5DYh4dZFBkyU4VCC8KUqeKWQ2gKWm1ugGf3at2Y4ALok+NviX0hg6Lf3p
2CXrQVp4A3S/+4i7pJTjtjPZPkVq/XgcbhYCJfTwqI6r6zQT2n4wigDTayr6Lc1qHdL5uUHRH1cs
g/K8Wxk8XsBtIHLufGpLL+y4TXqv5rg35mbm2z5JmqgJG4a7LBtbLVlpfKPSEMFDBT04y8YeXJCg
YW3vfRZPZJdFlJMggOw/W2bUHVOjPj8RoVgO1EoYZsETyz98hG3CBiyHxZrknMurzFQg+uuS2KwE
eScQLWspDxA9yxho/OFgwepY7ZptRnLrxIBAGjAzwpmynHQSVFFGTNLy4HBEeHy+fBWALrymAlKw
v3xY8bDV4CSsuL5VQERioGxBrs8pCD20eou4RS6NjJ3IjMX+lj4O7vwE7Cn3XqaeH2dSzoHg8+/Y
aNlkHAl7UOZKGV5pWgjwwwy/YcAs+xZePPiZFpaJyCcb8CJu5Dz6yhJjvngHIoJm55QwoQ0zR4H6
khDvkiSI+BE1sGdjmt0/EpsGPQX9g279qH/tFzdKqBJzH5E9tQI3dq2WuLP0czyeOLwBiTw7BTZX
B8FyjVtkMyOKFKiOJXpjVrCzOsS4Bz1hEAkApCnTM/yBR0LC4JyjnakJdKvT6TelqDUzs5tsMWyV
CW8iMMDEaQrPjvSx4dulEObo89XH1bwp9C0HjO9FemcJThi9SnpLkOoPctzy0DmB+axLV+eA0m+c
dGw9WX4zRQawrIZ/hJwxz4Ev4GHI5IGt1Ba8l/3seZJB6qMweguzqwyP2XIrfEd779njg9Z1k4W8
XYfj3YgocWAZU/NGD7n3XWUeCrggr687mZ0ixONIe/8hlerUUP5+GbQvIqRUVRqiv6RN/gK6VUyH
Png4AJWo8QYo95MKJeacyuviQz7ixrvhBrtFhGC6Qpomw2ESdPUte+/fz2DIDSieX3YXsrfOrt3/
fg8Tsy5B3+6gaDYJ04TIOH8kHJeAIUihnIdMRuYBIB2GtO/3Y+rAzXiigFo+qWiI0rZyuehIhI1W
GHxEFCw7ejjZB5b7gSMf4HFztTRn5cOOlT5kXj4AW0dIDzCc95LFizxX/gK8KeNUfjKZ/IPqJkYN
Gb1WCqPgXQB3CNVzFIGovCmaFTUHTvFOsg/D6OqApRweSQUJg9TNnY0pQ4mFLqJDQ4UHTZFtom7Y
EFiNkqN35NzqZWZnt0eMFbuPgaPsDdgqlb6jO0GOUiSHPqc002mlskZwTq2MC5738qHLGR/aH1cB
w7gfvsQGap6ymr+4BT6Sliu6bkh2B2E4nEjRkFbvwAZflTrrUkH/oeYBxpU4pwSOO57tmpdOWguR
HlSRP+/2VWuOxAapzNvgcBcto742yxubCUwVeykr0Som4GKKSzGf2cS2rr2/2lgr+pMWDS7YdPGA
+QRwCLNP5D3FnB/nM5pEJkwCL69bfYQ3D9KsdPqGp/pWiwaCkn/pIrInSWfUTXtjTHmCfGf2Hh+W
m9LfQHlo2CUYx8uzXPaVoeVc5QNueG8QswamewpdB6A2DHyFLjjckwLTYcM8BIiuCcwkL/jOWmyw
U5e1tYQvhpAxPt2KTlUxLQnF+JThmNgcVOuHycBjX4x+gVB+VkdI8yWojxHa1kajx6ih5jlIdx6+
2+LczVolkls0B8vECcNgTXMRc3CDJtarbf72fX4Uf2cjkEG9aQu1Fk8R727ows6+zEPMQ+tsKgJO
GcO7MfkFlN6gEpKoWv32QjQjwPlik+T7q/CJVmtm1RhYpUkpjZ3OdfNyxBKfffyBY7kTOxiBnq/U
nbZpj6YfSAAP4neTlqQqyzcrixTdBhjKwmYd1JVcCNQKmvKKpCPbw1d4MyUPUPqulz18KHziD8Mt
aPGLoOoUUdhzuEHH+SsBWjfZnL0tIAfSL+hGn4DqotFCFj/XxzPYtNhBoePuKkFh8axB92wGPpgM
v9AGk//VtIj6x1MhurXExcieO+SUzaNANryVQedU2NtASVxXyA7qQgDyCWPJ54MuhjQ1XV0VgVW0
psiHDFi1ybyq+gWTAUuhtAdRd8qrIe7bSichNJpAAJkEu7vyfGMa4aO8Vzr/1sGFh20ePKY7qGDr
dlf2VNZ2P0E/KPykpdfZbKBf1JfB4KTlWeG5n3P7hTFkIGCl6K3IVFfQAoftDpz757sIhsuPYqKF
ItgBHbP21VG1KdcmSBN/QUVispbm/FW8zBfjfUeRz5Hr5CUo82Hma3hlKcoICk/6vKPTYyktFS7H
Z/cZHVLfzotsXtkf7I2OYEIho9/j/01YuDsNNjFY7w9QkNX5UzcgE64u5iS3oEOSxQ02f2K/nTpo
ubOj/rrnJdxBA4r39Dl5Rs4m4h/aOjSSNvQlJ6WWvM3+q7UZGhGtt9NEv3vL+YbVBr7dhjyIXYYh
R406ZOHFmqtZ7QRWolXck7HluM6dJUsX0s4Nnv4KY6OlNoNQTmvxYJc8DlvsKHlBqtip/aCPRUQx
cEVqq9XUAGpN6QTjt9gZ0zsRLfNpyyGuDZg2HOjn+pLuI2Qs0LOE2wBEw6jgoqbgJRqCYBbkXmz4
A9VPKP9cllOx/JLWe8w047FKB/JJDvvRFujVrJtPOiBkJL9eWk1g3OHCal6OEi9iCwXZRIQ04WCZ
uu7Mj+z/ocE7hJPbcsR4n0h6BA1KkgxhA5D2BYnZbfNQbOA3+lSS+ICkZ1sYl/PlPG0uk5W+7FPX
Lrd7XKZ8XB0BfZb5Q8dHUwCtHyM0cSAF4LRcvkqL4LUFoUJTFqB94sIFm3GvjTY8/WoWAP8fM0jh
gRuNEnDfvhV1NQGfEDDWZ6bVcmtiCpbg2YAGrUc0L9c7MZGisG8GgXT+AkPYzVgDTkncUFqOTFd9
FQBvBaguHrhmlYlMCmSYtTUd5XieQ7krnDeMo7L1+afClOzq9UL98mkh2TgRvotcwZG33o/9DbOy
FcQ8WBZD6hXK7YrPkAeKCSQrL8NN1+0Bum/aRl2RP4tF4u+v9n9VCQ7OSXr6P+it/ktcuwMw5YVe
c5OuawF/Tk23be+FmZXGQYMVlM7fe9X7NzsyecpOkxTLrqwBYDmil9VMSFLaUNTa1f8dvrg1pP+k
GjBsL2siijc/k2F1xHk6GZTaYpEwGg+c1voyXT0nLM6ETc1wAGJN9qMgSjNzjsmKjppWGqUKqvDs
L5x6r2cfAxIvGNHbtpm+jGgKusKqzgjAF9yECSIj18IqIDkbYAUfpxlPG2xfhvUHpqLl8MC8SukM
G8mGUO9ZwYESnvRa8LE3IRUBjwuTNNpFtd+X/d8gmw5MX2qYVRa0LfCb64lkJxYVaJfsA+kohEVd
qWKQrRPYunhzZWZfWkhsKXrBxV9ajPD4d3SWAZVKEXoZtoLRP6laR/bE6tg9TlsFFrEaw42LpaQw
RYO8m/G/UyS3ks43syIOJRFezqKOPJ03jOFeQSSbKi2EJUj2se0QEGaZ6d8z42rhtrY9tWJRu6GK
b8K2mzjYq6QR0xD5awiQBjNEkLDuZd9mxmEAPxQnTueVYkAG7wIJQ0qGRWzNOUet07mE+3frbeGX
IxJvNhfVlW/VXIkzvnWhgiVkVkaL7dRwVabtMd9BLrTPPH2kjCdgrLsncatQaKDyZfKIGE7P+VBu
xr9Dg4O6jg2/mKLp2LgpolJlW14woKHgSyAC4yAaTCYmgVCObf6iDaZaWeQpIskUmfVW0R5GNEq2
nQ4dvb1NfKq1BH7+tobBGS8PiKR1GUHAdZWNc/UuKsuwHOcHvtkZ0N/nS0ANYs9vVz+zmtFCpx8O
V21wjEDitnptkDQ1Id+roAvtGg+4bjyuRDyK9NyPuGpcvw2eQhv051pzR5w2rDmUsq11q4ZfQSyx
SkJpRJlvpyFwbhE9mo7o7YAqx+flx/ZtnxKaMHD6tdxoLMsy9Y6bDTkQSja/lr1jiDrp+EtHQrlf
3v604kyqXesXMHQkAEk1jvKSr4ouyNhmhvpZwzf6P9Ui9YQeW2NzQqXPJb33n+BxxtKgxx1nkYL/
hpuejLWpicHsFWHWkXYgASps2Tr3SDkNmiVJvmbIlnZ89/px7mMUAN7Bo04WYeqytA8QngnrijnI
UR3WJlkY1TKgvn6PzZf8n6uRosvuTlciIjfLWGgVMZjiKB2OZNz/FPyaPENU1uIMxjzYKV2QkQ0R
qTEvJhR/Pv/DFciaNz8970nH99JD4GxiXQGqxJvvGcigW7cI851uWRdzG/fhkZ/fgaz7Odv4Mw2X
wU49hn8Fagf7euyXH0JpT8g/L+x/0xYT3pZdofG0WE4r2amqtXtREkUJc0ro4VWsvbiKu6r4/thl
aL6aYSd2TjHDE0mPQbqBWEvpmLhuWY12/9ebahsV1gdqMy6Ej4N0feLIr1luUeiUKjoc6ubi31Hc
aQQJo53W8xGSOXb0xMJBe1y0rReLd93iF/Lws1New5SfynHTIZdbxY+crfsa03gPwO+0fIHU6e9/
8iGExBAPIfdfsWqnas/BmPsrw6IghSw90zrYcHoh1W0dzUWgU9Cc1KXrNo4izVGgyqbtsOVcSwHT
1enUoz+Bs8wEA2HJRJZRqJKg42AJ+yVVaNQjW7jagKDzjPaJ6/NptExAC852zp+2wK7Svu6GNDAZ
iGF8BtxlENSatTwxE9yFgtyx9ICYbPYoi6kaxzF0qv1FZZfVR8KQpptJMoA/1L2InOhqjaNQjdZs
ow+bfNo5jo9Ycq4dqy5uy/aHGTXq7o7gprZtg6uBtXs+GLUSNJ2+J8EHzu1cdI8Lb5rr/TA5/702
BsuDtjrmgiP+UAxJsW3tnL46oAuY8AYptfo9/wg6gZsqzpuq+XS7aEs9/5044QrucK71gfScL5fy
99+05crNmN2nseL3CDwT2Edzt61mTQDzDHjDlbz9nWpitJLmpLje4HxTfwFKgec1Hz4USOpTSu5d
PPc+krKTeFBE5Q5QClNbzluwFHDbDPDZmHW0U6XyuMGWBVeUEJ4AM0NzSIsvbaHIvqARgF7Dg/bI
rE0rVWW4Hq/t/bRmEypk5l3Bp0ynf6sL1dINkxqOt770PEeGjf2/kmABZga1x+/9V5XoR7dVp4pv
jCivRm6dFJUU0IDwEIdtNHAxYZjxBpSs6sL3oE6QJd0CJHYwT0+baovzUULPPW5xR6pFibv/c0K+
DtSbhiGly4ir22dkKblsIE1FrYb2V+v2IEd+W2/EZd3joVycdmxBJyk6KOTnDU+WG1kYtn6fbR8T
xc1uTdvCnRm1lGmKGM0U5QaRpcLveL6sniUWwADjfbjF1bP4tEGaq1zm3SH7Kq7/m+PxEF9QJnql
AXWYmVuOlsoD4S1gvqL3eP3tj6TwVleqUajSaVQO/hpBiP6WJmPahXOb0mfss4Rk2bEvOlUJGG8+
Ad1iapQbWxDyRYSw1h4yXfnEUnIHAXPJKmMNYkccej4+uvJWiJt1/KIqU9HY5vphOBETQmqBe1Si
1Gc84fCeZk/5vlw+5KjsLaOf3d3uF6T31VZeTNxAAhj4ZecehpqaSADci+7iqnua28UzCuk9tomu
TZRUfzVbpETvE6F+1+IhSE99HbMo2jYdllI9i7hX2brkEnWAFDIsswuROftv5Q86YjbHmTTpA6lm
c3lt3zY45PM25myO6/otClm6+BxS5jJR28hcSa1SdG5ErIlOjqji3OyAWnP4CH+xO3NmE6GEs2yB
LQGACaTnzMVk+HusABmDBPr4Pcp5DU/hkVTc3c6QVprND2T0Qep1rY99sPCGXGGaXODlt9rsEiGh
aRR+NNO65fPzej6i6zzbBaQe0xNMWecKcsZcmRq3/odMlF7WInkzftYfJmTXEXAxyqdbbzByxtB/
EiA7vfx15lkxFRwnjeKtxNY4/L/gMVMtlY6ZQKfuoENP2arbE44qrFAcKa6U5R9yxUxnSZyZp1sv
soL83+ofSVVke3ys8gohi1+aPQDgZpKzAj5fHervuoybWbN5h6Gw9LHURYA+7iBZHJ7cSbrT34Si
g9UQVxbcD6gP1728NjHAHm4B26WL3TyxEOzhP5plrcr54kPnKCw1egZHrEvZtp057hJ1VzZJy1+/
HWei00bf8PIUmlfpScaW8pgiByOwjro8fRcvpXFN5xgGVvTXaDXvs66kwS0V69TOJPUiJ5GrjxQP
2DMpoI7cdOlrkp8gf0EztONNtnFXaMN//m9ctGGwC2e22iQQlXupPsGy0iZPqv6Z/JEAcF8YuuMk
QX6XrpxlgQqt40pyGk0ET2YSgzn42R2JtonOEs8xJIzaPxnwJTVBu/s4P1IBQcK/4c0GdxXCJ90+
Ok2TnvnLeKduNCK4YZaALYk0kkLwjjKN2YFHbT/vZfOnrX5k8XiaLA2tEIcEQC58Xy9lLjwjOga2
akITw10WxG3oAoWkQn2SQn4As2/1YWwwlrNebck1aP+zFuvq2NNETuX0bKBrEJHdjnrtnyhsMdlY
meGVs27uy18WtGgRUE9aqFmD1di93GpIPPkGunODxIXzAqfbdsA5fM4+Mm1xyOlQr/h0QkNLpmop
MhGrVPZJeOgUv8yHnxP1g9NngrEp9VmxuP1dZY/bTAK0PSePURmpfSIf0c4QGXZyISrHwLA7+XKN
dBX/HtQ9g1zNEJrwRHfe67/KbdwMKIdR3U99xGRgiC6EJ9hsd4RYVAH5g2qjZCpv3InIhaiHgQ+d
hTQQydRgJEbPD6Idy/XcNz1+FIh8CjJFo5u86Pq1hSqI0d1JUZkHbUX2Hj28YEeedDsWNg69+SVx
XD0/Z5izRG6Igl47omb9ont/NpU3IofJqnDsKTeZpNV6YUj5WH++lGPhhB+8hPdmg5jp/1TEQwpT
cVZpSYeoO0evocQH43E/i1HBLlc5UFF3jJsKWMrklj16uaJ9ykzbRb2t1EEE8JpcnaNkHQrXX080
q/bp6K3le15C5Q/tdhC6srK5k6pK6UlRe9Nh4s/3cxfabMhRIHAIdExVYxAYJ8Cm6zGYACaxkjBS
KnfAvwB3E0CV4VldcoxvtIkJVbMcZZHmHRlfahJGE1ns7ZZHWRn6E4a9YMRmT1moVDhcSbBVuCtH
qrmByP1CnXR6iPF6iNAa/jvtriXMEd2CUAAMppaMX7DLSTElcxTqbPM89P7lFQ7kTyCcTY0OYEts
IoIg3TmhlZ9bKZ+JB2QF7oNfAR/BNuo3YQZFD7O0+gZiC6AAiVT9VmHa2eeiV9kD/H9lfYLMN4A3
cApVxXY2Pzo2VNk0PYqTKzHQEotwSU7YSQqjbD6/ZL0KnubviL+T/0N8AAvFK067oCOFP6dhOw/8
FAZim6hjKbYYFe4CfjCll0Ev74gxdlZwGjDKfwXh4Qij+IMtBO/E02kVwKvvLJLncsQJ1ODE/DXO
zilWpQjHSfJ5ayS/h0Mz4DVFaPn80j3B3aBwJ0jsTEpUFAG18nhCqA4Sv5hsxhSeCZNdraIGp2D2
/c590Hyelx+th+QOa7hfUQCdiHWwcpP5iDtzqrHQRLUSDJ0/T7KvwEdOMkl7ViRX7mIXuOQ7KcQ6
goA2UlPy7FkLqbCGRrOCfpR8MAxESOBZDdYrqPU1jjMY/XdHtJg6dl4MGIBHm+3zsIC6TSvXXV+G
9he7d/WisnKN2AIfz3qarDqT0UFV0PfO7sKFx9kP6SonS4dfNwamCo3ptq6CjCGGcMNi7XPxYuRY
37biswNGJNy1rgkAs5iav2ajooqH4rKKGRTrs1NoAfurJYiEQ90slgTOvdGB4k0q5EfPZW7iDny7
EMqxbWiDDnjp4WR4wsa5VPAukCaFgY6i41iLjn2chltdorEOpo+LUiOLjEx5H/9i/5mMBPxpYXVr
gEoZ1A+qy3vaCudqLwZJjrlnInOoYorW0GFUwxCcapyZ0AaY+k8VyhNm6cS/SWDQk6/uMD7NwW3T
McsjHWW2eM/lX7twpcIEnNlntGY55TJHziqiHfblplNFq4AWRKbPJgzJPxyAzufU2QMT9hMF7MQB
3jlFWkJcgbHic8LGTgvW1E6ij3II6W3Hm74B2nbPRxZU0dGVqLBcticNJiAjC1d2KPNy9+iZAds1
0DMbTRoyBTOV70j3pAi6mbAi/Pn05A8I3AZLzk0W2GT1bYs1utbwVR/abNWCNk8C0Jm6XSHjeGoG
hG8391oCtBQXY5iNR4jCEO2TXsu0kaKFXT1Ru7EykjkDTX+REENXYt/tcr5n/+/I5xxq57ySNIpX
6RETUlQ54inxQXtj66BQzZa1q7Btg9tsEUmgRqKzPwWB6Gf9OsE5EzVDP0inuAOzPi9054nC1Had
IwCMfxGe/THb+wdb0C/p2MStbhQ6Z/gKmiDprmDnd7ZO58aOdbFDUdKkz5NIOA7uhM9DIDoIpkwf
uN/New4NLMd/ShYx+irHdIzWee4O20cnrEm3zwnawnSNSPLMJ95TS+CSMsmSxxsqhlMTljC+ccLG
E37kpFvP6mL93ra0QvahJ8FxEeLP94iLXlAv10yin1dcKApFbZ3MA7fUzm6jAfSIbB3QW2mCi/H6
iNfmXe6IQl/zAVZ85bSdLQpcWlg3RWqfjtcBy36Q4YPpxqwayU87I0WYyp2xVNWOm4zWluvpf+0x
ZUAteEblWY9dSdUs5TNwx2n1awULdI9/MoBhJHSOW2YbjgvZ364EJYiIE9TDM+L+yi1Wks2O92OU
F5AAQETQqNzeB5LEK92E00A7WbVStoMJmnBJYRKCVmEcrib5jw+se0aqGRY7hcBCU4iRnETIwb6I
hfB9H/s3QrL9OJfZc8u/KBT78wcsM5DfuW9x28IS1kK4eMWmMSAN31FFaqCgdy9GQOSe+69QagaR
YYybFWFwQdeliXfh2mtVL6d9ljulsB+AaxEfrBXvzNRCNDlQyKV4DYUC7E8SEoPop68IzLO5DyLj
E/fbX31FPjBDGhL2RmaZz5CULS4yZN8qCJpDvkpdT6oOdokgtbGvF7lOKts2GqdCe3Gqt+isZZmB
i07Jk0p0Cgrg6ITmHUIvVyo0c2uxBWHLmFfPqOr7gDq4iUAcXZ1MnIDWwoQHmCA+EOd7TvMa044m
jb4dE7RLjB8mXP/WzZ16vkPZu888rYjXR3Ezv5uyGf4j45oSFw9wgeBl61bK6rgtONsaeZSPwvyv
F9gKlRChHKaNVtoIaCSmmSMbU/jIwjZPjvhmhsqgM0opxx2e/Mf9Y6KzSekRpbIO/AZvgOcx6vys
lwD0bHE9NpQjol/3FjzZC+j3OhflQw2dypgE6stXT4uUXCcmDfUxBMqbZx2RVywyT+xXwXbZ3V8R
pWItyhQyUT+v+hjP7ZnC0mqiFDsh+0RHPWZBX2Fd4YwZSy7mEgdTpDotagkFKN7SgNF+A9cj0Y9X
R8FZLfiP+3Z9L76cXCBtcR4UzVx27q3BYvybBusp/quHNOVXfI4OTYt2KlEo0/6MVswObRxlnfp6
g7asO3tYdF2bio1KDQajpmo56+OUlPqG+hTssqHwN/2ZxYajBjkWR3AxXq8ATsZjP9NU2AO+//LR
DQ3gAukMaLze570B6b/YdwblypTiyIsdHlsZ/uQEB7FRacGV7B2hYtOZqtNMC+dUnRZcCGovdf5N
V1om+jvQPWQ8WKttVXRL1KwATpPe07ie1N7khXlzxIY2vH3pFQ57yNtGmHVBeF3ji/Mso4ydfJvL
66DH0ApRhRKUH+GsJVJgYrMvjwHTAMBis/NsnoK/tk+SO6lbYtLBkQOA/zElG7Lbj9J2HQBH2NiH
4CUVDXeBUxAIAocxsukjoi/jXM4Iw2UQgSQTdhePbffpgLV49GZifSgrHhFXwWLFSENwAIoUcois
/+Cg+sRIm03G0Ln4ct6g6ofbVLusr+7jaZJNBZZ3DugXbZk6n2Tm0M4SPjhwZ4fMHr8ZpZz8ajlh
EAAW1OdbJHsWMZ4pykIx7SPyfvSIVHU7IYty+/eh8gQH90Y10fBWaRLJAsr7z4q8dK/equlDeIiZ
isXPfx/JwEIcSVhXYwuVbJ7EXxclY3+RtZJ9agXSwTVPUUBUXHSrrJSmUcanNnDAp3RxOkuS7wz8
dxZq3aPOWUXl0tTutK16z7nX/WMJghJloLH+mwMccyMS8Qz0FSLi4bOt1JY3NmlIQkTp9WKZp7DT
3HJ46/6AmiQM+BTD0MZhd/aJGmGcvFh/SDfFUCfrLdDyH6thNvekWdtssIHlm1w6iQDDv3wGJaqQ
/v6HiRAP6lCCRwFuZFWohEUzrLxZaMx9raAFDdI+/3FnmpDDzQ2zvJmKC05JzYd9j6WV/12I3X9S
18NUqRLbOJwm7YwdWon+j6FKVXjg+W1DG8kGCuK6cAjGNP7nT1/eY+U00wuTeQS/2a1appHdalqN
2+kbDdaNx9Sk6Objb3mANXhm+fGeY7gb90/VcbqsdO4lnYqyfzQzAIl/TxEPBCxegHpLACVGVPbO
WGI2LmgVR7phutGAcyqS1Bh9JbRWNA2RZmrX7TSw/pXSFJjsQGtqy/z5u8U4YmlJXiq+nNixtBSh
RvfMl6hfHkiQr+BWjIHX/I8QRrskyjPz+D8xbw54EseQXQakhfiRRwSYIQtOlpE4T/GQKC+g2Ii1
e2YMwseY9tktQOPAqNC6PnpLJxwi4jeP9tLfR2uFe28oCaAswUSyBzSz4P6idTkncfwIH0bSq6C5
wjAqsunyaSONhid60YQiukyeSf+A1d+C63c4mwz95O9/8At3e31MakrAKcT4Lm4TsuAXM4/y1JFh
GRw53H8J/0ku9Gr7ywm0vuPV+/w9nOCNZeOwBRxa2nkVjGJWafMBCDlhcQcWlS+kBBHmz0+Kqcc8
MdTkGEt5FyzNEgfOqE5qkVG7Sq30AlKFtBLvhq/9sdPcfCnxEbdWpDfldZUS7X1haJmCSMhZqd0w
KH9qZ53k1fGqR5WADSNu6srQEyPQ5cdKQQsIJXFXMz6KJPibE6Ixw75+alBSR4Mz1ge7GMM2v8TO
yxY8GjMNKJ/QR0MBaPf67zjgSrM/CHpuUlnDafNZQczkxuQkJZ/VxD9mnRdL0TtW1qfKl8+DekdD
GY8/sct07oALQXHZKd+CerwbiEQFwZZ4XZWezmr91TBalwtNGrFCP1gAaNay/VCTwIRe2iG/eBdZ
ke97ArZOv1/sCB7tPnjHMKbiuf0kpGiZPFnH5tSAXRh7jbljCXo+Z1Oo/FiT89MY+BaUS6HISw6m
MyHDAUbCNY8ZOQOUaIlMAsfcOEv7mV9ciKemayCqGSrprehbT2xynvXNayyTb/gyDqR0wThy7z3o
5s5QEhWYjkPqCenaVMFsAYUr8Bi70iN6ocXaEIAOj7BRIjbbE5giFuQhjkJvVCDjBkmabmOHIfIS
pOkKQRsrG+6FrgF/oS52wBaydivyz5SMr/ZNI8MUIGYr9l97zHkvDnLcjOJn42NLEleFEUFpJy8S
KwpHtb7dOr9N/sWoMwB3p8l4bcwoIuCWpqzFH5KXojicYi4GGS2CWssrZFbExejg+6zI+9LdF0Xc
Z7XLr/WT8imVUkn9W+7ZFAJ/Oh48FMVhB46t8CU/3LzXS/vNAyMxmbCWR0Fq1gPA0uJIKxu65TzQ
dn9f8R6mfdG+k5/hCn80KOLSjCd+gM5W4ePOSoFDfq3vmAZrWdFgduEYneZgvs0IQdFceXy8wKvj
5+6nCbQrroYKqq5YXnfOTVz9C/RtLJiesXrJk00h+qXnmJdT0Ca1qQC1hDLRrBbzeXqd4+YN1ppS
Hr8nungZsaEFHwepXzOCkAEDUxJKuaIfAK36cWnCNWrlLCIputH/YG3qv9UZtwY9z5t69k7aC+J7
s/yM/JSyqR+F+LdoUFQRXkpzmISAs2EjAD5yPeHknLNi6mbt74dV8EaZxWdBDW9b6yMTrEU1nd1T
zz+tqZaTwyts3Ie37o65RB8e/CbOwEbjaEZ8KCJ3rdVZZj5aoou5yej7GMllNPsTKlAqb1A90eZV
cK1XYwaLx5XxyrPpz06OjW/LM5wFE6ncqgzRXoqaaewmt8gnlO9KlyVfuHE3szVDB14L1c9wIdws
QDZXvoLZiIkAm1Hr26fJg7O9Mkm2JtgGoLKkwbxnA6JOrYX1JyV2Zx8QUTa+nhJCX1eodXPfpg73
c3yoOZYLuKxCAnxRWESj2pK0sR3FUbVtKBLLksvIZzySL8UyCXW5aeJNtNxXSGgMnWW57Ll42Oou
+2RCiChg/p2hrZ66nDnWIF4mWl4g3Gqzl+tIF3eEP/L+/JUKrlGiBGfA2z4wui6yZPbwR1jfAboc
Cu9PDzcF14nNRLThL5qq7Vl0qfyp7wHPPINfdSL6QFFsODSlw0X8qZIAuw7xxwDqsbq4Gqars+wI
gyAm3BNDX2MsnnZ6V8pLey7dgMt0EVs79MDWnBh3mfh8EX47qaS05jrRD/5VE/NW8JWI3OZY3oIH
/eEPh7YyR4NtRWCTlR9+QmIfvXpLKJcDBV4r77TSbrAdX8CTqPbCN8WMIqxVI4FqFodevFNqSEOH
AU495oieYKKvBYHN8Q/zxlI9DGIHTmHfs1I/xztSHeDzkD2/5MhFyi314BALIWXnLqoctf6+w/BK
HmTVpkZOdGQaG1jarISm7Z2QWQ9PYuuqA7BfwRcu0USWvqXLrctrpJdrI+dTCpJS+qZjnpvHEzOQ
GuTSMnFf5B218bqHNVv6yiBAPcdTcwFxs7+roPq4IdQkNyODGuR5fL3nCzJmaJT8udaLOsoL2hGO
l0vyX5/gNj5M19rTcDBeT07iE+YBfn0ds0qTxa1641b9mI4L61dwkqekgIA9rCaQx26JadBI350h
BqoTA7b92swkWn8cTJ9B5U39DI0d0d02dFTQ8wymLjs8/nO5lsZVnOWXtwfLA6rzRV7T48Jrq/KI
Gu4/4kp1OVyItsqHva321ZDy7xAZ0pBUSm5t3bTWjFjhBiHccWnCCrDUHQtAj2OrKeKC9ThYYkd8
Ls/Y0L1Y9puqqEF4uX8gydQIsfQvbxBRkz8lX/L1anaJwezafGpbfMaQjh6y59TJpKX36hhcFw4m
GDXSdNFpb9N4nsDyGsDNuCq18tvDyDrU+gH0dwDUuHcpN9boepDHLioJOLZoMmIKuPs5tbzBYvgz
H4WjFxwZ6xqlpTuVtNsMlJ6+GJPLYi++uiIFhaBtPG3hyEYKnPQEm5Tygl7GvmQuzE9VFvpVE+Zb
NwJRgHSsf68UXvm0P+cJNXrMmymbCVFySmuRweTKW1jTX/+VGmbmhc4/KViGxQHtTcbGu4spyvjB
XIMl8IqkXcjHZJy8z2aLF+GxG30xLha814uiAiP+d0r0vq0+blOM380Ih0c7tp1r2fdmIjBvCcYP
ZMLaEglw1L2dfCvryS07fxb5P5uze+o9rKzt1NpBmIWK08yI8Pu3ybX37eUzF0KxlHxwSWg1RjDg
VqbZAoW6QfGSu+Bl2GSUk/dMKmAtsSnyIhEmOJKrKh40p7rZhNpwYOpS1vZcZXO5ITkg7hKj+k11
a2/aWrRAbmPEGZo5u1n0evk7JrvsQLPYVJjZmdWsp5jq/us9Wgq1d0QsnNXdceqoWjrQKC45ISVM
Mbn4gmw+SNANgd1qzHa4OFCMd3yvrQOQfkNsHbCQGHOTh+NVSggbVE3dECrAJIu1fobfC79dbXUg
pcvpo1tT2f+JvwJ+51uPks4H0M2jtIScs7uXtanZD4ToSh+FQjGCTd5JHJmMaBTKoQ5gcOFjdxIr
laAxLF/lYTDW001dZ5lJaeC8Wqd306WEETunUNWX67NNW2PbUFfqRoNRC/L41aIrzS7ktB+VrowR
FEXA1yQbxkR2OaQztzQxDkIvapf68ampRP64hH4f/4mJ5dbXoKgb6zPCeOzhW1WtotPrDPM2IBYT
lkrya6WJdb/j102vD0Jmi1QKU+GYiTV1al3jPBxHT+xiDjFggj3c/KPOFFFK77XrzmRjv28TalNr
vp7YWiFXTn42dvm1PURTmUd6yAhvAnicx4jldzbS/SwuvlTYUfPSVcZWq1kvfYsD0aSOcOBUamkg
O0GG4JEL5PrAItXN8Dx4dmA+zSzeMPmD2oZH9+TgYVceFkGNrDE73qxesnyK3NqxzDynkFp7N/5Q
wP8NxLvYwuRLmHPTmXDs49yoMJlK5csvBGVVQhqbuSc3U3Ev90HUvCHZX+5VROKPu9R/p5fAbFJz
XZwLqhAVy3icb0tXsxszC79Rr4Bo8iv/krQ1FqdO97ryGjAyZIRPzyjeQAtgd7LcsXM7uL05c4UP
4x2LChhs00v20jfF2H8wyz9x21t/S5yqGRBgnQVUM84IcKbw/82TNuH4IGQAOJTxEQJn131pv4zf
gPcUqVULqzVIAkCRa2KIFPU2ksGQtbo2Vao0qZfcSlUMdeZuV1e1eeGqf+IEiYBEDrS8CsDZFJYU
wMioSZ2YeYLIYXJYUdmZXR1lD+1AVDKIwn0j33zSX6cbPzpoHR9An5AjjxCyOWUpBSECqewXfueE
nKYKjcSDg2caUOB64H/lZjJSKqCWe/KozXJhwemBXvSC6xetZnH6VxiUJMBJlKhK65k3uWCOPxmA
vBBfb7MknMVBvOe5SlSgx13YHEqyBvZ2eHZSPMFA1+PphV+hP1NDTpRNEPiUO2RvG+44ECZqsqR3
5q07ZXG8efV2S1kXKzu3gIBdjuk0cE5R40DdaPfEt2dpRn5+AsQlAgYP9wDY3SsV/UaXDx2BC535
GHTwa6AxYUbceSx8qcqrm6bfmIVUnR4Zy2zYIEFcWg5IgFQdUsCbbPKoVZccR0vHlLUHG9gBZXeR
j8yJO35xKoxgz7iYO2W8p+TKJjuOjgjNt1ttWkVCchkUb2cZpZHU5hsBH0Adc0Lp99A/1TdQIOsf
nAiMVcyTZBVVlYlgd8VOCqOx7eoBbmWUjeOnWmlj0EBJ3YYVaJjUuearVpiAo1vTSoC5igAI6pKt
T5llzVukTBG8I7hycw8ZiBJNfyi6Mu/CDj+o1rq/s2Ud6AtKOPy3/fRECvc7CIMPpoKFWVFC1dfb
uTFDoH8XT8/61M3kaEejtF9lXmCxT3e8b7JnCNWdL9Te3QgxMWLVpatOENSb95YIGtxG3Lz6MLIq
oCxFr9l06yHzptdeEk/ikOxctLfmvZPlluFFsIfyYOo7aN9a7xjA/6hLZFpXvadTdLx8/6Nas3CV
MB+LMxYY3TpJioj5qVvoBo4kXMbw+tLbhbmNfvxFLm3hKcYu/8pDsk0G21KqShFhqd9QVLbdn4b5
QlqCWO5XQuF4gUUW4nwZm6pf4N9qoOCpkL6T8afIHp2sN2BTPu1Z7dvooOV0Pu/iDYibmYXZZAFt
DFwSMd1kQT8ZAt7BG9WYwHyBjUOUzWZ4twnMMqX31Hwo8aHsoOIex7XMZ0OVYhokOLeb3shXWMUa
BQsIQe1Fib6BCacyqOsXZd70hqrqZCBKyuW1mz6gWlWQYHUIGUGME7v9gFC5qXFoWjic487Xkh+y
GJGbLBGJZoARIynpZOEzmDWXjiY6ZaLwOxaj78CFkf4hi2xQN6menUfvBYpgoP9owdnZb1b9aV3P
vIqXVHkssYqbf0ROxXRQce2enTkl4iH3CkCiMEn7GpkfMCk9Sy/ARreygDjwBINhHHu0xc/Ksonm
3XVAu3E51Isi8mDpq08vWw2XJszboUKi9ZzrzZBqB392WpaIF6+iOVuThWALZL28KfLoOTbNW6zi
Vdp8ZtekBTiGCrZcmAWkp7TusfsURPmoabuFg59sNgqF2Y611ukA3BcMyc6FlNFAy5rnsPOmNfMm
w2iyM6Zwiwed08UH5sFFBTKcZTlYpWqvGzQwfkxUGaICsk4KI/RoPfo1fmXy0nfpluBxQdfRJn56
dIjzYYv6XZpzdoP24LxB4sLCKUhF4JgUGWrJipM3IF7UXcEnLLLLfWbLaRII494GtQgB5IgxvaUO
h0gGI0xEmj2KAHZ3ZhgF7KN4qI8AukW2rKm3rGZYR4TXZiB9GkKHhfgwnSSW66674AxrFrTAAUo/
gAzqaSXPlp7mlTgxQ9wxszZ3EJmb2vLy63FhfeTclJWoMlSvfFpBOVx5Z5efwVyTrekv4OkbWGg1
kmqnSNOtQy8e+FIh9qffhl8mW64qW4E7TlKOQZt8NuVk+Iqhy9n0EvO/cQLee68O1lXHvUTDev4U
MFaZ1/DFOfvy3bThyJqFHgWxlcD/2raVs/pfpEjQ7yY18kiit5eCVuo0FTmTwDnIu271WtbCbzfq
k0m8lYDQ7pYG/IIsdu09U84DyAvqxCy9eOlZd+Wam9gvE3fkgfnWtWcXiMryLWbCoxcjPQaJUhEB
swQ3ooSR+3mlvfQLGLdd3W6KLJWBWh+ftb7zg4dNWe3mzS+ThynQud9mDWgPXEvVwHP4AhDIw5Ov
Yy+i/FUyQLhOs+I9fgWJ9iOr52i+dfLaKqTJM+KEcKrH1sK0TH8yiJ892lh1ppsDRBgiho7I4s/q
YcyMyh/80ytjl1Qve4e71zFwlswP7LDr9CCsEyO/hagLATl1drIX3Nq/xl1j0vFUsSxhgqh4WWBd
HKM9qR0xEYalW5ZKaSapUZ4B1nZIs+tJNExfipLaI2vkwLhR6eAydB1+oOIlwCGeq3DFvhKdaVvP
tNC5ZtjFbY7QFeS6KTlHGuwpppGsGPNOWLAeDeZrdppKpQz2T14uygd3TnF4NwOXuRoresHztVJr
tNpiDBztpNhrsUdTeg3Lj5czsO3danQy3S8+RzUFUjvUuuNBYBHQdb0QxdUXnggKoTiVGMqJVNnb
TkICfg6jTJJzitXN+6TrkEJJhnFaQOnkaTnso2XWZAoNS8WzKy2QVPNgiFo33bMiGMNJncLxj6S7
NXb5rqdVWoDRUp3ExKSBsLP86tafK8GameVUUHxYEnp0BYZXzfIUBMTfY2tHFPc7V84RhJtAfHzW
vK/KtBuRKpAZxNM9Ys1r1ou9hDY4puHAc5pJO5qks1Fu7w7SafZgweCyrziUL2M9yY03p4895PnH
0vmrm4KRjrfztjn/Ta7/h1LoMT29HU6RgxdM5lTOReAGfc7h0h5I96FJoleHiXX74MkMDmyZE7/7
SbAbqIjB4iXjOdnugdGhvx/KZbDIf9vMvlIHHnph97zMJdYDXoqayrQhktfbh6cqJ8Dlm+8TT5HN
zWEOu9x0BEHwRiAO6fNyg0fAkG6GXN1RqZl02Ms0lVnp7CA2pSVVpw1mKuy2HgNzDzMcfok/m0im
oO1XAw8MN40AO1a4ogTJuqLfIwtXKRQUgOPwVxAMKiVC9MunGMb7juA6UtNX0MdVKsjVs35BkD8N
QAx/7j3+I3Achyoy5/KStCWAv3sxFYObnF0KSPvlpDKfCz/SPqRLAMTrUMsHOLU8B3E4BHrDScI4
0bItdQ2YVW1o7bycmsh/8aM/XqiV/vA86QJVjlYry1mQFk4d0A0BELAv7xyGrP/BB+080AxE16BH
L9pA0ol8Pjz+MK9wN26pAJTRq7a2hp7IMAq8TuCUesiTzTcaIJL42yvht5Cye3clyJQisC2onN78
tvDIgPQK1lORerfX3cBvjo+8ASfTH5FHsspjyY9dkhYI+gmFTHLcmZqeSSlj/NwQBFcBSCGzNbwe
HyhYj/lAMvbbxyQ3d7M0AONTjCykrrVIpzhZXU43QCo+b71glbhuxIm22Fuz8hcJxKxyHDGPLkd0
v6+ytOOqWkMC2io171il9lddryBexo5tCw79wJGg6nvnj4gul27pVb/vozUcO720xzMXlHt13rVg
C/+A0NiRiG3i7YzUreD+YdzN/rOQnfrXfcnCCgtqeg9Ix8+nTkPBApuucqM2Y66+1ycwar3Y2R8R
Etp2HQfX+UYp9xFQV8IBeyZHf3UQLPOOP1aEpSyoTXetBM1A+Bm9r7fcwkNVHUNWQEVxRU1yFGWR
l/Qs04bbQV9ayhJeIhgvNGK3WgOz0tFxk/Nh9kT0HPabBdPmzbvr4j7EHFpubIfsw4TfAO9PTzpi
q8UYnTxK7xuJqmudelVNQtmrdVK4eADC6fqSGE/ZMB436T6xQTW8U13PC43Wp2oNpQA2WNlom4Zm
PvA+lEjYtoiFX8VQ6bXPJZHobDwuCT2VyurgbriLb+WoiZ0sdq3kXaoRxs7qaOfdrSXuWJdWyU/9
9PnRuBb0ni3aaLnZn/V7IG2yVagY5xa/XXo8oh3ryEDFFGZaKlJdHEDmV3jMxos28CmIDr2T097F
ZoWRyldzC10EMoJYVi1ybQhaaGNcHXqjeYz/OMhTS1Ml2mRynt2oYg6XvtCEOgZgHu5psNk1IEuM
ia2kr0UDCOjgVZg/IbYdafMRDTtRc5rt7feL4K2b4CcpYbUx6iiCEkcqFKE1fe+LV2H02svoQ0j1
JYOsjbM70E8pCqN3Z7QWvVwHsEdt87+ovzM84rud3MzVqp8fI9GnvBrFY+xsX5Y68hk3JkW+pDg7
OvRAR+Z9HLpET9tFK3+deqGiilrEVPLv/6Yk2W7Axl7ISDd/JnRSzevcFy+BtJ+Zwsf+k4raYHFl
RHB2hjLFPsQuaUe/9pzvnSC0iqjSJabqwN21TC7UPcGDMu6H0+ChoG7oqTr94xLRBL7c7sutZS42
K8+BQo33OEIUAd+IIJWEHLcV1Znxq03mqpKV1DtRKC0lYjX4jhOW7jENxbt3fsqHm8CjODjw4jnq
4DfBl8eDGPapb1W5epqGKUOYI2ckEkLm5mHC2dqYeOtywh/lhfgc/LZE4WVJi6BLFSs0rrSVoRQW
4DcP/GZM24faHR4LnScZYsWSZKy91qHMdb3F012DLKNvCrAVHeVpTnM13uxbfNTlP4JNBCU3rtLA
nwKrU4yxsg5UoJVNGT/jGNAjKR8js9gnG2mmYpzSt0//E6R6y9r88LcfS9YySAQvj5E4cr11D835
OJJ37o9Xagafk+uawxubyvdi9iu771mqI9iGDvyYFRnLBj1HRvokzyGUKFemL7acjSGFoDDnyuxi
61baKzcdSHUahYxTwW7u2CTAfkkwYv/WB7xocHNfPCyKpss9ulwCt5vItmXFgsIk0wrQnZ/BiYZl
3rIDOKoUbU2djGj15WKPj5lux9edldIq7kkGqhFxnV4kHIBK0Fie/5i64blTLayI1RjZr9UVs463
wwdusgiemiGflTHOtn+2lcfq2W+FsbQRszxAnQiDbuCK9vJW4ZJdeUNawDTHnGyp16BCaIEz0t24
25hIMIQ2HD/CtN8VsGJwqGdtnJiAHQpUj/cce8ngrjRjb2dBr535xrMpeWWc5yKL4pFon99OuEyV
diL11PGquVNIE0HJWwGJ7ziXCAtBIQKjrY628P0SnOh1UZr8WKgkeupGa3fQ5pM3N3pp/SsXf45R
3YIbxg4yQOw5lHUPhUmFrXn5Zdn8IupPV+mFqvDrZQYabso0J4yZrLxzv83lLNwUC6vQyBWj1fop
aUbl0gdV8j5rbY/v8UOSC/QqVNyeHx0uZwSkUhBrQwgH2ynoEqBstCcLW1o9sLURDU2xiXQkytqC
ZLtE7sKsw0UzcVHaUy5/Z/e+ajNR9hgBme03K744lFkKL4ao7lfnWasv40q60QhmUv+MAfamHZSP
U758sboXc8qD2aTF9VIlCLuPnXW/WmRhNszkOpb8wSlAhzpt9Vw1u+JmxhnalzFcu1Be8/CvWYYo
uTZGPuL1Q2k3cIGVJ836pgyDoU2ATlMpNOTZ5bRX/sTj2bqqvNk9BEYpu63SScz6kXsc2sU6xuPt
oJD0OFffCPN6MjR07LgiZA4oiq6KcCMsDztjHJKHhLSrA4C3qtqWWqfUcC/wzosnR96ckGZhyj3Q
n3XgNgf+h5dOu8KLdmiTkTSTauNnD1B2frk3xCURMje+pORVi8ZFfOWvuDHoC2xuHHqcozVR5sLx
jHXGOfLnSr8aCEx2dma8fGdHnr4CQyv08qZHv9m3C5/FgHzeCKNyUWLHzcfJYaIofe7aZWgsGu7b
9zbjZjWxreaurl3ZnLWIaIR4RFtpixNg4C95m+xTQCM66kMbg654PzOnOg6RAdmxSyNPRMb++Cgk
fIdK4G7NEv31g2ay2M+B5XJPeo/WXuw8C4pwM2B7RRZsJm8z7ZDUbBj0Cgbs69yDjYEWYWQRlO73
juL+NVU1+cc42SfDoAi7Vmm+cX79HPyK6hZVv7JfP7Yc9Nr4QzxUw7lcI/TTmkhU/8RXumNrOQEb
IKPTeYFLbDjeDeXICNejd7wai0cnF6IJGGOqpffCo8yQbD4fmcX24ybVVhN5QDeemo76M3+ai5GN
BU8FtUaR5rpukZUUG7qdLusSe62YABqL6XoRHS3TJlxaB80+vguCmzM75p92YSMKZucIY9sshEed
Ne6FmLidC0OFyD9snkmABxINaziG6DCshVtNNIljh1mQxWAQa6NBCund1HyQ4WmX++eYvYGZwzn0
7/E7rYHEUv0zNJfDm7AghziejMWmIhw2ekNvB3hC/5AviZsaJxO0iGZlar+AimNn1dPyb8UrUZRi
h7jOOcySQd/z9nkySLkAIZObv3MUeTtiLdWKDDBe/NC86mTt9HFvVbGlVUI3vxyCEqLvxSJTlrdb
DwDWHkSFmD6aaaaSQt2AbEe/4d04u58DezWFW9aIIXl9V1IfR5Hmoyox8+8aT5kvalUEvWE+50bT
R5XOAiPE+1aVe6Ufim5/fWJ3mOkuZlaN+7IcmwGR7luigzPYza+Nlsd9UfI18jx+t0OrsIdmu/MI
2UJDkQPHzoYT8kQ7u9L5cZLPntk3fhRuaqhnYNWFowlddfyn1koaIF56r7MGeNp2oGC8SWsU+v5F
tYrei/JYSwzTKS+TrqNuP1RbUnT6jnQdjn7pKA2A6cknnQfTV9Esfy5u+9rCCpPNxbTdfF820gjA
cCaEP9bu3JHG8QRA93EPlqQ1/ZSDVMfa2j7ICpfCyNwswiLQvOumuRPj03q46v5CPFh9FRCFyQ/9
JA8ig9wvk9z+dHlA9KxQCdGqvAGEcx/0G6L4vk9dY0fqP4xak//nmo1mfsBOVvrP6a2lPvKzKMeK
ii9WAXvGGRM4HiFo/On8rySrkurX8k9k2x3FKMDLwOPcFr9jgwg2gD20DEuOkwGRVO2+LsJkhpbI
SOybpjm3bnnzSdQBZ0uwcxYzdHuaCuRX25qrmL2Y8U7TrR0SSdSPU/oh1Yz2DScXqK8FYYU6dcSq
7z4GVXQ6Q3FjaoDqGC+CFmQxJu2GpMSX3egde0sjyUTa+qE3KF+xI3PIKEM4+nJC7Z2Kffb2Jtof
wIn5+2JDEFyAVrFrWG3pG+YNhR1zKnxx/cia5Rwzfl+CfLEqvJ0tR59cNJSPz9WgJVDJ/FBu7REJ
BzqHQhCKVeR7TyG2u3DlmduC1BxKre81ahZ6/LQxsNg2yyKCt/IFbmb5WDGTDlnG9XzfTFLD2oP0
FDOE98xNKjDqI+SkoANuen3EiZ3BLaZ//x6/V9oFeWMc/AU76ycdIRHSHIz7rIIq/+mQM1seHXBY
mISnxOOEq2YaTzfSRqNuu8TJQFJ/AoEDrv8/Y6BYp5t7t5Pv3H0MSrEF8jtBHzgdFKOshsi5zMbc
zIpuBssa35Jz6wmyMwp7Xpxm7LRqGtJBPPOng335F1aJMJB6f8zrObjHNmlLNGl1sdIP28eCNwqf
a0GdSNJaQGKIcTVHoLj5Uo7nlmcFstrodf+3Okur9VSGcs9PRltemTby2A9YIsyXt2MWOkMW11GD
4yzHfpC7GCiqrTlw9caF8kIkGzak3nIAzYKXMmFVj5otOTNsUdF4JnyZzHtCHuZfpP/LPodZWxne
Hyat9jhQL6THH7aq2mTHZnx7oqVB0OA5RpHF6xv5BzwhoQZSGWzaQgQPTV64R6hmFpi4uBA5NZjI
8tjWdWbhpyY+Jzu1jSc4CvEyWXvyr522D7Gv+E0M1Hj3yyE18wDquOumFpsY79VPmaTK137IMOcb
6ojukJMGOcUA3Z7BB5OqX8qffIWvKu0RjmpsUqA2lJOxlAJ0tX2mxFKT94Gxdp6pOm4497pYRSG+
WKci8/b1XVWuIR9nS1p8HZ7CBR0HVRGJEZxZzNokb3Erq7PPp7f3fSK1kHATaWao8Lft0abfxva0
8STCuUkz6kf1sU3HUYB6kgUFwBLB2ocLglcckyvu6oUVKBwGY4PLvxL0rrCQ4Q9Abrx1DW60TbhI
LfoP1cJ+4Qjda0Z/UnxwzEljNnRbgJ8Y2cYkZEaS3hnY8gOgyjUMWZ+nqxqqM2KrmTUR075XEYKm
DFOZeh7dMnUJVOpqXvT1509Dv+HO1I5LhMXJf60OMBVt7/d5STG3PhmmncdLbzAFa5N4xl/rGpYr
6NU4nRvSCG3H5AjiuSJMoU5Lz5O1yx/lovRIO0kKV55R7DQYbeUfAwfh/HYcIPpVDzJDBtA5JPNz
s9ylomWe+PfH/BQUZvJcKubUzC58AGKyqjbjU4uUrt/WJJV97MHcsBJ2/eZ5BgX40QiZpjCDngXB
KAPA8vCa8LyAJcL085zwc5yMhJMEtEdzZbNtIPg5mh/YwThrhcMf6rk53Xrb4Q2866B2ye8Wwyhy
lhw3OKEWHMZuL81YnqZEaBtd6d90yVfIPFojgGHlJkSUVUGBjDscCFN674EbIZHrhyg/6wPNPBG5
v6ujvXtXBhO0qtX4kFSCUWdyMOKudzZrv1GIMazRqzemBeq9P6dioo9f2Pntc6RUVis/9FsFHpuk
jFi2BcMphywqo7YQACeiyFuJcSFY5egOOU6Ln5ohsBqyLJ8pr7kLRTZlgm6Kw+fyj9Ia2eMohPdW
6MUFWci11LYHLkkUvjLhUl7so+Dx4drOdHr2VolL6fMCBEVjiJl8QIIzj4uv00wonEnVh/WrgYcp
vcB3PyGhfbf3xTFLFRNWR8kugH6fPOSen2IumOOfKWQ1E4WJyz852S7iX95NNaYFxjGPaLZ34UtO
9/IhWJzdlAZ3pJtSflwRUjzYFKL+qMdRptr8B6fIS3n43KjGRGi+PqmhvulVCLAqCnuxPm6R5TBq
ib3dkq1Trc++XH7d0NASFg/zUiW+qhZmZUkMCo5BBBjUD9wYkCr+rRKULAlrXzrB8NFRPc95+OXW
JVf2wVeoq49aZivcG6ZAUqm8aHOX1azWRHN+9CANi8Dz5ST89xfzHUq7IGHgR/+SQLTtUZ3nmBqd
NOEBgb8AK895f6sqzvk0WdQv9OlKsIDfcjtS5xFCppqAbhdsUc6KmD0ebkC5oOqwMFlGwQxl+n1y
0ZUZtKzuGv00X/gmtLjkprOnRpurQO+Xl1luJKCEzM+vfEXUIJto2wd0EfF6STuAnW42u3cleqmu
cnHepvNTGZ51sD4w2gvyOWkqa3c7d5jmDmcuAiTH65ugRbuC/HLB6aSj32v/m4rfGViohsNaGycr
yjxkObs7FqQD10LHuuMN06CdcYD0JT2Mezflg5WlOJkzP3AaDzU78WnH+cVpyxK/LWZogiZ/A9am
HIjsgx3e2NHjQ83gNpTPuWEnBJ/dzSPMPnyjjziyiIoPdfByPDUjCRUHN5NmrYXvEPxXBBZ3mukU
MGvypE2wJZkn3/4dYjJAiRIiohv9BGYSKhlAZOnoJcHDSIRi4mHCXKJNiHQOhvOgOiY91re3aIPQ
EPjOtBwEpIgsoARsHvUCCtoiFtN5vthQdPrzpg4FpWOkodzrhUGMyy5FUpVxh9L8kC+5Hz7VwudR
lrRDw7VcMp1xu5ahFXXehHHxat8gLmRlhOlgQ1yF3wnIR0bQVGGGo+v+ZPEJ2dVJr+bkPlJrzI33
rXSXpY1pYsNhsRBeiqIOAbiHednFQqIpGqlNX9HYi+8JYVwxZbgt6lu2Bn13yTK1RGc4TpOF7oEV
YV6paGI5H8iqsHu3gymhYzpAGgaG5C9Lu/BnfeGW0MvuMdLedwcewOnsXRZk8l/XkxuxcqQomeZc
2A1OUkSxFIBZVLVkWvnjRvQp8YEEwJ+7mofzRX3e62eoGJAVy28s6JJ0pKBU/EZay8C6ruK0jV8K
U7NCDEF3cGMwFVeqeMzPgd50XgsbWxDI7+rsAJLUdCaHKCtrqxyYzd300AddhtcNueU2SP1aixg/
LyvRSWWbIhgb24Xw5edCr6NwuQTt2YJixLTrq4taqJbUY6MfrfZ37oxGfbJ5bL0rr2Gc0V8f1jtV
FThAEhMFppAFMdYFULCJFooQevs4NVmGnZhfoA4iSPth14ANZyvQr6eXlf6PTyKRRyl3Bk/vRKl/
cz3JvoZYDQljOoRqdqu1+Y6z5pSdaVkZMumVZeHrYERk1WZ7Nv6r3nyUjSnpy0jBj/0qjeoKYUvn
S/rXKFcXtPPOkbuN7mtp3OFKGbYiX2u8sncLfpJ3DISlk0sQcD2EP0QUO30ZFVokCQubiGOxMv3P
9dx+kFhDVqr6KI51yxRguAY9h6nSKMT25qN2XMwMUyo77gkv3og8UJavIQ8nA2TeS6qI6JminxMP
n8oMDg7D90QBmTiuWlJvz2oS0rrwHWPalMpzmCXUZ1YUQ1CSw+p189+q57oGcAOxp8S6wFINcsA2
rJtUF05Qb+8YtJ/4HndffpFy/NFXucbsML7gIQ/n8yUcLyu58mnTzmWLlckdh7cvOuWm573NEsmi
mDdazyRD+5a+QCmn+skfBdX2Pd5x5gvV1BRvNV/ILWPrvy/TwC2MnM6pX460WRAzyJadQ8wa8AIt
JnNxUMaEHapGw8BzXmI76liLNOtDYJkxslQdoxQj9HtHgEk9NwtCWUfsI/aNvqKPRSITm/sCf3Zk
R78FeFWUZZ5JscFXjjYM15AV+y6XzjeUCOXMU3Kly0KeeSMAHsFysdBCSHPc3TXKjpvmfTklClnG
qC6nUNHoSOeoQyzxFlLAcAE5QUoCAhssFuNGFf2YIE1XQZTkMYm2QfIXj+UULBhHuzZyU5vIxAzE
fPrcWsIDGZD2iAY6ybD/XcJZeJW5ZSCpRei1j0nME/vY9ZXpSRTYsLLqbqfWSrPxRtRKdsdxRcPc
ivPM27hdOwJg7zkWgV5P49DCWKSnvNG4AkgGPDnOmApWiDabwkzJKIer0DBDoX+hBcCCBK+jrRR8
a9gUw43i90l0ji6K+TvhdNjauYLH1d0IlO52unSlW5XVAKaDGM1AVJnBAztTWeklUUtJQCFZri7K
PFi2Hm+fj2YuClpFEZ9cuvVrMe8/IhyOtScEM0X756xaIWonVVNgY2r2LwQeAbeVKFo9UGI8bcFY
MGWOKAkUoRPGgSj2ZGFECi65u9yX4U3mxe7K9+mnZWQ4gjaqI7EV+BjWA3RpcJsHwhfGMA9KYXX8
K46iKsAqRtDebUxF2oFVN+QQl7LgRoXvb2H8FosqruhmbVDeUxOcpOl3wo+1RJCV1oI21uTAwfEo
iH8xN3gtMe1wyXYNSbUXxTG7pvm8wtlteomZcx9FTYcJJ1mmHjlqZZ2VGbSd4CE3IJzrs4xnaFk8
uNkmSZssBmY/u47Xn0FPm8NOnu5mrhzXqZQ/3f4sHTgO1LpnqBkTUK4neDTblcD63JGMh8nMo7kg
bLdLp+g5AS8sNPWtroxMTD7Z+yIjiGQEU8EalIdT8ZvUq6AJussF8EaeKQ9MuWYKZ4zAKBpNAeWo
nUsGSsOa26YDLGMIsVJbd+Xb3yfyXWuncM4LJpIU79yKMJ2CkyOdoIL/70BHDIJTjVkQSOZzP3+J
v+TXUZlZuuZWQpzYbhwQh64Ve65/prZnhIRinC9G3pUYpm251lMSf4oML6P/3UAE5vg9HwoQ7asZ
CBo0bO1s3tzGJR8QlHlqd004nRwVPsDk8ydv1d2YHKkUbjMT/SdMVZv5iV/U7Q2BH8CoxdGRRdb/
11fYMopCcGXS5WshjAQ6JFjsfPunc0DrMq/+1M8RBYYzO54GjEP8CGdXzEPVy5YpVU9gxK2iUAHG
aA2dgmL495ijhnXL7z5UtK1a0YEnesrzC5siSHAZz7KTyiKqb4mDxOC+flBgAwbNfHwNiameP0j+
KJkZG0XitMe+YOSBOlbvMXEnPFkwbSWsI8trg7HoxtGZvr2Q6uoAuyNtSvmhNxK3ydxjobLKzQzY
MaqMGbtP3xPDPFXdvoPWFZZBOH43nQv1HBfovGZxK6rERDkXheLsihcgDgWlzrdo7b6x8ySYvM0z
J2QPHZOnowUYY/5vtsFu3xDmMwcv6dDppt5bTOYfhnT6ENdPyQ4MQqCAN+Ai6V7NRjIqtVpu+Wwy
tq0KXrurhHa3SEhCOLswd9RZzcz4QobIBhODX1moRWXTcutTTvz1PG+gr9wvw7Ae2PmAWWaSux8C
PuNrDs8ouavbCXsoHBoaF7ECw0XrA1GoT0spY+E2J/5X9DYmIPatau/M6bDeBeAy6as/UUG9SgBx
ReZNMZ8nVeFRKRqGJkFTSsHatfWO1T64iSEz6Fv8Xuys+AHagSILzd2vfdyDAUSH5G+I3A/z9/ZZ
xIe5Hn/BbR0jX6LcAjDcTZlinyMS3wzkdJvMzyXKGVJ6/mkkMvgQJaUu5L4nuqn5VONn7cAAzmNE
lAS2AxYfzXu1zbzS1vMavAZ4QOVyGgnHMTKhVp67aOw0466dhh/GkPSZ6qkXnfupD4gzlHca51Yx
VE8eXGbB2YyUeKjDFxLcpf9vpah/vY8zQavX2wMGIxliuduccqZ/bl/7tqnsYaxNkxyfiOXOxOJQ
g/9VZyVcX1ShW3yjJXqBabPN+4ROQnaezXxTGLnAQIlpCBRttnKgDuBHwqInB1SUy7d6aIyskxHE
d4F66J8EH0ZrbhbTKa3m5pQWui1hWT6DOeVxX5IU/Dfbx0Hf2rbS3/N/x8HVJLxWG2GdP/6UszfL
1C7GyGcxnZAAS0zTj6XBxBIRTnqVeDvAmSQAcy0lHHvQUafxZfX928Ur+GSlJMivjsI5eQpwMzCn
fLBwaG1DCTcbYL8KHFMgauI0mnzc3D72xleqEYvWaFq4otPPB79aLjKQbr1+rAf8WCl+GaNt4W27
i5xemv2UrznJdUYidm+M2sNkWZBeehoOe779XI5fIT+5M5TMCroAJNSTP1LOPXlErKArZhJO74BD
sdlngCCeQ79MkZwUhlbDVkbCMZyUTOxT0GWvRPbV5BBmKUiDYQ1BCd99bMnpNV2rFgE7LynkL3eU
upfKTq97XKaqYqt3O1422ITJFvoDGlAyMdb2XC4ol/XNYmlvCbyD+BB/oEgxX4e1BJmNsiQTsVwk
yIWWqmDm841iJo3svij/rQTK+sAkm7ZjxSrqzNiuUCE16HNBYAb5xhvafyVfKHDnmUYDcrT37fnm
WXT4R7JuyN3B8fKHWBU6sRe0eIocYVFcSoRxISWcJ21w18yO6VeLsNajIQS+ggIJ2R3MslQnkCVK
9C+ls83O26QGU1gjP6qg04XAyXG+VFgu+SFWA6i7CrzSAhFaQIxPY4cfXPYd3kuDBSeN+tFRNe1u
0uFnPBgt9AJxIJOYTl1FQxSCVNe/kyhjOZw1rRZOcGFVOsAOz5K0cUyPy4BwoVqESuNgWNlYjGM9
56R9DvtE8aW3ZEgHiD0KUy03CXil/UrHjK5p5Vfn+wlen4LlavAWZ7bYVT8wuNZLg+3WI+Tq+n70
YdhmrRP4kw657OnA5TxvZ9je3hc05zmk73Wd3LS+4mRsp+DCuRwEGaulE56d/QwxeuYlr32XlIIr
uXqUxt+FBNjjQHeQ0z+kKJs5Y2vE1jkB4fteHmoYIrcVrGCK7efUajzy2fpt4/6HwUh8/ET30hko
9KApK1mo4fL6F0YJN2J1e5eoA3sdRskUaewy9bn4MeS1KxKpInCbDNTgEcD1+vfRtfnN3q2Nq6l0
3VN3rs1glh2yf7oo1q/MYoigyxc4JlP53rTY8vHC78qNXlGrZd1lxsQFi6V2Gn5QzN/KWuaZY6iK
UCpgvN4Xn94L+Xgc1X6ayIL74PoQrV1ypP/DTE8801f/2M98MnHE1zWKBFs0ZlVabfXtKNWuTdns
XdvV4BEm2wFxw0EcpLTmLEWSNAr66MZnWR7cF+K4M+NXXH2EJfu/K67LlecCYl9OcboD7lRLMfe9
x0P18aCgMc//BwV1bC8f87Jfq29s9CAKj7eddf510VZq7v5dKP5NTxUFAJBMSRzBl+kKspT1Lqs7
95tHXhWJg0reZr9XoQIlkPOrZ0dsmhv8hyKPAKPHeYaOCRa/SMsHmaneKuzyIum17xEdtzMwsq7R
xpqr83QLEu1sGDXVCsjDcMKgwOaz3x0OZ/tlQQC0HQGCN1WM0B0sv1xQ/6hN8W5qz/zdfv2rQAT4
u4JE7WUHaIU5gIyQjIPeBcBD7MPYL2XFK33onnpp3OooPRfuKTYhtFbdMpnBh15KVKLbZs/wGyS3
CJPEBdGEW8UcwQKGHvUq/hO5dlOMZrA8wI5fu2aqcgCtR8nL7P7NK40kS/SBPLDU9EDCJBzostE+
OOX2OJo7CQ3pgO7GnbLcL710f26bX3+VCGZU42xcdPCpC/VAF4U+jAvD+i9CQgemEZQD09o1Vifi
igScjWRuI5rWkmNOe4j6PjeRea/RmCkW8fSN450X3vF45EvKM0lebBGWWCJwxZzFIw+wSv+6TH0f
gAK17VCL8/TPMShe1MVHzNRGdcOGirqK80uo2Sgo2TCO4LYs8v+WgXQzxggxstIX2Xrk/nl/py36
Mats6OBns51PdlIS5Ugi+7Nvj1CpVrATL0m3iFPzYXLDAXkcYCe3kKYIEvxmP0Y7ZiPyr2yy+JFf
mLSPP6qkYLlkt41srTymcJ48iOrEeN9eM/P4/4RKL3f0OT4gg1hVBi/rttold0ANw9948P4OcuOV
HbzavFXq9cILjb9w+GTgbSUYlhkgPOlCj4q9Khmxlv8sj7uwXH5jlssVdsAWADvnQ9B0iRDs9KhK
ayvojkJe3X410ug510aqI+W6NV/gDzT8ZfqHOupkQKoSOOZWra2Xc9XCl+ffZL4CITeiNV2kyK37
JkvNgyjhvneD3Zp5TlxxYRE0WKEAuy5zWNX1YOFGOdUVPE0Tw/6vXGoa+CEIQ1/oNVHszFVCiNXy
faTNx36uEzealhVCaQoiB2wHIiZ6XWpemQ7Dm7lfdk7Wv5xbkPqYlLCkvNLcgCDN+4h2qLY5VI8+
vlsjyMcBLs5CistJpvTM2c5yMNcy4k2WT0ukmGuENDP2v7hHlQXZl8p92nJJ67gx/Na0PVOLwhDA
OBnEAgbNExqeJsbpC5XmHnMpY3J8xs8RrFA0SAHltHuNCZE0dtIQfe9Q67K3WBp6IJxNtNS0LVw5
OuuNxV5y+uZa1SaSqdARUIZhpauzPLCNa2wQzRWMo5PqIumGwcbsW3ff414HRkGzB7cNHMW1AQoW
eXJwWdUY4ek2SkPpb1roi9/HlGLf/ChYbvUlTTopFPZSQSXDsb/0fsFdPh1o9i56wcQh361JGSy+
CKQgSKDfQ/SLIHcMBHtgIAczdtPpgb7A1PhZxdL8zJGdEdROWz6eQ/av0F0Mmech1UFws0zQ1qtK
7yagAR1ElJ6lCovj3XpDeJlUvQh4vZxlTDW9zIt5XMWQn1FTXwPRnnakKWIwViMgbYWmeTYGrR3q
yqboGBgBaGEKf9BQgP0gOCxA3SSLiwyIdAN/LpFk3NZy8XyLGlwHSguYRgJyG05bNMA+ItaG4Ra0
r/QEuT5m5P5dw8BfxUd+csH2i8ElADVtACxX6Nn+LIrH9/mpf4ZWp7aAOKd9uZpf5fVkuRXQdVh4
aa7Z+/lIIejornbe66yQwBsBmaO2RSw1Ix3vNcgzdrEc+rXz7aogmFJ6aWGZw2d6WgDimBI+TDiA
561fI15zKN0JD/j1nQ8Rl/qOdEBJAJ0MCaXY4UnW0WX68fyRYgwoIaIDRs/4EIlhAvCKg+ucq7wp
kC1xxWqMaVPhM0tmYTTcHAEZkPncQgZxPKif89wqHR+zoQRUpK6JAOfsSrZ3moOq2GuXgLS58k3O
p7HY2xGGAhI0lYyF4jE+b9vCSf7oYwJ9AK5Mddw5nohx++/+dN2HE0+loHwx2mU6twdG1njq0jNo
JQ7i+AZHKKd/pMcWZn30wkPNv5cP1+nOtfhSn9B/uk7YMdiTOrH+bv0DRrr31gNzV4lr3fMVBcm6
ggCEz/FL0cRtxClBKR2Tw99FBmYYHOJqKjyDDd54ombnaFdkE05Naxj/+L/KPjAHnkgdibeFVGju
sTWwHFJzn3J4mr/Nti8TlldGp8vVjgU6kq3qiko98lVWF+WXsXMfATFPH2zuj/ZQSw6IK6e4yQak
kkVgUyzrLJEJfhwJRC+AZqCGlIyTQFQ0winpSu7fpMlit0Xr2w/1DfFsGRPr0DkXJuYNaX+XYA3E
5XU53v8eoeMnAUFP25YZn11oosVMnt/Rt9UZawgH/N4TFV3EY7kqspQaU/VtjOP+kFfk+hSwofOZ
5QVzydywB07R2rXoknF+6YANlPVVAKHCNoNL3wlVMnBny0MbqaAwnx6fl5qUgHX0aA7itOr/AhOS
mr/4R11sP8lLW2LqnhXWrkLHRglrQHg9W693fvd10EeEsMdEK239cYpwRKhUipVz3YPuM0neRC5r
eZIVp1pVNQ+/tUxtpsft32Cd6ZZyPCK6YxnyoB/Mu6A7GXLvJEczfBLNvw+cZtwctY/+ic4M1e8F
mVEZAo0kelibLe50JfmQMQXYRVm23yVaIIO4DwcsJNJ51Z+cmH0IPcme+VyqgzwbmzP9U+hy6UaL
FDk6yqBtrFEfkeFiRhfdCiaX4s3JeA1EYTgcF9lqPBCaQ1QpZPNZlhx5B8Btq+X6oEKg+Hz/+int
zZ5fK8K1Mv4D7ee9P8MjQOnvoZ9w+8EvImMK+LgD8SlNze8HQwBYu8HMjt9yqyA1Iy53tC9moZ4O
B6ez4wJMFJrRTN4pDun4FWxyF88YnJ6pm2SSMOL12epBN1mruaMsYM67kCLBFp7VMExkAFarpi1a
B4zDlMLML+1YzbqSVmPU58v3M1KlbETph9IqKR6xLJcmD98bryq+Wf/EmZkiTJRUM/8BrgTj92Wr
JcQjFRcD2Fxq+dcsqhr6JkoJV+wsmybs4Ehxn8QN9bCipjBURZk25ytTxHsgdOpNkE9FsZpo4JWk
5wHfl/WyasN6E8Wsn9WCprVmtUt97rRadzbPpw4QQC79+mURd1Vg0M2BtqB9pyKXP9+oidGqcLK6
wNu2ZK5Rf6wO3risUV8tZw11qrpgg7nFB158tbBBNvL7VfoC1a81wTdISquVw9JKWjITjCdMOUal
O+eUn/oPW2xmfpFQuoNWgPHOGsoVNJ3YD4jEahXKpmZJdjyTOa2HyWt1ZvWh5aaDXwEp/fgRHlmm
79P6jdfTbfwb4YVBxCsxRfLHX+ZNsaRyOgyojHyJIO5bG9Mn8K4qhWE5nR+LVKADxELPQszmtiSJ
seKoL5eCL1hjJ2ya1PW3OUz1hYFH+TzqcFzP4koNp2sx/GmcCn8Mp5ZPrCB1aaMjGQJpI9KmXeg0
S6tWT8L9T6rVweBE0G/fsyK29JwGqY4/fXkpkutEyzrRTBhKlykSDcLiQs9VcwuZLkb2FW40iusF
o66vDZgKxxiINfR5V7HzIMUxiG/F+C26RCM7pk0NLqxdwXinPgRaUxOXNbrmRunWuT1is5rDI9CW
NMp8xzhX0Mde+JTJdCOtSv+1OEjxvx4HCD9Qlw5zh0h3Efklisrm9zGRZ8WMkMFHXf9ZfCs8kv+5
Bygo8hnYB7ZXvefw6Xxelsj9iXJXf5XBfE8UwpgqubryfB34wGVmLwraeCi1v3jBC3Fv8N9XvxVQ
zCQFjJAC9Y82mxRBibOARvO6JaKdPpnWyGQSVNcbMuU9jZcFFGAgZoSkHw/BygYVfAPHZfiUa1xX
7PrHx1tM+ESNB31GZaY86SmW4RqmQRGxH+Mqyva7HzB+SsR9/qXcf5NfowWSKVhc7dUrB1mmgGoK
Q3Oik6zLZARbkmFLjmjk9P7j5iZhmWirBmTbq9mGb86dGEEqwGyFsOXeF5LAZxH7hSD6fHxQtyBJ
7fYitepP0B1qGv7svcZ9U3hgBKDO6yAuxZ/q/+twavqjBjgLxhKjJ1cCHpOr8gLvoSSm/Rd2SxKG
VGheXIRAYWfs/cPdTb6K3Whc98J6g8gNNXBphsAoY5yqgjveZJwv3kzk/lP4vfv7OwoIB7WiaJK5
a3To57Z0NAHaAyZiA1rUHhycHQK6mC/Tj0g4ErfOFqmBjQ2R6+sNM0HuZjZc7Y7JXkH7Yux5aGjG
BOgGxt6Xvy0Yv8G6lbFCakvn1E4v30L+ThQv1x7iL5Tqm1xEPQ0HpBoRXSj1JR6ncyrpSre0z5Mw
Jy1KNnblN0nonQSc+PXSIMmEfQoK8PY3t6skmpOcAd3kSaxXQl2eo4QWVx2rQAZZrKuBTWEVyC6b
gp8Dr80qmLRUXPJ1HZ5OjmnFTXkCbCbLuqheXLKx/VxTttNtXcBhoqfNZM4rz6hlwPrXDe3Y9ml2
7pGsHtb4AZYzJI48lH+L4XIloZj61zR7im9nIknmofNz24NnMKuypkLLSpdjZuLpMKcZQ7Z0Uv5b
K8Q+ZHL6PjOCURusEzIccjWwNkQqBFSZX+RWs6PQ4dRPNFyPTgG0fRKrSOysgiucyifM3+9Ct9Ea
w443015QZiBrLxYYLAVIMsjfUTeRqEWhEcmoMNG/vCaRs2YwtUgTSGbcUS5xzwRvYJaA5stjuQ61
czUqx3dxIq5ZaZ48bm2SyDKQ2hW4Ydnx/N8/kvcP/wTCYsV7mDKeqjEZy9b53iSsICSJ95QrTfxL
qFHIEtKEnh9Wq+s1WAmJyOcL7HB8jmm2K/uCwgxESV+r4SqrJKOrlRw/iDPQi4XXtSpquFHobnOP
r4aMtHOATjbRVXBQ/OcqmwzHujaEg0tAzdT5yRg98DlkUsXWzuTqP7x3qpgZafgxJmAJbS9I1dcH
GX+C1KB9mftTrUnNYBVc4UH94rNywj2ABocO9l7ORzqTcvgHSG4rSkabwCKjB1VvHXIA8iqoa6mD
HevZuvNDRCG5J7t/fkNEvIiPQtGz7zQxVOuAtI/XzTMNW5UgTY6884S2geJG0hNayu3s8oFCygyj
onoB3S0plEOCm7+F9qGYd4XnTb6DhOd4K1LQgPY3RJUXZ1LvC9cAdZKPPa9XTITtFVLzwxqGFDWg
uNVrUKkj/4QKKOYyAMXXnwkEBPEYez4g2CWxEmfU6hedmRa/cvECZK5ipdaoLO3w3gyU1arG6Ka/
y7TVB/YTe60igkOg0n1rJcdCpZs1wotFH3ZO7gRvGgAkGYlD1OD8KBQ/KD/8ftA4DkRsfIEfcyQE
hS0Shw1RImDsPF7cSJ5OPkjKItxXGuLkl8VvYE4S/Iau1zoldf3x9OSDHpB3et/HyIzY88KhnqXL
qn6/cPjr5VRvz/K5Dl8SI2LHq9LiAw34vdq2B1MDlpxIVtW1YryeT+SDkbbWm2QVqRugzms8Bd8Y
wXVj/4o32ZUg8f/iPnl+5GZsHs9WeeJG6vOu0NGk6JGmIVfnRRvWHgPVWKSLeqknKVZkJbTT/ZbK
V99OITJWgOzYED+Tblzv4PifR6ITuUKAPCNNSKA0ajLONBJYkMmBr+cAmWI+vyTnzby36z2UF4bs
/p70MU7XWAmtlKBgP4DIbQ0Wecce0vdsWjgq8sGIbqGamTjKZvebpncpIg7ofmLQL0Oh0YzTt5vj
bNu2g7eYJKTrg+u+7ynh1KpnC70CoLhraZ498zrYxAJIRAYa7iLOcO0J5vra+oSIj1abgjAwJ1e9
cRuXAVJVVNxD7futO9Gd08gmayJriKk6MnLM3fmBlM/zcu+KruH4g8YCxWUGJqLUz0cY83KGdpiR
B4lT4qqk5gvHIwb+TwKhOtC1a4Mqz9kYS16cbjEGVd/ywG5DYbmuEEzmUiv8Nj85dIAOOCp2LO0v
iyt4xDfuzp5dUyRovhGGr15Sbwqjnu6kXxdAuSck4yaR95Ivj1yKEyjbI+TQXP1c/2A2yaTx53Zq
5r1ZmpWjq7vQQmjFQm5MLWAdtD4jPoasmc2ZebXi/DNSLNPDWP5W3SSnSu4RMt8i6Dk51Ia6DPiU
kveBWgmibVrvArykazZTCM+0KQ55KILsQTsTO12ST0BoI86KgcCVZKjb+KxXNFPot3J7/E4xB10H
MuhwatTtdDPB6CSheLSQES9A8/cyersaoTFQj7ZxR8QBw5k4hUnuHuQcZ+FhGzOt6/LKXPGTKkWA
//RCLsbGi83D4vr5JwSxc1gsNtJWzGAG8zn0HBFsGHGmgyYIn22d+uJdm49us9u5APLRKQ6FRozZ
fMPPD/LLHnmdDY7mm8Z7sfqs8GLlaWtJkxC4ODJ5bTee0pAxGAj+5BcOxPZO97bV4mgW2T8Nt9yi
L9uI34XKBlz5YPqwprbu3Ubh7XueRQbN5VTtVQ3/1qNkwH24B2Pzf75C9qIuKy4E+aT+xex3iglU
Q6IUyG7siGPu1FbQv0l4P/xxqYWO1qD1g0cpITj2BPWFjL2XUnMNBwSmTUhlmZperTVecRHDJ1CL
m7BV9TCoWOY5Q6WKjA2bGGRhP5Vv0l/dqG/kVBuMqvn42Bjzx445c2YfJuFxa98eIaaax7nz0y9z
mPxSxs433jtgxmukQuBZx2XP4a7ziSPdbXaDJp0MYPlF98nuD9H8QP8GHRYo1utDsX7A++QwE0fr
vWUZtermOj+ZO3HB6npOkjAa9pynNa9c/mqoEKvL1H+avb+M2P2VHRAR4BKGxmPUz54ltCodnD9h
NajiYHJXAfeIS2+HubwwNKdAuZ0SqzFdFs5SiID4T/zHqHIJULX2CIK5jYcpszkHrz+OOpwwU8/9
esHf9ROOLyr74XJZ+IZjVa0OGWMNAMwgVNznG17SnL2h+d56czrT7Zr6ROa4QsXatJZn8gZ4GHyB
L2tpeG7BBTcJJYLlZEi/fchu5BQNLGmG4rXkReY6QlORt3M1jKeFK2tQJjG/jdTgWl4SWTWp7Bn3
ByQmZ5OwE5jyfQilVZO5XP1bjIZbzRSgsHMF9cntA/wPwVeUaKh/ffM7txqia2hk8Y2cG7gaj7W3
0D/eSp2uBHpzpeeM3sNBzELiYdBCELMgF3NNyxLbp3l+ji/vXTtGqkqF+uWK8cdfTb/QnmWSLzjM
aG06TLPqtoXmKp42s1NxMg/XNjc0C2LgsvpOnC/GK+vMqLbxGmdFfn2I9ELFamfTYqw1VwhrUlfG
9TtEw5fDE5DI730WDWQtzYtDfNX5jxE5i98wGJxFaUXn0fU4p20p3h8I79yrny7gVKw5DCgjfglm
DTp+6c43uhupMXVMEV8SSiKdsaTuuZrmXwnstKFwMjo+KW1/0w3Y2Pg2nSQIpZQ6VWEOQlAP0HfZ
/TDji/TLcY2+WKnI9+4ckKd2kwgVFtvtu53+xByLWIwdE8+XnlriZ00KjvDgUi81pZHJfJi0S3sF
LUlWtuCWP0kXyJy0lRtw1VAUQSa8advdGsRlKznyNJnmMwxWl+x2+LYAwLq5UsWhMulNoA9TfmAP
8I+OCh5S4Bro7XlEZNZ3oyW2vUR1PIb1A8ZcnEWdZVqm2AZwgcp8Vn1FHCjhi6QBMvy0t/6tGkUG
8YV1jObmtDv4WZ26EST5ghfiz26JGNh7e2Zc6io08CeB4+bql1K0cahawFruTooaFTyn+VR8T61+
2N01VngoHbQeGotz11OYMLCh4en3G2YOs0OqWOVv7MjydjFiWpz6LiUK17D3X1DGZzw0ilxgE7DS
z6iqoABjLa4ga0E7x64Z74M069C2C4or2LoE41i6yn+Dz7R8zzXRMFeBbBzk7h+Rp+g7kmcqwu1H
SMRMl0K1MXpB1R3k5PBozwwGjfuQV8kRPZtSRxISY88VHI3rtNTAJnENjwxCOYGrcRi+QfuR4lUA
K7R+o+OtdgfPi3K9sKMBHHjsF2nR8J+uhmWkeoxELpvt9k+B0XRq0J2+uJU+d4NobcGGvuKdWUdA
Yy0Xix+78Z55MwLmVrhopTdf4dq+2foqhv0RnZ6hilbIQJQq3ih1Dapn4BA3PA+7t0kzg4WtyYjp
ZK6A6RtzPgddgAc2VJWqYcMVEeqwki8BS6e9g1sHvOSzGTSVcIwnjDJcXTUnqAc4hxhYrWkldHbe
m0fRMRwY7KlTk+erFKVfVFAslFYM7HD7fq7ItJR7FiRpKJbiIdoecQx7fYShU2dOrWIdDbyR5gT5
ZhqXQA5s+YkaxvhpVJmdzlwdA6oZC/xPHTpZ9wVVnBMudU6g8juVErN0X8gwdQ8To8rIO1bSKKVJ
P1iCfVnTXBjbOgchlu2Za093MUK9Xp0euES0tWbWjgALljkkIHslV7ZHwi8VNzZGq7rGx3sYQCIH
dumbP0Y9UXJth612CKJPjneR86RlGDvcyUrrcaxdPTqL6SlcDK+X7KAWjzSGUjuPlgGUKcETbjGf
r8clubB70BX5CcoTMIXBfYFVQMFfNYwS3LNyAt6mMln673kx/gUewGHDu4xktTGjZ7JrBC32xaEY
WexvpwXWlaNRRVMSghplPdCsfmxd5irZ8BfiyDh6QdiQE1zaDEx09ofSW4GdYsJfriygMxiTdzzZ
l/ruJP6BBj19QT6WfSaA11w/2s7ik/MccW/ISQZ5XNfnZxv5OFN6vsiwt/SFfIQIsXItF41bAKFK
6ODkOt+ddbDGLFl/MeZl21lG0lZPJCOPI+9+ho97dQ8OJzGd+xLVZpM/klmB/t7X424BhttHUSiG
S3FowQz8JZdcQ610FrU6IyeVUfAl6VH9RLhe6aLW6LOEHQEKmkUGDUF5+NEPhekPkzAKXWA8nQ+6
bSSnksMquAggON3uxQGTscRhrZHHMiw8cJDM6qrqIKSKZtZETSesMvhzrQIAMu8sbLyPn014/W3h
ViPaDoCzZLlV7v9nxZuYoNodtuuVr/A7rYYSiP3P8PhrXc+qjLW3dOiouxSfmXpc1/w6QQPZ+8yq
h1V1F6duCCsHQ73ILTvQ/QpQcx90IGJCizEQ2VdC1CVl2YBqh1mDY3vgUO0PovDVRJD6M1KZSBdW
yhP+0uO0m93bEcfyug8aFMuIgu8Ewc4Pf9THDHSMEMRXLH1d2yaX8bg3Kjb3ugb6kgxNkQPPDWuq
3+2liy4ltGh8QTzsTT4iuswKC4khM+2cnvAxxLHq5XFLzYP6dnv2mcgYy41A1WYN+loqunoAr7pH
voUui4pyeao7I+pddJ8r1LmEWdAM7tTabLhiXm96twvlMzllD77pfWjKu1WoFVhIfyf2nUHu7p6c
274BblXxi4oWzjZ2qDnTNXBlVeaXSvN0tQPxecjjTQTYND4cqxIUeumYXE+x7Rftps3VYufrRR8+
PXOL+rInH8GMlKVxnBZo3u5dBKdOADwWOWAI6wrsin10op+wgtG0jMiBsWYVg+rGJK19vXE1u35m
oY5MmqDIG/liR9OZVVW3ouoplpawsf6k5RzPGXvwV0wPkc2WK3YwkwHt1P8JkAXE0oYL77cEjJLw
Sl6VlhxmI3fm2eBF6ybWxapTs17kuLDqFcBalb8vAedSIah6ymH0sxNm4ECTWPjlxejJaZRfY6bE
d0+u23Q/1vyvxX/QM7xJSzmvmV+ZO9URtastJfHStuJezjHvfziw4iH/Cx7SyuKSDl374B1EIXN1
RmSkBsgVOnVeKorVsJbxompEiM3wD9K3tBznhmditxZltqAz8ljZ+bmfvDCtEF/jgdkdSSph4SDc
5sfpaknneyZ5p5Z4KYa8fkwKBH5mth1q0UmDu+IHd8YUY50T6W93OeBLMxoqwB7b6DD0hR7+nP9a
QMkACodjDfTcDUF+TxJFGNmEVlw5l66NYv1qFcCkMfT2Tupo/JqOMaLNymEsYRoa7X6oSA9VQQey
7uwQroaUmXexNI2o1sm8nQV4pWKzXhVok3yLgG/uxqz2d3VajV3sUoZ32arxq7I6zMvVQz0fXvAK
3UkQ5o0btmv6pUDTr2kGbE89pP/NwfpPasbrJefMmqL0h5bA1XvCmZL4+yivbaOcNQLIYh8gObr3
qB37dH3K6mNHgqlZGiono6/XBcwajcEGl4i9F3uNFmxCXu1pmpX6xJFEf15jhcdrJVKEkSZRRJDk
krJda4ea+54KpfBQAKtE4bMEGzxfumGJN7szYc6RO1YgJGg8RBub3rrqkSYtD/Z7F52hEHdRn5Df
Ai1vIhxD6BQusDZDxbZkWgCA/OPhHIRFPzgC21uViOKnQ5XC3epGpmC0CP6UBHrlfwvfNhuhfMb7
cE0icGUpZUMoCIMrCt6ynQLf+k4/RfdPTD7tRpzI4zzpIG5bFYNk3BgrQZ/fDQVRhD+vuZisC1k6
jGZPTilZPj4RbbscDjPdFgeSVkvQneRPpINwJV1kBGPPXzhK9yZmOQzgB51cyHR2mcZGTFAPyhIg
ctapuD1jXY0cqRM6T1bL9KwfGuYah8OtcIoOTt1G3fADszX5bNuYkd08HsZ0W0bnPKdr2d7NbT2t
k1AU4/EMgmOhaLVbgN4kC9mrU6TMh9VcYkf+5LAzf/mCdOdHkSWdfrRIloSxvUVSjutIW6N6UebZ
s4+gj30jV85+erh2GtofvixEwKNrbDmXSF8xyzGd6MxfBqd1o8BiZCvcYdLZk58Qu1cDmRM/Pqr1
5x7SAqTdBbzibQeRD5HBQP1rCOOB3inGaLd9joC4nAJoKkCnBxFX9i1RlREHG9t/bPTzZci/EQsM
ezXjBznL9tKtNpFIk79ndKw13Oq4rgZWPlOKpHf/aGlFZQHwOUuVzVgLqZM80VTk/OFGsAW7nKcy
AJDbO/AjJm+ExmwutUh/yHWAKV5eUtS61kKIR3K2zttnFIWz+8TFNHLtCGesEZ+yIjOgfOAQ1T9H
DjkEmaOynGIexLYFii9XIyQTYwmz3niPk4Sj93em6ubWBafceY5gSnvHmW8e53JK423X2fjJUb66
o62jLbSIsmTcbpWcR9shJyCYOK4xGg8sh6W3S6qKbt7EiAXZDStg5YICiFefUpgCsEZB3bjx5Mxk
NwYwDxbNNmJFKL0IAkIUBA7pMjh6LLi7wDSAGqOhbwgdnkvvsuKPcJ8W+GJ6jllKxxXUvMkDAWHq
3Nuuedaq/YbcyU30hJSjgP5cQuNiT2ghBKTrOX+5SmgmC6S6EbyyE3ngTT8sjs87Hoy/URVbza02
ODtPWXscEkG5tmSaxilx75KMzq7/n8In9aUEK/p69BK9LYMskOpDvI4e/ZY3HYicstQr0nEsNcGW
c0mCOCpF86mQTbQZsuPIfPKssanBjK6diYAqlbSM5UuShjQyN4vAlyl/EiO4ooL7UbHIE9bGBYkU
XYj/4Dw/mikBusaAEUa/6v8Gn8QxwDtbi3Nx8wjzO/b2qGay48Uz2MWW+l39AQ/8yb9WqQXruhTn
O68CrzaSwYa2rKg/qx1YmFciPMuSG6vHB4QbqXi7nS0+PHGAvdFexh/zTBFa9jmcnJDIVa+thazc
XKuiS5JUtCuBoEVRb9z6y+meDLPyg9ilmvBRpQHa8z2A9pEGEFQodboYyw75fkhKtzvEbU7H7hkz
RS5T8aC7qIR3xVTRRbNMsSbPhcZyX6Da/VoZVDfesNWpGuEiUUOYoc84xhC5cBMK4Lb7yWKtdpzO
eVyUnDfC3n4WgRj8V5hkzE9eoXMhNpcYzbIPeOMy/DTXctiLCkU0SsZnqCF2I/15u0tnfm+BK7Rh
DJfgk+H3stJ67ucxrxm/vW+GFeqSB+vLb9NVtrzlgNk1g1O4cFw29qRFMQ5CS87dWtXRSXkxT9m3
gfEAG8k7NbhFblbl7foHGBmpPdFnH+6wLFL1juOum4isbVhocHCKhR4ClhARZmes1Bk8iPCkgajJ
FXc9Fa9+Pi6It4zAeBXqT86k5uL/gViLRsGlSm496VmVpu0XT7dN8uVOFbgzMn2YQRnmL1CrRASX
zbsBajYZTe7i76nib2ComOuSSl+DW8JuD4a6dXf4NsM7IUjhtFO46+9UJpgL/OZ6w/oElHXoS9Bu
gILjPnrLQSsDh67r+af/4V41eXIJusNjI21G7utOrwtcYyK552E10qPII77PiTqOu+WtSGS7ttBu
CkzRVSzPeTLnB/ZjvNBQrneacxkbKdAyH5PtX9RpHuIzrvF7vpuoqTLdj8THx9msb46vP45VFiIV
4CL3ZGXp1zyyXHJzSej3OD2KiIv6SjXj1z8rGH2Pz7yPY0qJ/A7rqzvZWnk3X2MvwIrS5dy3ZUZK
vshQMvoHuih2cj/m5Cpf2jU8Sw4C0bhaqiIStMtAYRD/x87OIAvxhapFv7UkE1pdoJ55dVPKrZna
iG0DCaLleNPTIYHpcc3BVA9ZXUzi19YWvXERivK9S5BoNxQOSZxek4aKPRWxochAUFvtzSWwc4+L
ulNsCEig2fI86O0zbkqf5fbBO1HrEKXwEHbBS2PcZuBXo7zBnU8r21XP0JxVgoFXYUac0U7adZ4z
s7xw5lTUQdEXqeQUiCM6ftKlWIaPd/2grQZOqbbKarL7zYutr9b3PomRWDT3/QL0mQz/9LxdFvdY
dDxju6D7se9jeWGu7+Xqg1+1AjVYxUR58P217ftic2z03s2A/0asnv9sMaLSPA3wo8aKoJB/3d61
8EtvRxuQnloLQdVf1neI1SYhh2qiqusu5A7zAkA6GaxyBq4fZY2yvJ9v+N5TrZSsGGExvi/ehRuc
9HhNhLo19hJdB7lIWGcFoyOsgEyJ6zdiFyRk0a4hoYco14vvllWfzxTndOXhV8Zd6C6iufTXVpe9
cx1iPWsmJq6ubqewVwzqSQQxGUWbT16htu5jM5IQB6Kp0XlRUg8Gud17MUZTnZZycsVc53fM1jBA
zTNrmjGvaNoK8vn/RJMldkhIpBCroDQx5xpFGw5DNNTklkvm/w7ghpNQ+1cr9LR+yZ0CT3S1GDa2
itgQPbzKbrzcChXOIE/bVXmMO2IotYA9k9RIT64bUABawHf01PBloALAy14Vd83RPufDOjmVTxZb
mOC83gcOgcy+Xdcvwg6o/OlN4Ten53ufxHWfvVzKZ1P0WbqgiUsF3skNUgSv1/4DBn5U7NTkEJa7
ZfaWl+tvYFtvClHN1K6xzkZkw23315Dg3Qu3vc6UoZNTTVPDuKxYOCSHw96lgzHWCVgWU87TExqv
EPwuNx8UelRRXcvPpvnQlBtS7RQxl4QPKiRCwEqsl7QSS5rO2npI+1qUjs2jRztdT0FPLoYT+NJ2
5h1YAhAZCxYpeQoY83+hI3Lqptyt1zsyNBhwx8gjEvgFh3rHk0OCaL9vQfMh+2TrrnxYXPvlPbc5
7FoW9NeEnLyKTDWAO7IqL34SEGUC8X/UEKAm27I0spy6vjbZxuwkfcoiqWBzSEc4qqcvF+EtJQtn
1THqnZzdTSYzIWs7kmvbDOVu2dxOmEszipe22rO0GmSwNyBEwPSHgNZNCoqzb7fVzfmkL7Hbz9FX
7FP0pjUQl9rglchp0AgDZG/2T5YVYNZ/7L1nhIcm8vUsJbCP0nJptemcej/NN6NDiWTFKU6ERImH
miFHZWmRWXZKTN1vlS+RBK0bLWDo1PAmhutUGyX+tif9Y3EON8gpySqENsbTM6Hr8yTUBhj5k/KC
N7fazyZmIi+3RKtzw/aOjkGWTm6gTi9nueYWLkMYHChp6PgArmXgT87ty2KIIxoyV74FGLLkArqw
R3mqNoVB/ix1wm6YCZq3Ti+nN7BrMhRvUpTgIdCUxE8VieQOgN5aHuZ2foAeb3ziOdHLPArdbyyh
BNZ99JJvqISe5GAMVBF3S1rlefCDZHUh8M4UKZF/uEBZeyqzXKeFW83vv708pRUo99VLiB/wxx5t
NdM/s9MwbvLuL84Cr44UrmdBu99QNAbGtRc7EAVzB4jfD4txuRxJGObnEPYQGzZGsV4+zJLXaYrX
yUzDRMWpvxOPdYE9DlU845gtSlArWKXwVeUgsBS1eEx2Drm7663mtTp96sqBVyQ8El6L8deIBQuZ
GNBUkTxTnAaotCDkKDso+RrQEvL+7p2Fr2lQh3T+7B1HKo6tcZUD8hvLZGH9TqDlVDIhn1srROys
YpLn/pj0HfxtmcO6b/9YP3h6gyxOouD728O/Rv7s8nDKplbCVr/mkQwFpYHa73YcfYKyYZYLo0aM
Bibf2j0yXRvBzpmjEBNneecMgHA4IY5RfznxTouGdqHiVwM8wOCz9ILEoxH1wdrTy9uLuGD/Xr3Q
/YBWNKh9wWFW0uY0N/KOviO9b6+jKRT7Af5VWdIM+BAcI2OvYPTQ9X/DjAx9RbHj41ywfyiiDyfN
pA/XCe+JtIZwjjSCtase6M1lSLAAB29mj3Cl2CR4W44BinJbOU3fsR+bJHYX5Dmpka/4ykUZ2Kcu
Y7X48IVRSZy7fx0f0jIzLP9gPCmt6wqddsXvTKCYIsQZ1dC5Wa/e+/ix1yJ5VxcqRhCPnhfbjeGn
c4tqVbsrb5saRTcs5Tg36NaKhTejmVyuDDwLdA0DeIX6UoSeDZyFJvrKvUpuAGDaiBcbm9X9tJbS
hTbWWxap5t4+XeI44H52pxX2BlvfY3hHElUasQ1HrfYQb4buua5uNurGcPOIiP8/h0/Bw39ZNDVs
w99mT5Lfv0BVh03/kVjUCReGbqyPVuZgh5Rg0quWTOgA0UWOPgCqbyH8wAhp6jWJZj14PJYDo2wV
2mZ8BSqR7Uq9lQpF2gZke/+XBKig5VFkVd1CQJBbfYeVg3gloKhJASGzZ3R2c7GOt4hmiDIuCALe
5eFELWnaMbXhMngXbxJ0r3I91d+tmp+ldWXhQm8ynOkXWmKpYjSLySXnSWRhE9qX55Oafk11Yx+x
+4JXWmlULFsj5sxIbunSnx4NK8EbnthFc3LwsK2MCKm/xhBEAPlJPQLTZslaZ1uYRyYnFC6zZY5e
tGMbRy6ohO6D5m994x4fMKaaJW0Ih8hTFB4oRmIQ7u96ktncgQVY/pdcj5rjsyn5S6l7cNEdssir
9PyCML9I3A33LsK5DfZjx47hZvllMLOzoX0ve/gQ5yA+xoUidlrc9gpVWff3i0z0cZxzxX9rHoWR
rPbJ2qP74RLZLcL8XOKjVN/6WdaqJdioH9/toLp5M9Zw8MwmRYGW7P8wPDVKRDrlX4d5WW8ZDzok
l7YAyf+nNqw0/o3Hdm+cBgm7tzfxOEbe8HwPGGpreja+3LJx1dQ9IK4UA+Vq7n6WEa3d6xpz3zFY
NXXGXhIGf5upZU8cCKqWp4or73kVx2Oo5Jg8G50mS9LKEjpLvIAB4P9zDoo5A8euJ592PObSBxNW
l8/xjPA8EXx27oLJAHB51k8odmqGToNnSB0KLUDeFk6ShhrRi1dlM6FA2fiTAebKIaWytDMiejfg
y4AS1HZ/tiqlLTiTAmXIHso9Fd4BmMbMnWrKcknteP+Ym5kzO4vujNcdL8QVLrRj89iCYJc1ApHk
mhq+1Ftgn+K+Np23+N8rWx1B2riRa4hzqwdO3bH3SLULzIaMIPM9uJLfq36u3RhhyTn9VgJRTWCx
CYOPvUj4yShm5MftVBG5ty6khsQBxSAGJUHD2iWqUUGmqo4KqDj+4srvy7a0HKO2fBm2NVmLurYw
uVAseHaSPX3htNlMktZ8DKwx9rRoSFIOWv9rOiVzFFlCg3p2bNnFxzAmhVQTDmF3xoScL/Z36GRA
oONunxHUugislISr9SovTfmVSCoj+uSFx1IS7tTVcwAc8WHJ1omSAaGbZle76Y/L4gcnRB0OWmFX
FlYicJysbfyPOQ7VdQkK5EFyN2aAFlXKI9w27WqkAQXaZwsC8eee3meZaWXpbGEoCYBZuM8liiET
ygJoLmvt/U5KEkf48zxYunQHoM/tsl2hXwMRs8RfXOuTmoeUBxLqLBzsZwyjGzoGj0yGUolptLX9
45HCemWATAmEmgLqo3HSRBKbVeWLbz/8gbGGhBo6ZHPgxkqtQ4+/c5D35vU5iiitNax3RSaHVLiy
nHa7Q1GifAGZYYI0TSaOxvZxYTkvm/2vMaQkIAHtpAW86k2Yf3WEULq9fubiG6y5vpImgqTYLOn4
Xro7/DyYsbVXHNMT2949fPeXnaYHDJp/N/+tqlb6krx1u82VV9LCYHZubQgSWGAOIPhARzDcHDZ3
nDtckypGO1FKF3QcS2XawPV8FS4SwPa+0BO8BM9htHg99iFQhw3emFRmVYjjvb2oriyIa5xCzK8R
3Yp8z13K1uRc1eb/QdYLWQWmb4bMN12DlazXbJE1+CaG9+bnxI8OktioPhF7jgY+9Qz14K+38fQn
IwM5eKcc7GuWWhQ0Bh4SunmADQl5YY1mK9q51VcdxDoSvs1WuDA/tyog9qMJKsWKRghC+ZnHji1R
sfxWQIPR7dob+P6Tu2OA0s1/F/xe+Qr9BQkEcPpuOS9wk0Ksfq5mm8xwh8Z2rvFtaA5nvAq5B1S0
fdS0gJmv/SMlFB6XY8E80zQjeK2HHvHnU8iMMP42lP2n6gdtbSxS/q/LbmMtVM/cUIR7SrdVjrlq
nKWaBt+a9IYCb6V+vB36m8Cnf+uUfNbODdFjFd3MLm6gv7oFs/ivjHUz1dNu1WV61ANSZ2oOATTK
UCb9PCRGbn1ufuJwUE0kNSRFDm1+VNFwOY8+EOliVvwwZr9gt+dVvqQ06dGA0s5/gzrgCCuuJW80
m2l1d7EeKOtedcF1KgiFolfHyxozuJvdJuF0qQ6+PWrNtkPhgXuMj/Ne8UQKo1UnRg5yAa/wb5XE
wcM5pkkxpk2xoJpE3nPZ/eCln3XDGz/ak3ksMmUU6uraxTThNLXejAaaa/uFhDnb31ZnncFyf3uw
k3M8C8rll0oFNt2X6kErbWHv1tft1e83QrEJarTH9q5xMLGLV+4HKW1NJVcwZ7C+PQN9olljfzFf
mVm5U2mDHYEvFsBJN2G4E27TE1ld2zefcCXMyOspGMWk2rbPV097/MOUaZbatIR9xtT73wVkTecc
tHBOpRWyfBX2LUii0qpgbLYrJSnbMJJghShwX1FpnV+DBxM4zJY2DiCJRE4V4oLzfiUM0sNyVr1D
FkbIC7YMSCoXw/xBt0GjZB31dyLapE1PoJhHQnmgsJdAWqkeXEnOsBxXsHG/cKBxllkaD2ztNU89
JEPIO+tMeAcWc5y9XZqoB4ys0r115OhEhonF7IOpA5TR8oOrgHRNcJ1JGZ+ytlMEUq4+MvLPJ7Yf
SQ8jovbLRKW9T/TEEESCX7DB5DuBuuz3kzbWNEW6L5ByRNp5vcwnAKEASZhWMahagIVyiLQig/EH
wT7KZKd3rf3pXOJ/5WWt+n6t729NkRrZMvDAWAVhuQdeGo0zYGWau7awL2n9hYn9hLm/RezlrXw8
bh3J1WPncbnXW4OPNhYiwg+KQek22KtXfFea/KaaAfg0SxmNfV56br6DLdSO8wAwTG6CzKbtor5p
3w98behhZGs+Fg9xWmBDPlART3d1zgHBs+lVURnZl1mQlbL34Y9TNvlsJ7wqtBJ+zAUD6Rk8AkPI
9MqjuoOyuKYxokDFVWw8rqD8ALIDJivs36Xm48dO0lTbDux5LSDGgXRbktZJD7Xijgk4HylE0Kyu
K5uzLif5PiOxyP9pqFrI+7edkV16sa/jGzKuj74Rv0MtnaKXaoRBU/hRH3itS5XngldQk9AzIrS7
TrfakDzWJb8PKNhbkkgiuQDzoYGi0y5A1gzk0VASmd3OnQjQpxVrT89V9rujLJM09C3KcThIht5P
740fQ74jgNWVdPCd3Opk6zZi9jNZHqzCNYSEWkvCkERFTGpv/u6/n2+bNmte6O7IDuUUT2buQx3R
XijdXfhzEaGMIVo5aS8OVIEiAT6P1q4fhRtAPqlyFh2iFGiDtu4V4latE1CSda+g2qwgSddpZSto
E0Iwy4qBBMpbFiQQjDHp0AbO5oyoiJXOvnromn+8LrDlg44Gj/KOk2ZJ4S/qOCkFF0QPO8N3AsUQ
jjbp+EMJpZDJcmjUUYNZ2oekjJNzPgCaFoIuJKTDIrDDVTOq+o1pQfJwI7hQV3lbxi71eJOoz7gF
vlpMVKxk55N0ATakhet9y20gAJ9Avf+NjwtIDkKDKmmFSm8z7N9hDxIIErj2c9xoP3us0Bto6oiu
iquK8z2G8VJL2pGZhdEC6zFHuQ6j0/4owMrK4mYbBOPw3I2B56eQMWTQUSToi14b4FAy7OLq+L0z
ifcxl6Y5mIHXjxVIWPjsfsHm5jL6dP9JGSFhm4UmMd5aV3bppov9Mww4/XE2iThj0owH1gsNqWJK
yjTZaSsM/II+nfzSdkjNYIl3qxs3a4spMoBhygrz5tx9DX8E5xiEbmNo1+yWBeijpZ1nfujzsRrd
p5bd+RfjhhbqrwKIsmxhOsQCckFGKz5vU0+usc94wUYMPZSUObK/GtLStCi76rhXGZmGYPpWYBur
H231wseHIbe/0FkUsn88zh1JX8BPHJcUlkUYTjc0IgSRBRRkkQfXc3jUSZETuU3x8A7XanpO+CwU
sX2W3LO1bBNnb19sOPSqMVPwTRigEyATWuvmPyxUgXgH9ZE02Ps0jndPbHT8U/Ic+9tNcp0Zh04m
4okL8HhskQWc++gjQLhPHOVdgFd85a6mj5DEQoTAbQuGKB9kGXr0Qn9iGqf4Ix1lsFa5iNVX/syn
GPvgAT/kT1W9l3mhbinpHLVV/xYwDM29sYrOc+mFx3mujzYr0xC/wrv0IwfNw57sCp1sJoxiGRNx
cjkZwo+XGJwMVkyLpfgZM1J+swanLkLZRCEX3SdH9k8WafdM1xkRRrH70rjNActGhCG3Nb8H4B9q
Z9CjqN29e7T43XpZ6sfWdzUNh1X2cZcz5TYMuWtIveVpv7a2HjHYMw5wMf3Yv0tl1Pe7RQLj/y7R
UxDVXTdNWU4Q/2RMaSE57JTu0VTFX2hk88KCgHX9vTVaqAWAKLM7ENq2385ljlPQp/VTsBYYIJNb
ZaeFYGRtfppRT4LfKDsi160bBCZlbnF6jzoaeybkY1YzBNy2gC4FAFdhqyn5g0BiCTF0lGusoSvq
ndiaNWg+Q1IKlcSmVAoptGTpo5eBDB6QGv2P4r93pbV/37VcecZ95hjBJbSNIzLdVlyhRu2OGuKh
Kurm8WghhxuPVlF5TLR1RApy2AvmWe1kjYf4DDEKOJFE9wsM/pnR1pvL7C7Ed22qca9V2won+A5T
neu0oduiSCa3JM/+/ftCI4z/QWPH+hMtEoakJvppBG6d7ok+BH8R7je7RTEwuGsv71q5qa+hPd39
Ujwoguvc7cSq9Z6h6XJ9jVOdeffnLsXV66CVztcw8Jr5C0gSmHKlqDDhyZDt7Az2U13b1gRq09af
vGXu9TNaoNLHac9JYqF2qiAW8jVCZ8oLJzGhktPYZmiqSClkNdcJOvL7ftrbZjEgnu0w3JuQargd
Dxz1BgSxWkBZLMEyONiVWF7qlztN12dtAUGLuXH4dtiKjWSYGsZmqTpmptnaTGn/NdTaI/tO4LJr
6es+ygukpQd0AZ3AmRBdS6ZttqJQ0GLGxn6m2ZEqdElsiBROFzOChER9PNcVr8sfqpBJgXVHt9Bt
FGM0CrLGF5GrkDNW42CjL4lypkYfpxIUsgtDTCVhkLghnlKmeaAwfvwxZNVQTiPNDbD6cKxElmDc
jqp1ELYfinTNntLTWnQlU614R0uYHEs2h/HcX2mMaqzU+aG1S4kKOkIA1xdfU/hwfIGLOIEkFLko
EGGLz6jWetc9JdVyeRqgU1gAcK6nU99OxBLUpivR5m9LjGp0eSMQj2Pz8uqN/baycRfF+BWFPjZB
APh160CKIZtgCtmszKXhy7Z64WFwblGYQ4d/FpfWw7JYEY0Ob8mhbIMc9nX2tDDJ8DFiaxbvJjB9
IftIewhSL0CAfFkhO3gJEUg8obc06IHpUHi3F3Hpn5go21CD73KE1u6ElRb+nWpQ1peLauxUk09/
0BwXXcHXbVnsiqk+8qhx87r/8CCrKD8VorT8te3M2+G3GVjovv4qgboV2QJAa0qP9pzTQmfGQtl8
f8zN8Vr519SzhG17dKq9+XQwNn1lyIId7DvUxISmRDRuj4x/kV4PUwBg6WCCG8iW5FpwelEuxmZ6
oIIwwGVbJOpP6KAcEigFzKcIKDCvWDV2ZUIrLvJxcAtdw1fYCGfpAiqfnm5v7Uk1A47H2kzH+Nwa
VKJOBDVVYFK4TQpvhfMVzhXB/Kq53bZbhAHSrk60lfkOMzLCGC14HkEQkVBc1eEBKoUhHPAtVKkW
5m70PjVZLIW+QdHNnJIucGzcKsv8IdfxAs9LOxL00gbVPoyro6wzufi1t4t1vGrQHPqnCdG6VFJv
n5dXDRG8/dvDs2pW0BVPbi4jducJZzBIN1HbosefpzI2ngxzfoi2tuCxcwf68W9Zhi+aJ4fk3VO8
XNesEVMbuyFTGN14PRscLJxyFNWFaCUrpmAjsVEVd9CbT7BMAgBSoiF5mcw+iPQFL32Loh/Iq/ux
ivm6hp+QImQetMopAE1FyhZcP8RMhHR5yl7uZH82YS0XNmkfhInpNJkOZ5b8zT6X83hIZQPOUj+L
BDqAB0jOyJ6U6+u6il1E3HZkfgwrgqnMMGptXfkAnbS1kAUqv4Magv08ku6nm+AbouUEUCCOQ9Qf
TsShaZIskgTB/4hYUPpqX4vEv0m4+pOX0lHFY6yuXvJ5UQGeNP2MVjbbJtx3Fm0+mpElQFGz377l
L9KmlzWL06l8l51jhGrMTlAgUp6PmjB+kEcGkZykIDQsjFQaLLl7H7u+6bHZuwpmQZNy3TYb4xxt
CzkKozECyLL4RTilRT3mblEcEWiShul2lusaXeeYa0un//ZkNSZOgFV/vHXo4EA3OWZSREHr0ZMe
3t2iwf1vJFngBOkx12q747vtRAVbPRl52vzbQvmxRQS7WyBvyN9OPnxMzi9gFtF2RJj8SpCVhXqI
HIvDtzFYJ1fC7iXuTnuvYBqnduwe/lN+fzdibU0fULPvnp8TXCwgkQCPXT8fF0jnaK7mcyWrHHii
h+arv1dRMIGNK+VnNyOJFV5BKIIEmJ9KF5OZ/u57k7mzzXiTJuYWjMdCu6NBYRqfCSN7Hj1hHySG
KAIZl6c0SwhOrIF9OZQPlQaEr08sGXh8Xf6tOYcwaWcb2JphyvfIgyOf6f8MPhtPFIs4/LI5p2ur
4e0QLMa8Z/OKeQ+Ntcf3d8vncD7cXS1RErxB7KtZyPI9D++FV+xOCdnHkFmF9/m1jOuULAKkgMGM
xXV9UNSgAugQRypn30sVduUdg1nKU+m2wldv2cfSrka+/p6sJKHeXe3HAuOKiM6ONymgLvguCG7I
51xhQqKCpBsp2mo6UIjSvlZ6w9Fyt97Y9htEOZmuDy1UmIXwZ0RNv/ouZGeJlC8FFlnmroQijP0x
0p5F/0vNNELHR43piP6CnGo6KRxDznxbePq/vpoE7oNMZkV//oL51/2T+z0ODplrwh5Q64zOjFrM
gdcfc85MtjXrqb2upykF5WN2rFka02mtHso4/Wjzpi39tixl0T7Kf/d8lPtkDacwfcF/iSyla408
wx8yTloVHssNgkWusM6T1MpPvRmKxAuJzPIEcHxmLabRWA30pRIGvvFfmFeryzLE1jBy2JTkHpun
Y1QWUfGhjYNDop3V6B5haxDOHu6xYfBLmJOH+PJXiB8tqexQ5AcD1ukGB53r1bPQXdB6wz0QALbr
ZBQ6nXRbxPckvzVfpuA8zs5aYIj8d4M0A/0j9BOYOdeGxZvEsC6QfClsOumApCuSH75yujA2RAm/
CZn79FrAeGjc4iN9ROfqPmNfeSI4bl5ajeUFHtDo11ZmcpcKR1AKnD+Zo6iCe11KGkquYQqlHBdV
tv/aKkkBiXyoV2CKJ41x6ds/zd3JXSheONtQqvKeQp4XcXrSB20eeCfuY1ktRHTFpZJD7vPwOs2R
SkBnnbvm8z9sU2QPyISOALM85oE9SlYMBWpg465Ec6UzsE3rSaFk6JL+NZIcHDAo9GFCoNWDI0Vb
RBWhmc9zRbBwJtqHWG1ZL+NzHGXnd6wBnnhF7iZPKBA1UYlsfFnZCcWZZf3xJ80P9uhATsaEyf6C
dRuHOki1zY7fsuXvhEfO1ZxAvxjIT9wQr+HB2pOzVYNbD0VakjjpLR393Uc2AEoBBclrHjDHO1gZ
7me3zzBFO/ienEqEhtxbKp52MTKRKYWuJPXbMgYESemo3lf+SvA+CfHLGmHIMnsaxO0YpDeThCsx
iuqZmWeWV3Dizm8D25bN3MkQ5O7KBZErExH3jnIGjiL6VOoGGKJAdg36tuDF42w/h4KhO0eJAXke
qZgwcQ7sxeQPUPNnqDAnV4LVKcr4mbS7ieO+5BKRHcWaa4AE/PwvxDbuu4PtTcne8VupQfpHCD0J
fG/BW53sjh3u5zOj/bAPosXT8DunqOS6sajTHkkgVn1xQE4yGWeWX9Cs1ckqLknit5ze6EIVxdbl
OHIoIexAZyEYc/lK39dQ5Fb/rjtphAJ50Bjc4/QOkHI9GfBd64gToCES+Y+QY7g2FiwLnwZS0VMo
HxfSr10IKLmkOcu6mBnkHVy8WE4DRrkfy69FvfccWk4ZLlyuOODUIIOzxIoE+x1W2GwGtbyJKYf4
/RI469JgIwQswRCUDhMmWfI8cdrd7DJgOj8EXzsL14qQjSF4QX9JHbvYRB5IftvNB9eI/CqZyto3
0dGFqGda0HPpcxUs7D0ewxio5LT5aRlIkBraCfkTMvmPpgoWU5YM7aAGRe+UKCfgB4EREHta4S8T
HQDMl20DhrDmD+QqveqdPKNi9jBt6lmen76Wn0UUdU598gFlGatMtEk/I0L0xu67meoW3C5oqVpp
czKnQ9WWY8sCJbjJb6S+5ha3zAm0lEHxk8rNlXXev3kntLJs5fk2Tv+PCYGhYMQG+0BMyqpHUGX2
6OKdH/Gle9uZ7PrD3Cx9k0qFusF5QG4Tfyl4WJmstWcua8lkMeQG0vm8sb+zvkTZNyqNYl94tU0X
gWPpLoIWBQqmRk8d3qk7VIJ+dNZ59sNoEFNT1S7/4gVSVNvbzHEcaMunVWIPnFDZiFlE/qS7MH3y
2f4WJOJqJiFsPTF83iOTxtRgaQQ2xgAT00KLwi38S+kqO93G9RZf2302926Squ5xkVGLtr3Uwtd5
nfc0V7B/K4nxIIZJ4kaH3Gh6q//1ETkzCDyGDPMs0+JhITxhZIKrihmOoBo+aCcc0WDLAZjMJ4ce
lhmco5kZvCASB1duvzn/ZOnIBFcyQFhZXriK0nVpoifUskeHdCb/o0fHcgwGjIMeane0SwNJv2Ug
BzXMU/ok1tC7wM2Wg/rx2dpQtT/JLSiMl4Lv+vCwsb77jyJi86C9QNMStTAiLiI+bCSuvyi/6H4i
IocXy/8OjrlVLBlFsNMGtQr7a5NIKGmNseUXemiJM4UKUkpDQ4RtYOmBhCsO+3LnJYArghLK+LTS
U50SwQx7lrf5TZALSdpBx4YTkN+mBCE9ZYyYuuyO2ZZCXQh1TQSKrrQ3JCuTJ6XtiOK1/CD9FHIM
ONrs9NjLE8kdoqcFt/bSSU9XrwTZ8fWh8uHScrFgWU7s4mynndcRGlsNMIoMI9jqd1F19Tm9luhv
lIpXPZGQH+o/aYCSRfjGsHiRk70V8ZL2cT0yCYhYIizSE0gHRy2fl293pV7T+NaeBPWhFhN8I//U
jEeNvGGpX+Xt7YQNknrm0J9ph9iuvJsSEnff0gvv2SS6kSbmxMnt06O07YxzjKl+j/IlHrmWsnVh
+yOWPWg/ejESoboer85kpNpi2JEe1un6br+l4q9Kql/L/ZEU34kr38zEY2Xcts1R1jOOZkr+c5Lv
AHZJunJ8HKN/2uMa1RZci5t6FmNO/By/p5oFquWwTUdY8ZzhKyT5tj0OmfG/sw3ji8oQDOmdGMuQ
pCQ/KqR8TwLyU7CW6YcJFvx4VUDkpn9FX71IY70n9DLqbQJtEhjR1cB92e6sClS6EKh0M/p+StIl
hTqvuolT8yGhVeXQMS8EcHuBY2C6OKPp0PHSpyFYDVXBkBTy+Kv7Ssra0jv7x2b0BSqgR6T8NzuO
5HM1XL6doznJTgCW9cHlsnxueJCn2zRM8aLzP59OMdNznq5+24HRPbj169LqBGaLEE2dRywfHAeO
gNvA6wOxBBM9HOrCxAaIeWRmMhsow9LONe91yan1aTdCmM7gGM0pVBKXsZC6Cm4JhQ8wZU7UQCS6
CAIt93iTII9ZngueZoJvOZX1uN8/pwR1Tz9d1a5b8alqPxWOrHaEuiMikrG/qaL6EztzonA9VnLl
STcrhwWisjwWZqm8QZbJ1WLtycoHc0Hr/hFzCIbBQWSMUo9Hru4GlMdJbI0ajo6S7OXaBXyO9mfP
okOvdHAgie7dsTnYsbpo2/B32T8D2AZ+IpZtX+fFXSx6TSXamQPNUDcuqOEbGUnBwUKlwSIToXV3
x3KwdKgW/VsanXHCm5hstRKFVMeC4ll2S+2vD9Ux0CYocJxCdZ53ebavbjPHHqHGmlHpJWazqQHI
/HKRBzhqi5fit4FQutw1ex1nk1JyKjP5JKeMDWk3ohP5oBFLkmJBzZ6O6EXNSwGFEicwh9bUo8P3
K1mT/VQKD6uBMiTPYBMHboRU9ei+J4sQbBgPO89vAOPy98Ti5ZeDOINL6pbxxBpwEdye5TDQVmRA
fz1188z3hom3t47Lrie6RJt6/wsq2hXCkBgDrpeM+y6y0mmmb101k2XWVACSSSF97GTRicNxrW0h
i6/pkBSTqbrTVSADJDcaUwdnzJLkEjkd9rZLTF5zXeF+vgyl91JIeLa05YwZs+NDEqPlKkyOyEcf
28XvYgl5o4MvHEqtM7eEWFhBUOTEMz7sx1pp/kebgn245/GTurDRYKrDFMs1+DXVVoWiQAzAzSv2
njAwzIPdKDoNbNoltYSd0lJ/cBoV6UfEmZ1AajjDtlhCAVWOLWaUpzfy9/MG8msMxfVYmJ0vS2Jc
PZ33P1knszeI7EPBYuSl8lJewvoreW9+Lv/H97LhLRLjqxO6qxxwUzKs2OViY3oDuqLOYpZLlWlJ
2tK6LC8P5dinenfsXE14rjM4oWzHG5cwACNRGvRt4Ov+FosAsfv/CVb5UTPCkiRTPsI5NvFNJ2Pi
IkTfT4NovW6dVMR8kT/3Bhs6IztupCNgY1mrfC0/tb6fcVuPcT+gSXpS6YxUid7w241AmOuMJ/IY
Bc0pm/PQRhCnHVa8plDqk2hOz1ItZi0tysOwYEhO5Rv81sYl7IY6Fbuxwgp4SXQueR+rMZwrMWO4
erDqQKCeay4p5WCFEGQ60KR5TW+5PA3r2ThgERONdUjdJkOu2WfPkdKETHxeqCwSr3hHDlvHx2vB
4+McLTikBSf+1IHQNJDJ7JlBW63pw0uMUzzmvY2dePDFi7/auqr3JNP5cJGlneeyJzq/y/W1TqKZ
fd97NqI/Kt+BgDphZdTM8fre67HX7XJGGawiUNQVpT2k5N3RPFt+EAFTxtNW+CsY9CzyoVwZlVKl
QkVVmRCmFB46eofByRgYjtkUkW/FDAbdbAoB8w7v/5HVrSkA5x6gVFWuDhPUwE3bwmP354ndS/Xb
dGjofygiMJ5u+nC1088ZXg0cxCLipx5kesuYewi4X/G8uFDKA5hy7wab1I1ZTl5hqbwS3lwPUEdL
d1zc0ZljpJ/q5SwuYLKMqpbcIMB10Q3Lk9c6aglQjKvyygInsipbXYtBOhfc+IVAKUeCoLSVmtak
etvnFhBiqzigw6iasie6YVa2I3dJvaIAvDMz/Mde+kqPD+JiMJNioNBqrS0hqeMFJ/pS7yPbO7AO
f8gmjCqWcxnEnYwB9UbURbScPCeddIyaDn3P9HfM0F8mxaAzNL8jc0tiEE+OliOtSxuRkTA17A0i
11h9kox+Z9Ij0XLH28Lyod3C2jsNxtiKPmTQJxqbw2YVtklElEyJpys6OoNvMB3B8vzVh14WQu1O
XVSZq3urnMfWoLhXZkfibVq8OiFI+qVFulbhhqHc58QhvHloM3J83B2SsYfSXK9RJ5EORPsjsrsd
A5JhOfCd/3tWlnfrZV0gnd/SDfCgP1gwtAzQ48vuVIBiGj0W3U+Cb6eytDqVySAZiis8yQcL6IwO
Ot0trG3VgN9BlWsJ4VtrQerKJPAR2uUWYqwcURfzHcfh3Rg1CWZ+ieBaxhSfUuF4JxzVFWE34FF7
gKuDBQ/C7fT+IEtnSTa6bnIT3eXEjkkTrxaJa74evUtqzYHhCojU2X/jqH6AaCyqdc36TEWys2PH
6KfzBlnUBYs2hKnyjW5zIePwFz1DuOr1i0MoAi/JfC5xHRuF4W5wQ94eCBqf7D1avwFiHmWfsJfk
E5tPRFXe/aYJJlxkkksp7Bnfo52/3REo7DxfQWB2rPmlgQxUASNo3V0K5tCm1Q+atwacZlkOtOpv
h0pSI5U37Lg6KNCyDro9FT2H8xGZZDHgypBuF0gIhC1Em+F4edlHvcZE+DTiCjyh8DqSWs2rciJo
ukaT5PbEWjSY10VlIgeweZqTDfPvxUC6/HacB/cLzY4ngYtVEX5072CvqefJacN0UmOMO2s1PS7v
QapJkf48CtM5XVhUHPRXoVxrMmesVIBPskYBzjRNlw9y8PGr2I0KFUUgug0A/WfdR/JZFG6tA6l0
aMNWjanYneVtmwtyAmQA/XRi1gx+bWK6lsiOOMZpwSWDeAtE6W4l8BwPKr6w3FmpLizKBxw9DV/w
sR9EuUy/pTBRbTQ8Nseyh00YQuDpPUO5DQ3WLrH9ALXAth3GJdxiROH8ayNOysc9uYOTv5yOsM8q
mKmLhCv2KW5lSUzb3G4xTE1iGpG0NsPU7Uxp/+NSWu7V4qwxDjUn8/ho5EMUb1TO3caiAIZE3Y09
Geneeop1dg/7TPWRXJhRm7bKky95d2exDAx0HTNhvVAyFQtbRzZfDK9i0bfvJVMfWF6u2RmhPY7V
b3RkWhYG2Eonf0JXnsbhaLzF2wAhEPu3AI0eVKnHKESVzfCrFTAv1uv9lhxZ2DPpxiOE3Y0dH3T6
wEi65k3chkr77TK8lQ88N7EVSZyk48yn+FKjLqvKPPWt+C33Vv5dH9xnVd1XoGZwbZ72e8Yz/OIr
bkudsTrNasBMQ/L2AyJVjLJrJbD2FLuIMkhGuh46RFsInh+z1i70mbIZlHUwhlipUOe8fCFsQXs3
fri6DAp3rtrkUYakWBFjgsehkdVL0AxPl+8mRi0FbOtTlL+muWpruzN5T/9cDzjLwmlvWEQKa09H
Fjq0U4O6lboKVIGs63fJTqrILDqXWOngDaofWqYtkyOPoj0bku4oi7377M+fnScJQ/BFplKyDTwT
Z+/O1nWDCtXuz2xb0VBlAIkp6VcasRA/BRIy77tiFhzkMeHaENKLYf58zFSUuHqHRq3YfgN+OVQa
i5u/ePPa/JUm3zuMijsuJqXYt/ezBiy8+BKhHrf94v2kGUxps1CJUcXk5jtja+IFxq7mzWuuwAvW
P2Z49nmMpfK8lScVBBwJFV5bZsHJ6xTnDNXnZo+UnKR/fvVsB5OAsVC+B4EkGED+LKxUR1avqqpc
4wM00LROFPynWyP51Z4JN2OULyzWvf2gbrAnh90akvCldgJMu1SXOGyRemoeTcridxMIvbLdK7k0
Ff1t+B18xpjEsLuSWx6cHhDmU/gpAsqKqLj7QbxMcs3Y6CCZXELNXyWXl7y+TFRW0/wxCIhB4JGl
P3d/BPFSbn+ytzQZzA8X9y7E8PZ4wf9Hb5DanFyR3z+RrjuoBdumAb5ienUZnUtyHEpcKw51c+Bf
5AxN5eYSEee72XfmjuXNzTT8Yl1zT6kGDL9WDapp6rBqgxM8h4UV3n1Kqqpcu0cSkY5J7z9Z0WlB
devyMhaB7mARXd6NH2jAQq2aKdSirEMFt8VuGqyBiNT+1JpBW46nIpGLljf5XYWRS08vlzdXGWtq
dOxPP4+hmfcO1Suk4i4atRJh08wh5Ee5c2tuOFhbagCYiE/k1ePJUKoeqHBqHJN8o+pV103IHrNp
s8rkZ3792XKrr48xf7sNC/R/2Z1FhpYlCgPubCEdrafs2JCeZSX5rGvHFuHrQ205xdEYnJsKhWB3
3vNPCu5HwYvwGEILWtMPN42TGKp0TCyRMA0lHyxNKRMBkXsLNdjnNEPWON5XQhHO597OouAYD8K9
RzA1C1DTonSPoOhGO7SI/nR9F3Eopag8ENdpFiY1bn37U+5w2h2EBF0MDyPuPZizJL7JyMqanMo0
l+JkSafdySME1ntNw6wTQVQ45czvIkF1NY+r+LKR7CYJtm7N4d/rYeI3RTTucwGQG2DtaW53MWyX
iet6xljLdh/pii9BKg0DtVqgDN9026mLYXRp27fAjxBjzwOtkF83Pa1OoEpODXDbYSe8zp5M7yf/
xDunTsjmnvk+2h9CI1NPd+3My4XwdjkCILBtri9eDgPKcfDnrVwL17mTAkrVGbgycjeIp9fhi7N3
M7ZHf2ZiQCJ+m1E68+Ohe4uighUzEVHu/jij3nSmxrFwW0ARbOh0T5G+H0wCjCtUGmTN0SsP9Ae/
TLcb3xNKNfJY90B+9pmnlmPFEh9LgkXX2YpQjxliFVuNxY5u6Vb4drFlAWbrkF3/Tz454lW7xxhk
41lsyAmbM1vt88eRA7r+2JTMPj46zBtBqvsQzcVk6vruTUmnkLeYU1R5gpXYwj/rIYXoVCpNO2+p
MxzxRtLBv4aNxgCWWb2YPJfB/Nw+Obx4A61qQr0r5VJX7nUK+qZAMiFeyO05DmO1WFVsBHDBk+L8
IPOlhEj6iEajSewwsLnDo1vp7qdmXbKClDP/vI9agOdHI3gIqPGO16JnwR28edFZE+ECa+KMxDd1
jf3R8mf+LwTKCUcI/Z1q+nD3kbQZg5fzlKMjw2NO52cjTqeFoG3gyh8wP/tIVxI1lGgPhJxRu1Vj
czjeQQFHcIRZvEWEKKc7kw/92kQH8v0iKvaNLcZrFUu0v+78OCkbP1/FfrrTuhnuTmu3tLoGHlPc
mW1W0UO4gbMkD8J5sU0/ZMb9N42lLCGpQTNVzdD3x8Jpt62lhCTSDgMBXb5S4TCU7DNGoPm64obA
nH9JtCL+ONWGBKt9K0PBAFgVa+AsxL6JHpnuf4M5J7D/i3GefcGwYZR7Xk/X66jrcXKPqxk4BG3T
EzcS5BrLNiPbk24nrpWKm2I54R6/5O7Uy8p6zVuse/SWpM5SaCJfBd9RrnKPQZn95zUfxXwNiBvE
bwjm0IBZT1y214LmrWIioUEnwtayUnBQrp44f0yDEth9+uEP5pDJcWWLXW3sYwtWn8Xo4VYuE3Pv
6BZlzzvj9YX26oPoVcnYDLwbH54o0kQI24/n03PT/zpEhUJN0Z9hc+EhjUtQODSwSau6oBSTEt28
xs0Joy0qDHoKCWTaTATuP77ltOG1K94gYWZaRpjbPufGZQpLlyKZvsY4UFl2YJwi5qlyPWSd9kej
uaB3hkr3QUlpybKMX+9EvCjqV+vgiAUYnEum83vnyj21JwgdnSD4D2EhdZclunJ7Mu/U8AUR61nB
PtY1Q+4vUgAFHfNBipemteWIiNvYJtaCNrSmKUbO6zzpLLlKt6kVeD5BFGMfDXMwSftGlK3Zjloy
iLnS1Trdk7/IoyI8NqzX2tmbNowLZa0S1QZE4+8iasDMvyHm9VU97+rAsOemLpOX3IjRWMtHe+A1
UmG9bZzJBen4eaYX0NytcvETByWi8AsQmpBUvjheYjx+bJzgBn2I9p5azwayquwJU5zsItsoJVnZ
iJn9OM0YI2vBxuNrp+x5bt0hlvv55LgtjrBdb3ASMrfvmV34eugbZUwYXVReSLW0kH5xguEN2TZs
k5fs0gtwSnwofmN25YLf416kAEGp6QPCyc7zHmWHFvOhhkHS5tJcFrMI36it49bQMXtZwicx1W53
mTRksfIgnV3MvyEHd1OEn4vZlq0qqmCJl9DszSB3fjV6ZYok8AfsqAftg9UBWIEyudLqCxKFgFlj
YlL/OxZnRXaBaQpOGBco6dELbYKFb91vaz3rj6ZcnGOfnVoJ/81dOqT03Hr1x01FHOSyKOe8rWfW
h/mVAUOwt6XMYZ16kKnYpzZuTzfp03b0p74n+vQxLEUyQ23anPqPObhKvYrNpV9+5CgPl1MYoCgm
f0bSmhVPGIDOpsw83BLejQanoJXgGjBuIQI8YD9y47cl4I7d2x6L0NwxMJ/VLgVcHwbK9lPm0zPq
lHYFCf7vsN9oGGZS0EAqiGBbTMBnPjQjmisNWSFdyPqjDNi/kIY6zsSmT9u8h2lAA1C/OGHB7aU7
I1KEoUwsuF9C04cpqrYbzXlV7qxZbOA1juJyoahzSoThO4gLikmGNWR9j/uWWhj4jKK5nSumLNw8
2ZXdKM5TOzPvVAvo9Xc0b/JwxL59SIQf2It0pTpEKSt9wsXZFLhBhdGtZ1k45+IEUad4P0t5gvKq
lPOr5dDdRp81UHtPoU5tMKo4iPfShPU6hIDroCnu33EUP5FEziFUAkyH386XICJlMCIwnRGUzy15
3moYPGZJQq689stYOoWkmAC8apWaTtkNVwolIGY3TdKMh1MjYlnnExbHJfNww/8p28YbTxzstwNB
23VPJTkaaTsyoUiTnUWWplt799VWFhiRun3Ebj+El9ZESIbuNuteXZmKPLHbT1m024uehhoN4huH
7fL975GlA4Jco7JTUOcII49BXyeWl0hZ/15r6jDmTqmn0wq9CXKfUX1WasHIhi0tJxw1NgkpAEoe
lB4YPfop71eP9+w1cYZ0Bv+sISQxGtnjM56bIOMAdEVwe3Va0p7nseG5ltu+aV3qi70tnFLi1bBE
N1hKm1kGxL1Mkd/ZwEQjpkiwmOKCRdJ/ANwmNEsyxKWFHBUvH6xRETpa01oYlfGU1DpvxBtXXdOx
quNU239yGfhXcMByaR7ao8RM4aCybAZGQiZMq2CI3xOK6i1XdVLjyiRCZKP7hg3pVEDkkRdJ6Yqm
Y/7oaG1HABhzvCNpvrpp47SaCCwzxxu22MeHPlKLCxNKvE/L46wwk25NSYEkJ7l2WN1Ustq+xHBY
k/5S40V4LLgAgP7TzhNQ1Hdg1Ps3ASlv1xTOHp70P5QFPdFBRWAQwjTUOoB+fxeE8QXp1GNvkrKC
3ljwUkrP+8AMkkcF5EjX2d1b1daYHgJ9t7pw2UOVZdaQTzs45YyHTbchsT6W36n2TKRko8TYPUM5
Z2Le+MAgnh7pn8aUeQqxGGGAktTxSU2MdGy17ijyrZ5cLjzsA58mDuPCFd1TDdteUoyZEhqhdGNv
x+xCYXzutj7PrEB16/zk/3Z5n1Tb3yAAS5rlqvYTxpaMB4L2qRAHYZTvOnPxjoanEWrwW7GopWZt
DA0MbeoO6XKXFiGReDHhm3XU5dP2TXZh2ORgSFA6sFZlUrqcytCytilu8od8V9N94/MAtBpwVoni
Xs2PAgYMEymHi0gbeHGZSV+x40Xcl/kbWq6/0e4CeLC1IFj7VqTHHPjKKNnTdR0r8AGX9GwOxCMB
UrXtQ3srqeWmyC64ErobIKDiwgr3DM90igAN3qcx2HDCZMCKlWglL60wxYBhPZOQDWGnmFuOHG4X
/zwvNJdAEsbVjAp0umqhroci4+zFvHYECIvUySWfbePKoYqJ1ZKZa+Kq6RlePlrHMlM3R/1nn+Pb
T0T6GXsh6b7IYIKafbT94GUZ8MNPRMienN+6YMq3f0WpkObDqhxtfPkB8S8J85zUWPsx3P0fmJNI
1MK36o/wrmPo7dKSMoRm22EyZbpK+C+bqFNG5IVDb4Rr0zoFSbGPn1Yy4f31uJ5kccWkA95sIZ50
nekQWCGzHlXW4pSnuMIilmAn1l/C/C0TGssjN3+SNRHozgTOdIJL28HBPfWKPahS1U6YOvfrQFuJ
0JYWj792y7WcaeXl/cQw8NT2bp6iRSWc7dumqG1txcA+MAWbuc9ON2M5XLtdDEuJa+I6yi0ojHwF
AkQt7wOsOlruFMWHLhWhxhspWoPcUpQD1WP/rADvDKW6kAQvdF38n6Yg8kVNbK0QwheSALMsk85o
PpThwVnstZyK22IGRZ7WerAVDzT1KNadrEDt5Mi+z+zAu99sxJ1xp09PONLdUcXcUJ4g/Gr1ezqY
LYESBq6e2nXX+mRx9yH2uoWzY56U7r1JjcXycCq2NkVKApmXKJZKrF+Momhm0027UF/+2YFZ2wN4
x5xy731/pVn+yWk5Zk+pYcqhR+r5IjSEh/W1g29Mm3AH3oSRWqZyBbHX02fDJVmB8JJqJZb25Ozo
blruQp0QHMunN2cWVr4YavVOOdJpO3VJMv86zfVzOb49MLcRTeY/kz8NQKGrsOkEEJmwKE8+wdSs
xFEeE6EENwTcFoEyrfwk1LCU3yK98wbbQKJOKYmObwZN1sZ7CfrwnIaMYmwUnZHlhRdZjcrFKAyo
WNybQl9mpZGbJlWtQMnTZa77WOwpH6rJdWF3hlAFe0qjmTiqOxo+N1aL0LK9V/AmVR7MbEryDnCS
vZXHIyIVzXs0SCrvaY6m1Aw0pmHEtfCNoDbF6+TyT85gUw0JYaqbKvcB44dtYjOciEv9Z/guzMS6
sDr8BvCwo84OxK+sFT79cU7H9lYdyovI3icYTtarFIQmLsZte+FpSNMz5hEZoDnETPvkkGoGGBVR
GPH6IQfpfx1EhEaik4EECn/VPkj0ZvWp5hrs8F3lrjffZPe6pDksZzj8Moejy6KCEpSOkzojuMMQ
vbzEZw47oi02CD6lTcHzsilkSTypzb5Ys1V3ybn5pQyrs/FUmNgntc53Vn/NW+43bOZO5fb7kKI0
+jJF5ezXTZ8uEbmFbJ5Cj51OJIrTq1HDvh04gGROGaq9AMisO202+dFBeu/Xn2j4nWevosNmoC7J
WRwh22fWvtzFqCmYi4iGJAH63pmma8GlD9oE46W6+H2tDLyq0I7QIzdPJLssbuckW2kS2DKkyMwg
SOiPhW0eTIHG0SlsXUaFGhlubB47jqb7gWOBe0dO1NZsv3Ri2EgTsrMHTI/CA4Aar//9Vannw8Qe
DZMz/Vx/5hqby8waxoQshsBZrpBJgBZo5M/BrfybUH4jBZJcipuo5n89lGgXcUQGpfiBvpjMm7oM
X4JQSTFjMfHFc25ia25n974CaOtJeMArea8MjVzsgIB8oKQsxnIs4xQaC6TVrA5V2ARBCunX+3Kr
syfj8QNkdFG7G4fE/Y0rv3LKr25Y/kkiXCN/MLMwAn7aEMqELlGF3OBcY1zi+N1Os1s61KTnzavm
QSnAaIihHW3Xx7V1GJ/1yFJHPtOGBmKZqbMsjkPYWYY/6qxgrHcD2MCSPMumudNFI9K5FzwTF9ie
AUoj7E2EMQVPH9cNAyCe6jXxQaEnrRRxyg5MzkAHCZJwSXU/OBr0HOAqQ3AP9bMa5B6ToMsX09E4
9lGVFYlZMwTL2n+RIYWV3AKB7lquwke34GWXDDSdhWQPlHYbNbUlClK0ExuiHhNg++RCVYIlGG+S
+CPqcmPHEPEoA15+ExthTWswrv9KycdcrUNVYS/tzi2IMQMWc6UZ/ERC2NY7ZhYHXcg5SyefIRMm
DuXiO4wXtL+K2elUDxnZ96UKZmiUIr0HcgQVzbrOrrSTEeAlDxEetBHfDrolrDqkA50oG77iShwC
21AMW4Wcz9jfQxcFk0O3r9oGr673WE0q5S+6lvehjaTVTUmCW+Z877dDc166LpM2+CtxaCz9EJi1
6kKgtfOKHAx4oQfY94DNzMzx51Q7Ltaq3Y0u70AlcYp3UkouMVKU/dhECSKfAuiVpKt+/rwBFI0R
3FEW2xn3x+br0o2UyURMmjtBuuURXGSZhCLVST3aL78swdptUdC4KF07qUD6rG9sHH4m2pb7wIjp
+o2x1XGqWTdQMErLknBxAfw+5HgJwc5oM0knMVyq7p0tzgJYQYD+E0enqVkhJUAOz09WE4MnWxxL
MbF5OzDxRA6q5hd62bj5ZTpN2stGxP8eoRarKNCnIm5FOcrx5ok0QCQcqnuCuLx50t3BlRuM1FWc
VPEqAxMQUzBLIlGIdz4JyHLDf4LHjCpL0On4+VHPHv3Vg0xMOPOJDhdfp9rMzHFWXqZt0eA5+RUc
eOnoeyK+/epZWqrcOzLe5mhJujWyOGh1RByg0HsHfPNBoshvV81X6f6M49wbqa6zEt8251UthQLx
iyb1mdX7/v19fmp1Kl7cJktrMulbE82A5BAtL5tZiMm2ykcg/ErewgMQq73QRDHPcqteKYy+koUD
gH+34MXnHOyiQ4YfxG/iDpgwkFihtg9B0hv9GRcE+CO1+PNxGUv2H+yfXWxqn1p0Xj72WL3zfgYY
b2xCjUql/JTACjGb1EVxghrOlLwptycYH5077YaHz4wOOk+xAp5aOEFSjAZC+Zc/vuhmLb7OkrXv
QtwoFOF7mqhuJecVifEigD7NvPCDG4uDESy8+/5ocfLpspMS24CtKOeRpQbKrRMgXuDhUf8nYkQD
Yb7WMDVPEDVm3A1GAH0ehmwHtVLgxKXVBnC6c+VqPAvLt8xFI1CQhu3B6zbAKRPoBX93xB2+7aE0
GvMi2PKi6iPOMSSY5Ag3scApVsWu/g7o2RmJACcxzPb9UBdUyZ82GZn72uTtR24iVEVejjYF3NII
0eFwxk2M6l55NoA9RfmynsF+pZxPleEzvID4nmG6dCsHtbH6H244Y1AAP7R7RYSn4r+yckxYrost
gxlNcQZCZo5R7SXjsGKT3MAlspkQtw123hlIVFJxhvm4g78zSm+csCbP1lBPGwGHASaUsifPiqb5
j6+aR2RPDcqQPjJXuqTxfEBPgiTXraKIevX0mzCq0Jhk5UpDj/9LbDXVFSvgC3gNRW17PNbdo4I5
w4eStiCZMyccmm/1BjGtOwEuWs9r69YmHyaZiJU4TXGoEKR9se1rl0cAEQrUjpCgC2JH05k7x8Na
0up9rdnjZopgsVIITvGd2Kb+PP7qHF3LYBRdki6rb6f2/Ht0TJpgUzaQM+ZmSxB+vHBxHHlrVQFk
uWUaqtlP8BK85Cea9SO/xynVVNWBCzL72GKW0c3MBedH/SaZDZew2U3UOvbCREO+1/8wWmQfe4nD
boMUFRUFj8V0HRu7wYdQrmcrinGNCekOPQjn/chylqVtHo2czgWvgG7DpIJoBDl2mXEthenkzBB3
pkeMBUKhr64NE18UUbRmakN1hcHM45bDfs1G8AxO3IbYpFqnNFK+NHsMO2ROPzIuX5nYJ2pEDSLa
rbkvdm6vPNUNDfDvBy24ttfAR2fT+H//3LpoxPIS7kdyzaU25mXsj5xqVN/5KIAUGic9+i1C1a6h
E5+sLZbSZy/yXz2X3VTJitvZSOAq2PBXVrFa1VuGLmMi2EFtoSuMbulo8OLLzUD6UoeiQz0US5VI
OjAEG5YSu+3HKtUVPI3ie80eNAz7XrSXmlRIi4e49lialykovAqqtLAVu3hUStkvACPBcxyQO3WF
Rya6/9pkbRXjWCBMRYHjKgTeXAjE4NveEZYhojjmfGt6m9yv9qKOpvj1ZpY93iBG4psxHbsd/kaQ
SJZU/+gxXNyWr8wluX/8n74zUfpMWVb4VJD9DRX5N8YLwt0zEkdkWwSI3X2qhatp1L2j+WhVmEJY
6V68A21t14xPwdlTEef3GVBnlAfCb5STqR2Fn7s/j20Do2gushHhBdrdYXesHdq/74OMHMhK0wp9
b23LV/EE0IZnDAt5PZBh17PuIWZOalEoMyNmlZ3+0YdAD0poG7hGH19edHEEQjuDTdDEFNKNS428
4iF0wqE3jnXkBXohiJrA1KmpageWRxoHfVsSvpq1/YjQ8PgfNOAmq72pigAp77GiXiwXECHZSJSQ
qX8DPmrbknhcUb4rFnR6P0J7V7dmCCAelKo0wkowevP/HTVZlRBhazj3/TCMOyvdEz1z95KG/5bH
XHV38WC1XvqB8voTK8pFF7KcE0naNAEa4i6h2w2nw8GmW8pWbmgeFRb5jNnQ/QhFA0uT+9Oc2Z+l
/LmCgcxD/T9eh/Lfo0snMy6K3KNhBLFyONEMoYS8n/gqY1KN1Z1L0OT5U7WKvTGf+xh+p6+zYy4C
hetE3/v53AeeSndxW3fesgQU7gMCWjeu9sEqLP+UUV1OD328pgsfXSwCo/irj63PaM2AYw1gHUFO
IBvsCvsWGFRH5/e+obbxxRIft+WhTCgDq0yBwTIGspHMEqYHQ4WgsCsm+kCOiyxDMT4Y3nZC7oM2
hegDmph80H7ecia92boz2clY88Suv4GS9MpHic6jS2BmSO9MtWKYUUYlVlu0p384K+I7hqy68eqK
GNpUyTF6MxoVe8Nn1HbiDKlCmeQs7V6zxSvOjRr6osawWuTGkluIE++cHAD8Sv/ZOfyJZ2Nflfwt
qEnklYmNc6r4xTssxtCsNMEGoBa8tzQ8o2Z1vYZ2y5rDgleFiNRfXBtYWiM7m+nSEI6liQURXhhh
bju8X7Mf9Nsi1csoJ4ySn0r4CdKko++CqhYCD6bWp1povJM0bzZCC4/pUAPpSEAxfsNb6y89cY9P
4uco6QeEYKevIq5xlytt57bRJjLbCviK9dtLqOmZRQ7ZI/REu4WrAds1GEht9EDUy2zuqvmsxX2X
uKFZa124/+pFPj8Gq/2z9cYPlxzvfSXG81wx/eAu9dmqXdmu9tuF0aA/jtIBCM7hRe6EkJJzbvLY
NHgcn+iCDL6KUU7ljdq/GlGdMSl5I+xKSqZxzIY9vr9k5fHT/qEfeDYdxCRTjFrS/5trpWUcXIlf
UEAYUTD2M9yDr4GUerIHD3/0oQxBkjfNZPcgdJXnzMrAMQ0jOFUj+KTeRNDZtOKNhWJzOXSabBSZ
Ij5VXmAnzYSUNUjlLOUVWwN8FbwYwWUh2+wzxC3lbJGKU9nKPevY8CjEH/fl0HMcJTdyMDBwEj5N
Xo5+yelAXRRy1N3RjGeK4sIIAL17pdBhb9roARzElvjWcEtvPsd1cjIHFQTkXtSZw+CsqIrzSQ5g
Z9Hf3XDmzuIxcN/sTxQdzrkXitCCNwDDDyFlULXmMdX5DDMX6zwK7mZ/+DEWZBaIXHw3mq4FiDmi
bfa7W45eIdSNMhflqNwMnu/7FoHNxu5KdCSGZUZUkAU1GsoRCCZeIWG+rLx/5U9QDWLnlNNY3kEo
Ar2tkaC6M38/X7VKoI1bs25N3ADbGorIg4fCN4Fv9B+0eKz2beHkYj+irn7ygB+GyI7XjieZxzdq
nTTiLjscgOGPwFatjgbHDPUkR4SGRWqE7MvMvqo8nZY5oVrnZzQGjyo5aO+tFiW5/BZWxY+/4Imb
Vp3MMLa7iCNZzv7p+dOOMS41Cap5zFHd025ED02RzIjq1zkjsjfyFVOP55/6cK+DvIsrTja45ffl
9AGOkHz9chmq/hOg/aXyFCZaLwCuiOGRISYcac/NnaezP7skIDM96KRz5w44f2M3FSuxRZYwrP65
PiwHuGxS2FI455qktKgDAD7tAP6mx7ItwuBkMcPHqS9NA6YoNs59UGif77ccaSLnyfWp/4CXyg7g
8UOVHunhtlEe759pKRPn6YPr+7AK62G1b5dL1tUvDSvTuEb2qZg5JmITT6Wdx1da60UTvi8h7R7V
nTN7ZwM8u+0m+E4S77nqzs/i819bF1KA4k2W3j/F/4EmLIsiifg9Q1NjkPvhK/qiQpmDyWmNVxBD
9yVOdNblvXRjeY/lZ/7F9/nD4Kwxyt2kCnKVyQ/aRVKVINN66soMqcks/MU8ZIsQ/s53ZvOsA9RL
m+ED62rBPUV6tvqFRViYXPWNw/pA0I4xUHQ2x0TMXCwATZAb8qd2z5FC6f5fhOcMlV8iTE4f52wT
SPJaLiSPGryBTCtBnXrs9faeXVHL4jjkhIGq6KyI/t38q+1qeFWs+hiaeWFKpV7seW/etqJz+arE
1AF6ssF3l8nZhX6QHPPbI9vZyaj9i0vZ8t9VLVLNO3lLGgEH4e7uQXWP30Eu1sD6hZCBeoWU03Yk
1oGu9smAr3aX3DH8f8+/wshZPvtv/gzwphwEtn8A1F7zihJlYMlHcoxuozqkBtofQqAjCJooKj5r
nhIyGGRvdPIzm/oVWhToTnCMCWtML8TJQNdfEC6mAcPVqJW0lpyJ9Gw3JGiCe3GLXJfJdRoHjiIP
xzxD28yoqEUmVgJA1wWLIFt4JUIuux/l/CBgooGraDm3dwVvsjf7jUpQTMykzigMyA9PK9BkY5Ay
WuqKFeGuSsQT8E0RRbhkaEJ3nlsWRDeq/MfZW56AOh0/fYFv4Pmt7UVWvqgKm8LqBL88ybD9IBJA
UOUYDuNesoOKOCpojCY4Jc129gEdfvrxGWLyyLDKxOfdVeW97Tn8Wcqyxvrm5jgzunTIG2rEJNmz
fuISRG9W4CyQddt9cva3rdpMYOeE1nkUKrK/0QQmoT30il767sL5hAkdknnUmagg6neku6BH4z/O
d+j9LZt9kH6tJdcvZOM+/+PxobtEyTCrjy7D3ubd87mpkReqOCoPGV3N3uqYwfWJdi0ytRs+tCLD
ABZ0uT8gaI0Iz35+HYoZstPw3Dwe6AUYDgCvSEuH2Gm7E78O7iy7j7YHwU4GevGTkoV7UA0egm64
c50fnCp2tcDnCudoAN2/KouUuRv8xIrqkv5wfKUUhifpXfqZxVo1trB7+lajC1ssLZLwO1ge49iF
fqFg4HOtMQWGxvtsESkXmQAas/DKlfkVVWD+Ku1B3M3nYZgdJEZ4a82ieVgdSHD4au/PVpsmjlS3
xQBgBIPf0W0/2KBCjw9iRHJzwZUC8wkwlBHvXZLt56mnBkUOHFo6fyaf5j+vxZvbQ10q1+uZmOlj
X45078mT7s9a1BMpGeU9PF6pTpMgGkaPdmuPtcUkdAGG4ymD6Fa4idudAbW4Knl/wKNhYvFtHN0X
BVPyjgBfKCh6ThZmiDBVqP6AZ8RZzlLl2ofhR40ZwjnmeKju/ddnrCfu+snU4ST8ZrB0Joh2ZG3Y
amENJ4ly1/+NGO9+yLPpLromsx4yWewVntRI2Of5TWNSjp2sq6V4l1oxIMKIbbxZZZqXaiuqf57P
dyYjlbb7TOfFBCKwWybjF2uNFv64G1VarCzHxBpi/I4w66j3wmDvQ4CW2BxwmpVDQfCKBVu5VrCJ
VY4SciqnG7W+XYFMay9b8lN2EaWOHMHEdXdOSnkH4IQ+KyrIeCcnVg1FwHjrNImIks7LSq/L7/Q5
kInmURjEn05EGhFUu7n13jA08WNOICznIlfLAAQDjfR+/bDgg35gE1MGsu5EKGb/VuynSEwXR6DX
gmwNM2Usu7U6CNJkIT5sRWlzFYuq3vn/wQzVS8QeBXurY/mbMOZxT3cGKqh7LGcgwNPYrT8ENFyF
izLA4X4LnvgvPTBGJeeKELjwyfL6Xq0xjNLvKm4z6my6sgnRX78dNDOlQYOtTQ8jIBeV+x3YHYuO
Q9WUk2u3cQmv1gHMoYIotde7goS/yPtoT1T8/DrpWOXcQHJRPKTnIK+ZfACJxP6cEPhvdalWfZvR
sUjcPVvIzUXNGPsC3BuvJQcynI9+hjHSxNYL4ygegjd5EIrV5/yxpNZXrKiC/3gzsNcfUGM7kIPu
txFPZKSgLjkPyqOwKVGYgvhTdU8LSSK5HUMgh4aL6F630XBxtS1sOQtkMA5+Gqylr9PNhxdNIC3h
NogJSftJGPQZJkd1DfuTWl/7y4qnv+4xzKUD9q81GthDZ0UCtQhdfzKoeLV+INWIocGyn3y4csMs
gjLHQLvZklrMBlxEFFa83ASiZAj2W903gPyUONL5uECDtFrXSyy7ibyXeU7m7YXPjC5mqjiPoxRr
/qka7xoAeF0YqBxidFvGL33WyiZ+zyU38Szcyr4lPca5BPm92F7SBTn44mkpq29MX8Uu3odzwCp2
oDpQInpijX7lwd6DoCuBGECYm22vG/uboq7Lo1CGcZAwEMtKg4qow7jehqTLToRLwGk3kG/b2P4g
7HF8dNdxnu0Gl7Zi8lqszEmxuXnApLo42E4AlhDJcwzcjqLdKtle2yTPNrcpAO8r8gE/jquGE3cW
iUQePWSiuIppZRjFObPBkfzMWZnbi+YBvi/ZwdB7hBL/kHx6uCksNNhvDUUZDvpVc+GyZ4CIfJg6
LmdaRm09f5BfWfg+L+5WVy+ukGT6x+6qLGKvC79EqWu+Lm7X6NloURZtM/AXkq4WD1GYlmsTDa0c
8hBvfYQUGkLuELopVZFNHeqssRpKnVtnfkEElA303M2PwoUdwXvKMF+PAQECLnkE7AX7fRwTNt5C
hYMaB0u34O6riZtzsiGyJxxMsOBiMZB+UfwzikhpQMFjN5tqYu/30d7HU3L4vAOR+3amFxEiqmw0
bfYCLlkRsIz5TogHjlLKAeYiOSzv/Up7yqZ+KGimVSe4xIVqH+ePtXHKGfmYWTbS9+TYO7A5bWKP
cP/K1G9ezFSBu787gc5KYXm4WUicdano3+Sxuq0kgMkUIRA82OEc7ysc5JfkqPEy5PzOGy7W9PRb
7wzAyT8to+YUb+rB18uVfT/Cmu7uGf1CX/804+DqB4RUcfrHTqO7F5zgIGdDKm5ulbwoJ68c8JFE
AzzBtNk8QTieQpz0lb3jF5lVa697tUaHuxfjXo4/rXwvHBYZvTENmkphDuNE583cIrTB7EG/ZO9g
8ikMznlEJeuONVY/qCLenPxzD8eTjRuOqgBVinT/w7dYVR04stlM4TGaNy0xzWwb6t8YCB8MUCGW
FT7bopWiMhLrz8Byhww9/CTCW/R9pZPSaoc+Sq2b/phK+4Zwwk0fm8UdII+b7Q/asHreGLlCz8Nc
bxBHwioMwZp397/Dq1TzIfjLS87ac83f4lYoEnKnC8OF00WaSiIcvImLiTQTx7PqxBhkYEp50YMp
Y3KPiAxSs0hPlDIwltS4bZEvQcVQFUYxUEaTWXOhQwoiw+VkvOtd8jRX5HN8SIQqtxhjZpzFvoq/
+Ynu8xqLNf5Bm3inRtagieGdvo+kCYdLjv3iX6jdrCx3D6gfo1+nHsIGv3ABud7Z0VyYvk8QSDfv
msf2bXPS4grjX3/LpRIxChR3MOaiNc6C0eRc8EdgSAtnLwpeqHeq+VLtC86WRMyLBZxxsLRw9Y2V
xlTdw3KKSs741wHtOFHDmtLDl/ZDwMj5ptk6N5B4r5F5YiJL66DKTWLXGHt53NmouGc1V1jYFD0c
SaIbZRcujmXWlWhbtOwxrkvCckWTCDr/1K07xkN1dNVs4weZuiwnIAAVR9PpdwfZ8cjJq/uRmuxu
SMvSSJ+cGXC2e5jRmkUPT1WOqiQRb4ywzkWXesEIhtGVMlpc2XVSAdBa3HqzTg7kEruvvgyIEwhq
+wqjGQgUMrg5nphAW6pcCTib5SVmPuYZcLDh/5wsxsWmIVso8PSqSGmI0sN+Y+Uq5Ha9YsrsUG+U
wNDSx+Lv+6qmGbYHaW/BzARbor2fWiSXD/O+aYPrM4AdXMHCmTNbADIlt8oj6kt27Qxk8PozqSWY
Jryhx1+opcTdb+umoas+evMkTmPLgB/bqThwFllAeCf06cvaqC4ij4Bz4DHACibTr61fksvPhJbR
5WISVLr6Gc/jW7DBhroiW1Ln3DcMa7cN1FC3bJmkcBuo9z4+lqJSrn6PZI2vdDKaHFemuXJfTepZ
GAkjYRlFn0QW53m9JY3EHz3uDpcrF7zhEnUNO+GzzYxvuTWDB7c2sS00uwF/NPhXFr7GTsXWplnO
PVLhTktf6b42wWK0bo6hoEKQwZrpI1vmWtvVKPX1rgzlj37zreMW+OADBYNq6vk4MSw4y4BBliBH
dyT5VbtMUOUgV4wRP6Gw/a9SI4SLLb6q7RN5rdECZxnwGsvESG02CUPcaMJrGMExOApZe8sr1jBa
YXpOiRiJKnTeATg0EL752RRTvkZseRhpafgTUiBUY/ecMDd201FOZeFD2Eb1dCB1D7VSMabIPsfY
zOa/Et6mhq4EFFmfU3A04RP6S909z3FIKhQDXXB7xQJIXe1efSWhOEIP52E12QdueKZ/JuEPCix9
tKdWn+1WR75g3cth5Be3oB0BtyYxpSSOpr65DHByLLgs8k/ANb94CMyK7me2YIJMQpiYQ8tQCEqd
iUYW0fkDYaSx9XoNLLLhcyt9M+61I145cKe85OWSgg+fVzM4pIBxFMZacyTYSJe9rQlH+wea70F/
EtoMIUdVfMCV7bwd0c70VFkQzC2esfmK29PBKy8pRDc+D+6pvQgTPhY1SHikMlw6h+7zeio7jj/V
FGcZjcetzaa6oUNVVvOJhcW6/rVSy+GIpfQOKwRJLV0sjIDeE0CwuMLYg6IiZnJqRznECdMq/kLj
rUJIIbBc3qQ5bLJyvbRZLrsfEwIA10B16k+0LUoMMjuhVM+/0tQTSWHonJRSiomwnbiwc3ugoTLe
He9KqHL6hLALxh+v9CL5AoIRX1bGXaCCwjZFF7cfwIBbboCUfm8aNVuYvxrwJzF5BotCZOGpGQx9
N19m7F58oD/O2VWGsQMbi6t50/DWOr7O//lc+a6IP7lu5Hq1zjZNGbISh5x3H4Op2FKuttkwnYoF
75LMoJuNDWGg2GpGGof+4AgrIvUjeFw9Uvbsi68gCUI+rWc3B7U1fDBNldH/hvhttFcSI2lFLvzm
hqqJHDf5isoOPhGc7tnqgwFZgk441FwqBP1FyJwAlRWM7eDlqWwfQvT49nRcW0SKXpQOC1ZBkYWt
fNE3d/0gO+7RvBKPMlqL1YX0DxnRSEje3eH1m64A993wAcJ+4B63fsiZeddxbHSFLf687OZ6OVF9
rIo0hQYdDt+KprzSXQzIXdaUoc0uTkDQZeIpVtnimQc08SU6UQy8aON7KSnzTe7iKYB4Fyd5Xgee
GwZI6wCLRABNJ8iM8MR/FsuVs3bi7cMF8MSOY6jAOA74z64cp2vAEAqgWorqP0ZbJc9YR0e+KC7j
8AlH8Bw3bIiA4MNzGkivFHOscIufmPBgKzlL6zqfh2eouaZKw1mytR4XxVUWKJeP++RJBc8Uo6+O
VTDh4qqMWEJ9c4H/2suZGImsNR9ewNRmHxw08JPMr0Lq/LWr/gujAhvsDmHsrf3FUIAri7SHv+2f
7tDnJ4dnTZUHI+VLAuRuIEQCRyN55brpcN2XyvqBppAInLsuKDNPc6L9IhIKotSVxl8xs6WcfyLo
z67/OTjtBc/5Yn70qxaIAO4lmEwQxcugxrSUgRNlWtNXZtKP5anfDfeRKPgRLZzbxzSeGALLymJn
qhZ31u8rDCAxCPQAMOxAT3rcE7eYla7D1/hTXMtHporgN90dfuekhZVPAVZzOUoC04r9OmqgBYPV
mCaws/Xz4Mh2FkzXmZ3u1MJ4tYk7vZdHqNrdhpUTV/QcEbdOMK6QEvO30SP6cDzXamhENUtLsK0g
LLDRdxO45PGbIvZQix81wxAPe3jL5mKdhOURWc2Iq4/RhpfrMaLTGRVUCXF45O0AskfBbFwD1ttQ
vbGltheGEyF2LMVw0aDy4duYqbH51c650hTp04YH3SRFrg1uW3hPABTLRjaQlWxVwNFteaBAhhgx
bzgIfHtiY/8bL4+A28Cr3jzzPygjuMn78lDngolo4HjLOWEFiToVABgfpbhRQZaIGTE+9253AGuI
MYY3m3EreOz2cSPdT7ZN7rMIBup+5vUe+V1ZqxN66LJrM2s3KJrmJraU7/mbM0tY9RoaFqiuSOOp
YKV5sX9qwNdQS4CuHW+IJTmdjr1hmTtytDZ5+fzlnE6CMussPPf0/uUv2OKmZh3I2VlQLuiuP5xl
oyjxh4GtJPfvbJzOPSjKDAlLdT/uTfgnkjQfww0DGmGqCEkZJ6mUC3FAPX6SY/w35La8U86geliB
43t5DTptoL/D9/m5qyG9OUZaeSqPsL29YA2FcaYPqkFboT4+IMR6KPjy7GAIHmPMxbsNXVabKf6n
jTmTVpeE+g3GBVy+Vy/445kZqO9uoS/sMPZNN8RtKRm8e4nkaVUcLl0IOM6J+yNOY5wH/v2vuMKC
e0jd6cUzOzbb2mz959ifd0Ppdw07bhIM3tL0ciAuNVOJYEi+vBzXPy34One4rMWGlf4SZ1U/rbWm
nbLzK3mvIV+1DE19/0wOn9RbCo+Jv6caBnsRLZNryyGuDo1351EeZAKXuMzTHCg+W5WlyQUCk8aT
Al81vIIisQFkP5h+xW0Rbjeq6SfE9jOKaaQXM5u3v9i4DZIrSxcZpIJ8gy9z1D6gAcqOALwGFh17
SHeTsS63NnS+qbEo4LiO/NarFSRuAt8kgLrX9gcFAm8VekPXK6FxPtOZMKRhycUr4gaqeLMbQ46C
ZX5LRPCPa6iH/F1YqQaJbgyjKDBhxRHGsaQEcAF3mlUusIoG0ShTPkCIn3eTnnnZcS2Fpwunmrg4
LDVi9+kifwTaR4hiEhbcj+fsmvCEmY5GDFyY7Kr8sINuoF28XGp8hagNbcVRQfuzEd+dEo0V8MdI
kYvmdvrdS8C1wsatkTU1CFcTqGgngjtTVt5QJHYIB4XRztxitojC2m0XQVgByrTaxwTC0NESrqNP
wRsh4kslOjtvSOZMvjno9YQP3hAU4wiZOzRmLR5TAaplw55jn34W9bAGzC07heGyrlamIOywmItb
6qF5Hp3N1IaqER8De33wdrtV3ON9PkBy8HSdNb+J+zLkVpjNK4Ni5OvB7zNDH0AtXOjpzz6QLi+T
cpb1cPc7hGdFvOE6HnwEtEh3l1rUZONmFvAc++QY0nWNNnb0e1cX0wkq9wIY1cm5tDrR1gB+viyR
gCdduHh3jYiZJVeqC5MN4OewttZwgno8a1n7XjWXOVNHRCrxzwukbPKgv101pLIYaWFhpGHGj2Uj
UHOUy4T8Yz/rHJ7yDdozeIjbtD7oR7XvrBhEoT18LVxbVBYCwc2Gh/IDZKWIH3+zBLPSDJicSsdY
UNaXBHxIxledEpGQaia5jr2gVl/OYHeXvC/l1SxCsmlmWSUt4AQelAdExSU2hTM4tb++0Ojxi0PD
4/qUm0FljNvA+wx6gOacQTLOcPrIoJRgIpiKEkcm2jVPt8/4GCteVhQp4NNDLkNRH6iFgj1x1VVA
mRuiEzf2HJpXdtqIUGfq4obFI9yFW3AAmDopX7eZIO4llAcDIRTGIjOcF9Z3Recm2FY8J8ckc1zw
B32aDAro71c3tD83aB7NE5GDnOAcDgh7pVSO2SWqMclLXPUV7KnknNosIuDFfCohT+JzYAz6pQkf
17r04LIgRAVOmg5AgaQjJFFhcqWZ8vDZ7IIZ36Tf7FeNHe0TvJk0FDA+HHoZ5PNtHRhlmqTO/jgs
8kdV5qE7fd1GHr242KpzGeyt/VQdreMnWsJ7kFusiDR4qSyJzdDh/pS7vyjwChlbciPMH4OU5zSX
HrBedmwu5Y3FlM+G0AqQOUSrpIe57DB87aoswEL172uZ8G+xwWa8R8I4/05r4mTdpyZdDphX4o6a
RYaSBVWDlwG5Iez2VJyg3jyYRn8j2NInlX6xoxJljl1wiP9mdYb5P83rDApXDyq3OSWgX6sTnujm
gvrWEgUJH0n2mPzmt6Gyn2N12nDEbYZOeeSc+9u1IvsEX75O3pXzoF7+PEt9a8m7ELRfxVKzPWTK
uApJs2/PuIDVSooxhUiJwqqLPGmgs6N/hIr6Xp1fnr0cbQoq/GKB1fCh4bNPxdkEXZUb3cEAXgk+
anhMaOmiWPYR7hPdq1SQgW7GhtTUs2xm76IKjRl8/vdKySiqROjFc3W0CvqGZ4QiS3cjzqzAy4By
Xf/JE4xdtOgXpBDgeHs0MFZ/mQGhh4V1ORGi6KAuyyI2uUG1AvlROswD3R4ECYTeXM+C8U6vCvog
WC6/U5Z2LHCq4dpibZF5JzGioD4MC1zgsEjxxaftu8lOccXbcuWsXjmdlM2cPt9uqtgmv6ItxOn0
9F7F7Fq/2zv/uEgzrWwZEKTr+Ji4FKj1W6a85lVMYB1xNnxwsylcT+U1XAbCst6aM2dwXQIU3rdk
Crx9gmmSzj2I9jlqRGR92USqvaV8JUGTasTisPGrhcsTzPWhKAI4i1y9Bbn4A43eMouy+AfQQCfS
FnS6JmGvGX4Dzx+eG7cKAFk5isKMklJQ7W2CHi2P5MXR0s2KMCA7BWIU7ggak8y9drGmPdFjaGbH
30zfdGm4mnBLHSaCMYtVRFXaCQo37yhk1ZDrwiN0Oh7AsGL1Tawj7vYJp5wC7YVr1pTcDAvBjWFF
WyJxOhAF+HjyGtbcCn4sjJp9KbEtKSB08dI0/XW5rQe6XCfYq1jduFFZkb8Mjy1E7+DsUHxaV3W0
qdljzScYxn1LJnsXv2B+RwiA46Ebs5vKLd6GMhES+RT2wrP0Aci6M+ycbUr8SjzCGHmZxgVHyjku
rpKuwBpHaDKjzoBxoavehXQe4MalYH5ogWNyPe5g7FD1kko3fhhI4rftgN2fPyC9RxUTZijw76RN
QJxY5/WmSMPjxG4gSrz4IjjG9EYzHJw+NAjZRPhenb6mQRyGQGa3+eGc2Oph6QTSdWK+UcqtKr68
LbmIFIVwVw3wg33vfwZqOcrrdBHK7m7URfkVF3JUqNq9tKNuJlJH9myCRtN3QhpjPP4YdrEvhEwU
TIme/8bp4OLbDIY/jtIDZIOS17fY/+yw7bigRApmlsMc1YWEdp+YktrioscJo1HK8jacnQkVaWAr
Meh4HvW20sIwl8OXrj2zdfelRhmjPyzuMTXGvga31gIplfxtQ2lECT352pEdnogf3bS+F4Ss93jh
CAv0QfIa2utidbbcOBZMcFK4jw1FvedbGM+Rg/tNe7g9dYyP4pxSsGWuSrzX1V3llJaGKOGe8LZu
nzOipHr4/Y3mQsHbpm0Wg+fgLgNZQ9n8UQCZQJKVTEMBTUk6uzwHea3/j6IgstUfC4/Nn4267VFG
8PZNyzPG8NyIME9ygCbE4jp4ijpx7t0arR4nXE3aQngX9+Exncx0QXOyCbSza549dxmsuFKPycpQ
JsYO3BCSo68tcLzxwWz9yKnzKVGsYCNQ6AOXm0fmJumhZz+xIKGjsGluSWoz5VUndFmvbSVWjmJ0
wdZcyXGeUfkF+LQyONpMOFaaSPhSYiuaTU0OoIlukX9Pt3YJjyRs1P5DlT6iQFQg1Oj3nmsULdSc
/iXzAaNWKnIm7RqAxs7A0iqysSk1ol3cpAmszLsQUH150fhxSdlpNnyg4GsCX7P3AXld06v1nL0I
PSHV2jLzU8ZxmNV0q8rOaPdERNtzKFmZ96VVO64dUWKeJu+rDr8zz5/z7LlC0QPkQWsxWjLgcSPS
Mwbut8wOpWcNbxLSX62cVMrprxZhA00w53gRM/Zu/8SEijUzB+kByEpZpT0unc8TY2rb/nWhAG28
lneDFsjyT54XNt6Jr1rB47QYrtZHYFYJFghtUK8LK8TmFY7kLtLyyDl2SqlC+PxGdx5DtrZ3RrAQ
cnbfTl3Hk1kg4pDLtCAhk9eVbL5DdMcuzt2bfZuR89UxRDy4JNaCw5nt+v2qvz27D+jbAATzeH4H
IZL4xoD2EhUPyBlPFWQkG/txpCP7cKKNsZAKNwCiBq8IELiiEUFzVDdrLKL4trYE1SgHbxszDRGS
RVkYFFdZsC+QDiNCsLet6E9mnSF3yqMY0NBxn1EG8ICuyfjfRa7dqP5fxgTqrS7lVbOnuMkHuDHe
Tn6SgFoMcGVamttdiU961HWRZZdMpYJG9Qoox6kBCxwN7T/7uC6+Mrty0g4RuJchsjKzBfLFwqvo
Dxoxf0jxavi41EyqgzhErFmthHp1t4Gk0tYRTt8NqA2zihcwD+zq5j2xiIS4UColVdorcHPL1hWt
YrRqopB53odbZqjllyksnX2YO21HL+V2wYiRmwth+GgxyPrmWtlg+KwhqFtaPzGt4L4YpmR2cugN
YI6dYkXSvrCXMZqPAdsEzcRRup9l6XmGWYNTr+rvlp2fT9K6CmvrFolrf1BTAr+Ouh5ecWw7XtZ9
+hyb4+YZUsoWJkhiDhtgRUdg7YMaXPQrqBe6ACoMcETJWLhU41aagAS4o+XKK2/ihXUoM7xN0G3d
2cfD2M3Db8W853FXeun5cSGUhP3U1HDo1krZRWJ8uDsnZIRu5sln7YI/0JabeNdzxsJjBAmlhhbD
rywZJT9zTdjg6wWKV/wevsVhago+HhMm66w1S+bymyNrJIuW5RrPd3GvcNGkQWb1QwHomg9KtDge
GZpXy9zWGwDbaZ+BDab6J6iMoaie75uRifdUKIgsB7/OJYYhUwBG3DeGqU0g84jGbz7aYFdxZI5y
qxyVkoOYrLBHKgUerDNt2KOYn1PVC4qeHrD7JpQx6jhOynY+yBDKp9+Eo9NEWt7q1YrfVI/tUw82
Wot3Jzh9plD2bKguT6rvZDssiipYsnaT9NM22ey+UHrU5BmHq9T++ylVb1qpHRvAyGPP06ScV9qb
K18goe2qviKQei54+wq5EtioyrxtVbDZoGhsWeSBPtYdfQu6hsPG8HPdEUL3IS4yCczXNU8ZBaMa
OcsF/UiT8CRJUCnkgvMz6FBCmWN149YEhN1w8WGmByUbkQ019EwqlyYpJBPd+ZuFewjQWZ/NIfY9
aisvEIqbt4j9FaJrl1+L7wTZk0IrUMs4Rt6Nyl9N+p2cilL+nT+ci9dL7iFKIuJCIAgcDHzBDFvT
OGVNQ3iD8ghILg4JtNsoNp3iMsN3/EnQmip5nSvy2fzl7OBSpwf9gHzUtGgc2TYwVV2VSpyYF9P8
ix5LN3dEVFfzQM0r3V0PJmSmKHGF7WAWitHSGi3iZ853ZzWTEtz0y9fKT0da1gJLjFP68CQQSrjd
UlBRaph8Vr2jPtktaaOkhbRnLgjeJ1Aj9uoK+7ntLPjYc2iKCdFtqi/8YVAzAEuMM1GmAc0qm7Ol
q2qoCuX+p9zkAAmNFWcwg611l8whnJzcRDGKc0avLXplYuUHgztLIom/+90mThBrrPhhPqtQKKue
hUfoB0pqorqJjmZfsP+SCVyJFMLYXXYKcVTRsPn9XpbL5N8pGm++eLkrG2VTm95qmRpKpjwEHGW5
FD5l2JmXzbF2zNOqXTQgbgcKIt0DfUVFZJVo0RhnerU5NveiKz7qNOwZvoaVSSjlJuFT0pQXYcN1
XvrbXKAlBHK3i+awTrdDZrNgJ906kbfYyra8pakCFx+2HBUEHX2fMcaRm0NgEzwxgSx1/dlxQiaS
mo+xizCf+hMtYpxYxddKO8FMaOXsUnue84TxUX3si+hlkhHVza6d4bp3EV0njIwnrPmlE/pSm/ay
HjxnVef6e1LNXl648mwWgy94tEWfDYrAF3QOFa+ZMRLuwIvzCwk8yBAL+rVd+Tyb0E93V868S8a9
YurEjbo1gHTfpt9R+0kIY+8zOL1pmlQuqm9Txkh47H2OAJglrOwEPy2OF/Hrmydobn9QySITcMEs
A6VeRKELsUbKghjn6K+GadJk2HTWfi4xE4nCjqvz4C7QGuVq2vn6Qn9vo7tP2OBWfsxevmqmeUkM
DpjkP3bhHBSk7ARaEgjGbzkRjX/p5do857Q6UuBW6zbD7NKGLl/b/cauvyGdaGtycyeNE9rZ3DN6
9RIkP7BUOQ3BkbUqMdpVoFjVcWLCsUb1VdbL8H1cNfK4Uw9fMEvZAUAtEJh2YYk/4F3xd4fwyugq
8JXrDaFqu29yk+Llp2Q5B1ZUUGutBEO2bXKA4UbfNCzXm70cZxHebghm6JxLGf2DqaWA+mjaaOni
oo4WGBTLSQn7kdbif5R3+oWpgbYNzOtfH6fGfojsp7a+tDAFMpt5eK7YH0adf6K49X23dlOHZnA1
sOsyB3rXUHUr712MvZ8KpNjCfFZEQQGnFkkHMaIVfVVvf6bvlDPFpv7ahwgo/p8uCek7Gra6BrEH
5gbpmm8uUFmpa+nOpFFDgRxieZF6yKvRLsA1z3s0WKTcIe3ybuzGBnagzGcWBOtT084JtyHoNEp1
LfKYhNNZTSoPvbxW2q/MmGuBaIFueulC4Gw6T2+w3mKdea1qy/gnaO8nGtIcTnssDK5pPG4Z4BYy
B6tFyb2smNaiWdd6wKe8pxmhkljLC4QZfLji2k8B7zUhdbzuXX4vfoMNOFoZ4FHY+TXEYAX7Zl3m
92eF6nwd9u9JuCVHOAVWl014AEPechvlFhqOkJY7DgFwlFG9O9EkFodLBww9RG2yR+N48dbM/yFg
/vvTsFfjEA65KvFmO7d2vUYp+GZsebpCO5j7Vr6iuoWf/kMt9oMDyBupMgb2CB0VakS0f1IYRHvq
Y9N86WQ5lFXSz9xayUQTNzfULZWvJn9BVv256vlaLW1ORr6KSwjF12ANZb/2qLMDEzslETeQEwM7
Ws5COWlQgaEUacwXVCeCXiecX/23ptzLGf0qf6VVyhsQldv6YUg98rvw68xXUzmXuxGPOeI4FWSh
tNwD1rRCZEC3I76aAmzD/Pqm+FJkXwKUL33CxNNS8XoioCIUVlfMexf6xn2PBker7j1Wo9NFVKbs
ziPx00BrLI6RYdXB4Kx/G/GKYWXKmoCE1JkrvBYTib/glsp6rS6260Fdb+yog+c5yVq4MvCz9cL7
5V3BAjFlLZbnN+7F6/UVLHOW2kAgkXFrIKeK8dtPH6VK89ect4GJYmaRz+T51ZzKQ3uPGr8hSdyf
Ken7rqGAmYYkF2Pxx/zQPrfcfw1SYQYsMpeJdo/PiahljYOJtrCzjhKt4V3m/9S/dtnDFbxMaTda
SvRpGgyg0MFL0b+pYPEGzQT56g5l9RghhWpeUs3iOX8t0JFTbHRnL26Q6Rj80o0PpJjAJFlhBC7s
jo2LD4zgbGDBCu+Yh+BFd9oEgR/uk0PoI8m69X0UVK/Ef5jRZ4WhjKNjdCZGDRUZBRkJxQN+tCn5
7UCHHT/qjgFYThRZHM3/0B0J1AEqZkz2MpsYsKCecIB5+ytfTBWUprw0SC5Uf9PF05J7cPzjvhTd
bAkuGOFwu97zw+g23BCvZG1MMtZukZwUehmzOxiPsEmpnqUTBeb/hsyDjbrVPBZFtZan6idZlR95
/51hP2d6j6g5vpWH43GMcUh9ILhJWfgkhSS9FJHrOwnu0cYuKvjmCw0O0vF7z++jl3ysaLA24zRy
7JRhDHawTJiU5cQYzJo8qbQuLcU0m65H+AywKZzCbVig7LrUxpC449RBBBQeMO35gq1/MFoxSUd9
WSWsUBihVfuNkylNt+Bk1zyo8Fn9buXTMTdJ6iplMwQ8G1wZt+EW8XEl8XmGwMumtCQsB3my3/BT
QCu3b8LefiLCDxiV1iZ2lptbp8goA4u1LgYcESfXTh5WvMYUmbjZ1Rh+FthjpyUnJocKPfVmTiif
Ym3uCu/h21k1nvsNEkbWieAWg4OuRdPsET41EjcpUz9DqHTerC2erGF+m86/DO3YK6DhX3DoE63h
xV0XceSTF3ixaVDgKEty2tMf0H0E4LOz/HTruJ1v7XD6N2OBYb5WoiBwZynvECYfX6tpkZaZaJFf
N7zAcnVECwvhu9oJ70qOUEboUjf5Jwsn9cCfPl+nrNSFmLlGCf+km9q2ak+q66yaxdk2FoK+8w+2
BRHGUhk+PFQ6frGA/UKbW55T4P09XSeMyj+ND7CQCixZFoKQskaZDWVD7TnrGUoy6d6stUWV2VFi
F0oB4rN5/jqUnWTy7f+J1cDImC/54GtoPJeFLulMahz27+s850Kn9Q/so75Cd6Dr7XGPaG4LFyx1
IqYzRDsAruGQz8LbgllRDemvLaR8e8Qr3zs0bmCMP+BL6yGQAbivs5yXL+Y0XNM8/LPRTkzglCOO
aQk915qWHrGtZyS8MLNsU2pKlRuG7a+dHzcjkuoT8/JJ225vC0ZiTb5x05eUGG323SozkZqckcHl
Wi4FOsg+7OVpOBsK9LbsG1jqWym5nAVj75pzucDY/vPMLaR28LnJZg3nXYDBRbvJPWcuAzLRTgWW
XOWyUWSyJMk+2+SE5OzXeRf2g93gfV+uknuxY51SYu3BBZtKdCVMnv/dvOrNJSzjMFQUMcPszoZ/
p6dyP64MXwxKvPW82hy2eAKFqAj2YU6/kb8gwn2ufe8re/enClV/yYQL4noSqwTCDsjXTR7tBKtr
uVjDRuJ+UpwR6OPF/TyztsvQqhPIc/mufrLW4GqUn1kqFLS7wpEgNKAN4wS8RvkXeBR7tlH7s5sc
jnZr8+GKPL7/n1l9zxl4mQUggqLIks4CIMUR3xOrwaam6kCM4K+IPL3yCpH5VrnZ4uA6CLXZX7DT
153lAQubNkJGEi24B/tJ/1sPKXUPQub1bFEGfxEr/tkdbOkfBO6zP08k8C6hdAnqQyznulYt+vQh
603yJ2ZTBQktQJ1A0VwDE+HWQBcJkKGQa2d6MkXXr9nFAv3ePFy8+04CqnJh3xImw7QQXR6ejzDK
xMKhql1Z0faEbh2+kuJclF9lGIXi3U6pQL+VD/GsQVqMJwbvv2J7GQy4Yb1Chun/alIxT+MtrjF0
JqUUXRL0/91ywiIHqJFOjZ0EoDJVybifRSub/Ki9UyY502Ss+UaUEWZUwCMBoDD3GZJZ9D9tw2dE
bBQdhDLdmZcE5z2jX/3yqU7md4WdzXuuQZB5QFIimApBtwDp5NmdKLlnIMT3Y6iF2vnQk7r3864/
dfFOiJuI3i6SeSS/USY3QkmsIB151sI2UBWiCBTDAm8S6+w7mnpn+vF2CRuISZAqCK1xsDEARYzl
ILmNctKrBZlPiv3HYo7+NssUbydSBckg3edyhSvPu6AThPmkqekyHwH/jhC5B3vrFTY6j8xBwe91
sSLRuHc97qw8lQBAOV6tSZxjomRmszKmOFvOPDcU9GskFlJZ5WS+iMiS16UP1rSLDswbzT+GrjUV
FBTMnKtuxEOUAGFZOl7upCQulVAQSZ+4dCxpEjr6GUzY5dw+hA2D8W9iQMLRyp8865+Is3IZUpml
rw/sgJUUzuA8hjB4IElZYcrUikL1FUY2gTCsKqr4zypAhMWG7v2DEWMVGh0L1B4EEJzbiJdl5ITP
4ZuaP9nZDUF5pUAzCAK+62kUaUZnKsl381BjhYhefeQXImSXmbV7FY4QxikqRWGdWzQJ25RWQZ+t
YsSVSvQLAY+62514QiQlxiheZQ4QEA9RDR4rc/DnznkFi+ACq5CiXOFOerfjjSwCp88KeWFRzuBA
NMy8SI801lo1cco9o4XTk4AYUs4zdsVlWHWI7zPg85McPatdIN2ohl3uT1KLwQ7qXO7y9L54jHLf
xRDPvNNntfYooq9UHbvJG3HzMk9WwJNxov2U1Yhz+ZQzpnVQ2NWQw+53agNPBOZtNx6d/78vNYSp
zqD6WmiZ+u8zP+Y6vxVhSlBA7rjWyE3goGqB8FAu3E5PNpzvZeTBXEXqgNFF38IbNzqxGpTQDpYM
+Ftk8yx4nS26p0Gd+PNDwmOULd0A8L3YNYSUHOsg2wGmSbqzlgjxl8fwLEfaobmBm5+ckEFRGvJV
PJo/9z6vUEYVQn1u1MaiFXITyOLWMtUQsHWkwhr5oCqwdpf7onViBfoMNHpR63gXzKaCnzC1rnZM
jXYJoJf+7LeDldjSaMoDMvU0mj1sIXQvUPgdj9/9RCDSaBUQSAuuDXn08WFPMfcwdaU0CEgiJThk
+7JwEN2NS6BGud0LLt1kHOISxxHxYVkK1FmxUyKcBQsFy1jTKqz+nYA6uXbAnoRGYbEosofvAQfX
K03j0O5YHl8JtnPrWyV3LQpC6vOYF5bylNM9O+YanDMbK7yFPWkdGMT4xs7YBhmS88IkPoFdMCB9
i/bydCvUX0q2KeiRY79lET8Y2hhtUO11LpNL6oyRUgFNbGXBJBjzfb6hNhtNI/HoWiGY9uKzz1G0
yir7J3F4FqkOelUgQNWs7D07PMtPtu8u0OOWx5/FFMN3yoXCrcUhseJts0J0AlRaZBX4T5auUF06
D9DHfjd6WU54Og335J6qljpxg+hpjrxscksYDpukNQwMv9NxJrxxWJvIVtSX6n12gjTEBQEDtthD
1rhyZQ5SeXHsA0qrNTUfFQ5WgG5K4x0IUCysH3AISyKo/kCxsZHcQ30iY2rRc6PAm39f0SlKY71e
5vdygri4LUySu+36nxjMcpnSDmGu6EeOWx0hMvuGOLHl+G63Lu/IFF6xQqdGoN8h48JEqe13HOc9
yro/zbbSTTOp/chbSOXIue6lPPR8fmYPlORXZHAunGbE+OfU3eP+sb42V4V+NXOJEjrZ3wfzdVzx
lg4/ENrVTLHGsQDzMpRNnal0469R9Bzfj54I0mBM/sgPPNwbGvN3AfP5RWEO+1WCd9o0bKR3XplU
Sg4wOubsA/bxzto2ow+qYoiIIJgPjhdNnfozeNVXHnnZBfQZay6byvoFCA7XX/ipxTLUm4kK5whh
zv5w3ZPcZh0LndcsPAar+dAZqygryhkElnMgwsA68+hl1SOZ3dvx3dzJwT6ythz4WkSsDQrbjW1l
MLCiAXVXY2q6zRgHovrWWDGSVcYN1xvFtsHdV9aE9Z+G81jGRH7J82wfUNJ/ofokqZYTHO2LrKHr
QP3oQWFXNLzKux34IH6qHvZ8ZUTdExm2wAinLyFDLW70+0gNTjmo6dnBWg2LM1ATsMY57MC2T4xR
ASulFNTiYAVSVuUq9E2sPHWboWHuYYPwoW1WM6ZxD3S03g77hIwGF7s13hJ7yvqlzEoLW3aFpf7W
3N15sJq0ctdo70chu1KuqKNG/kT1w/ZMHArLilT5dcBqPUFNpOh+bwxl9pgJR1DmWuGQfQ+GMBDe
IMPp/mpKQ27eKYl2ucMhph5SQhY63pVvmjEW0wXXjPMq0U4I0toW0MFVdi+xseQ6MowrgH3CuSyv
aGKE8tQ+PBthmLmDuiG9yxz5jdV7bqxao6T7y+z9Ejj4CKaTylIhot1vvOQ466w9azkQEV1vuwzq
a/bJdyLhsz4V8T3lMXx/RVy1h0RR6MgX7DaGjywNDMZzs/JFTmTxrD9/n7QVcK25E4pCiXWftbPb
ZLyKTDe68DmQ6AHQ/MYYjMV4MJBZaZSKCmydeJCxEvyX2UGBwbnQnGHhsd20GjNU8T8VmDYJhmLg
2TX23hX8+ZndcQsHxh22uK7V2bLIO7LSvG9QzYDUIJXLpK8Z6Sp1YW2DWclcB+F3jV95ghC+FLvo
Tv6qbJpynr5vlQRUio+mFys0/MBUe2oAXuyPCMnSlVLS36fwV6TbwSBaS0SmsitDfR/wPtg1hUCF
IxEJx7zLRZsq8g1Hpvia3uGsnMKZS05UHTr6sZUWMjy6TU4vHQzJBZZjrw6dqATIKyMWdf/lGCMI
zRNMlKHCYhGVKBLkLF0AAEMfSb08jihXV85Hpp3nsC5f9XypXFlk54NGts2TvYaAD7kHiH8DS9uK
VcxLQv9m7ZtpzWt2GPled7ULm8s7jGtKYrB4zTToD4+XE6wJLd9i5186vIBt1cJ6y4YYnnvVYdW0
MNfl8AoS4N4w0u5SCcl3Hp+Jp9lpuCVENTrIIudm4t/TZJncURY9wYkJu1juJEBSpWMVu6lJbVfC
wNL9c+4ROkXfbYNOel77xArffyzKyBh4yCTiumK9M4MwEs/gh6u65XK3wGscVjz64ltdUKXkz/oy
ZujNGDLANo8gB7CUlvHoDH2UX/8DZWwiWmA/Om1xVMxfO4rZGzMipCCSSEcpTbL7Bjzr+9ZIykHS
9Omg5I9BTLtpYQWklLrzDsFqkHtL6HM0S3Juu7Es29mMKm+JHkfor40z47KBEtmdE+mlUaU1CtTH
YMnU5JHKV5ulZgtdq39qU32mcdxRD5PEhqgBdmLlwUg8CyNwwv1cWWCNmKBDCvGL+IaX/1dtbiEj
7ppEXwkwPVQIGwQX13DQkarOhuWYBB30hlzhxDy7pTAUEnweSXO+V5LjuVWVcuytqZNZMEv3iHM8
/f33ZvmAJVaujCCrKoWYKt9us0zmfvYjAsHdx3xFAoP9Z3FhkdFrYWbeSqsdajABfV5FvMFvIZw9
0lgq3bM8l9vZ5K00GU4yLTDE6lnfVzIftOGp+CK377fz+a1uWvTrInn7PDaLL68GiEvt0ls1H5vj
MkqWewn3yJqBU+5TC/gEgp7b3IRQar5V0YjaqNUPGjtth7olzm4V9p2MheY6r3KzjsDnXSOPKRyv
0BzPFAqRdDTxqfTSg5uOgHXW5drPnhAOSmbiSH7AUckglMqUXVNM+oyAk+l61l3vcocxaYu9a6Yf
pXAEU/NyrXYlDrq2MnEkAQGYzHtt7ehvOuKDmScU8gC9gBDBJFcb3xhvYdAVyms/MltWErt0EHEU
yYiiVkoMRGV0WJY37Ci4ZzgGvFtvrkjtcHYMJRxmC6NkxC43eBzCx4fM9jVr8i0HlL4BC6nOIP2q
H35xUJSW2VF03yvJDqZ36vZlxDdW3qa+NCdR+s5Tq2ESopu0Vt58JbDkV30GMeuW1on3U44fvESc
V74nGKSEjjSr2BovadfXbb3zNoFvGXlm/4pT9grC4x6xRMzhszT++xe3IGtX/jCQm6tdVL56TlJ2
rsUVdIi9WnW/0Mb0UvUG/DsqDyoD+dDsNkzN8In6NSJuzzRUSllCwi/sl2cCN6c1akRXnsu7c894
rLFxDVHCtLmgp8ruZvhtWXE+rJeTOewE5fmDF+uWv0vuNV1weoa/OXZYw0GoiI05zXieIsFfH+aZ
gAznC4Ggbxp9RzduHy3MYARs8d9UsaRxHg2F8QKsCo/aKYbZm8oAEpvxNoi6U+nb0UvJHjxKK897
dcUn9f79ygvmZ64jbEjtnvdUurRlfebRPJJIGdDTRofwcp2NBQ3XNo/8xROd0cCPuJrGYZ0v9oTc
FtXVdx3OnMa4qHeBRU36z8Xjvm8v9GuTHIBhGY/r5PzauK3tlQl31YI0IO2cn6bWcmKe9WSdXKI3
+eYtwrJq9F2/yIxAwnGB6wNjeJTTqZj8W7sjyAV2C0by5sjSjEA9j9Ylq9CcOe+gc8NKOAFqrwWM
Ba0OqwYCNcpx7jYmdI6/IAcJf0/MyTw4DC/6BgBbXrhkxidMHMwoO2iazKuUErZLXcbF9BlGpIUh
TxTidgJrrix3/YKIQDsbsJ3QqOiDXGY26D0b1NM4srMd/NiSoQzsAAsgsv63Qb3vQL9W3DPATn0a
cHZrPsHp6r/JKNEOk6PPylkfWDxaBiOOmqkLVgNI8WhvLf7EoGYpwMqVE3kN+iIhsOKUNCj0L74R
zIS/Oyo6QIO8bTIZ0+QkCgiDufyRwYqUUYCflQtEQHB/10m+usL9IagcAiNMqumAQfVECBf4Gi+5
O5WEzJ6S6cuxC4U+LRmAlGdpAku7pnhg7W1gzOGD8Cn2ZZrc/vMnYunVePXFTP7u43CdjsUwUQMv
QYCCkC8hFGHShg4FpU4Gy9DjaDrubIa9WgUVFkljZn9BZRcQsJ6p11YWPwfyhLzjkhL0xq+cOvyJ
pudHynSUPQbIYwWgfoLBrno3J8GH8BoEtipMBTbz/gUYFoL3odqHq8gVpvdXkayVTZMmX7JXgUp6
Xye3wDsUAbhd7BxmXoYNzr0vt4kxTKSrUiukABkMzmnCtyYRykuVVLITaRCXDCK4JwtKIE03fmRq
SmSeVwbzNnSIQrSuZDaDlzw5XuMJc1/QxLl8ncvx20DS2e6EhshGWqbazAh4FXKf+W4lZwF4tkaM
BYy03V/8/ArbnnBswxYYquhCzs0HygGGFDd5bpS8H3A6CgqmLIecsat+diG7YbAEQqXJU2n3U/Lg
hcGvPtvGJhUyoFDFDDo3s/t4LspvVEnex0YkxVk1QVJpxguW+/jdl2zvY1u0aXznlAerQ7Plc9zH
/iHRaU3nfKP2JySqUppDJ7DDYzl4fWpya2S84v8g5ciM5p5VH5YlA5gj/PAPPVqCp9jGm7znOlu4
USS2hdqsNvfbNO+h5+OT34Fd0EadIeCwOXmbI7d+vKMfr7cVsnmmfD5gSeN6nsekBWaB5dFdSdJR
uQYJX3ZcuxKHafDEW11e0aoyZ5DmEHsoLJGSwlR+R4kKT+NrOsDKfGY/SqewEGiHQxBVq2bC5FO1
zPfxftOfWrtBDhTl+DwAU1To36GnRsW0w13NcyK+EqMImBvQ7m5t8/S7pFHqSII3dObD2/KRkFyF
GLOqykSYSvdqrBL6/j1AbxDBGt9Um7xIawx4rvjxh2jQ82Ap6l+UBLWjVbPnHNNaLGD0huqjLZQP
HoovHN+YyY+reM/twMxPmDjKjQjfK4BS5vgxg+HMl9Lv/ZKSlHD3d7dt9ZZAa++Ujkf6yW3lJzF9
fYdjzCFJccQjAhySZzL2ohL91PthghB5BUvpRhonZhdKMCC86bmjeEyUX+bzd/nhtVFzhxpk5scR
p7T+pho+lnzdf6FaO58ClBkhzJ0icUhZWO07HwOQgGa2nuzI0v/HA/GAxxCahStjyHcTR/jjB2aD
LolH/vBf2M4u5LN6BLO+VVQocp9JuzK7dvrn9priLDRuKT5wP0eGI0MGPnXdtF7FtOPlNmWZlmtz
HFqMCSKDW7p7aonrhmAxj5DP7BcJeJ04n5BwnrLg/DW1zCRFy6ZRbENvbhHF1e5/VV7OtQwYVRg4
WgCIEN7D3vqeQnGVNSMFHfoWRBss8YTOIkJjheQozgEXrCLag45/yOoFE+XsnblGg690g2WpJDA+
gp9p00ivZ0CsBUr4QleWz21qUovEoWywiGD4eLv9nHP6yK0OoiS8Q7iCgYXi3cbYRSA+2/Xml7AO
bggF+3XZY5kwO/CsT7B/2iOyW0lki7yartwZg+7SngaaoNuCkzbFfzvArsgy7hXl8mMfkHOKZAWk
D/hiBYP7Mc6yStwyWPEe3k7FTYRPSCBjr0eDVfLAHnmLS86mICZ1b2dLCNP0HV1kCof8so0rsBmg
lWoCUSemtqPVyjVvojAg3d2c8IOX1b6834gZJ8qQJUvMFa+mQAZmGseYw9OfNlQdNkHxKTkdSgvw
VYaeWVZVMNrgb1bJzWZRk/5Mc4RZczT8m/CJ2IUOmvIqAkiToiwq13HxtNedXamtbtRrzQoMxBlG
am7GYLXFWgXrwlI8u3AtVaTqbfktZPa0X07CXRgDMrmAtvSZr8ks9Xq+mraNJTS0iiT2Mmowfuqb
Fs6dkgzf3fRI4Qu9HKRt0JAMzLvSJQzsXrbMw2luyzJ4EZjcVuDQlpaybkuhxBkg8i+3MNKG+6dB
XlWbQ1vkKQ1CxaY297j+epILibCkUoVCeoTPg6gbBjFutFz2xvmXMX2a+FVmvNYwumu8jlC1jEbl
7XImvNDrJs7h8x1mrmoqsH8xu0Ydt9UlTH1b7X/egkxJxmydQkFtEOdMh3SpvMLPFoXSPBLM5vte
zjnN91ojJS9eeIQYPNNfyW6VAhMVCUcwg83jik8NY7p8w1jIp9HkdI4dqFivEEL5Jz4JiNK7XG2t
0GtlM/Xxm5sswy6mDmiPevD4mtK1/I5rpsDQE6CR9OPyakixFt0aBQlIRn6LFdr13JeZ0yQWuByb
vUF2ofkxcu8SsnM+6/97gDhUYRgLR9IIPw7D9L16wKUDengqb328aQEO8O2dEvF9ItOZw3L6YdH3
hu2K9XKP/b+GnjK0xjziYhPf0ooq4EsPZLDlFIn//2+vnXlV1s7q1ox+oZUWlnWY1Vf9dryy03w3
ukBNdsGmdlciS9jxmTzpQP83HUQREE0erIcbKq03AgRL1LeZwHv9fnijZlMCyM31/KGQaR4r7qvO
1WZWkhyWi8UxVd4iS5Fi/6Q7m5Nl774u+xU5ayYE4RXkGPcjzEQeiW434y4JLv7rx7PwOtFOLryV
ROhEE5iNlPaaG/M/a2ZKtbR83rG87AhOWonDA9DS9HCPTEzVeT2A2vIzDNOEbLAIjYc1XSCkjQgE
yJEcdXZ+4Y7OqxHYtRlqkELxt0LT1DyqvA2X4YEc3NJl3dldDFBPH6jwWXgjub53Rjxi7AVrmDKB
wLjt/j6+TR+Wh2qAUe7kK85J9HjQeH+HyyliLE5OHL84gV/OgH6ZXzt8frYI8i3Ruhrdf4grMpp8
S8NKplFs2sdtTTOFIBMc44ei7w9w8Eqz7OAT1k1ZpOWsbUfpNTz+vrEA7zSZHi7BljamnpI6HLew
jq6w3DyMqZoBWiT3sovUrDQ6lZKHcV+HRXe4T/xlpTR/CVuRZ//1D6nbs2u0gtcMx5OhgllkOP8W
r/lj1kQRTJnUcg8fkeUnGgA7oid3nZwSLTMxLwpqhEFV4QVLco0cDDsjQzL7yGwsc9lZmWHJN9GJ
0xr3hFkDi3Vo8TPByM3ypjJiEdge93MUxrtotUU1/Q0BZ4YzN3VuXNq0VyfU0R+r6sJjpWSsEKi+
ZaoPyCDcUb2O5HU7jwxqYOG2YBbGqiE5KkvVK329wGdWMSrNXCmilnQcMyDNw5N1YJOlqC+zhXRJ
+tj6oe7yyywdUlMD+WNafgHRWkUs0uUw49GQdQG1C8zmh6XkYLRG2UkTjuURR0ERR6L6SGI06pHx
kFsxmrXNua0uxyZiYBkgRsAmQsrS9WNIORc+bUKJQi1zSi3J8459eK2gzhpFsY5QIho9AbF59pq4
8YCm0ZHIg9KsFI/uria5KKia1vRSzU/wSFIdpdM/y6MeabrYFoshGhTOohgu/Z7Mb7GZ1oSvpvSm
7m5wAxyTxfw83bqIMFTZAM3CQ6YGtOlIHhfuZqjT352FCJ2Wwntn3l9ikHtfuhXAWZyIEgnTsZYe
pgr+7isFtOHIkTzF/4D//BPO7X2VKctVpl9QnHIFPJCVb5o9eBwUw5ao+SDd2JkBosOlwRnTHXCq
gK9YFiQN0y0cQpLpUXZyvJloG4MKtTviiMvcqD15S+FBKKFpVnCDlAn1QDgh53DWp/1WH76jVocO
MF1vC0Fj2fnZKgKmt6PDr395mKJKdE5UY3i3PR7aqgfIP4lJuUI6FdhjIZp7pUSArvuufuHytGXL
FFbCkFEpIYalKswDcOiPtlpTE8EnEqaVYLmY9otRckSIxyqAtv8ZUzNjVS7nxYwWtvtNyQR9OiUg
sMaN3vjRfih9VQhvIGqiOwDzxuDpUP8cdecWBRplyxwMtegAw8tAS/aIYsuuN6lUu8dQPmubi7c6
2kar/BsoFpCLed82HjrKKaeI+6PRAsSop3nXTnzC0w+zwNvtG2Y6TZAPP6bow6V2MHLxRwPMbnLO
B4mBcQYfBJZD/0Cdn0I0IGTpKqmrgSCRr5FVGB1ecFD/2j11UlQ9iL8pxK+bSuYtXO+IQ+54Ab+B
DjmePcwgVQGxI3rjC6PdHILtDit53uBTI62oU3B5/qDnD7dYMIfip6XQmSnOpDIGfFhvOfqqA/yb
xK6uyBHtcqTCEXDYkZHF1rgl4W5ZINP/gS3vygBW9CYzJsO7h8wmBYaSbKE7aLV54+DZIdi9V2Lx
FHs6IHOpFaJtg78hs7tPqNwfk7J+mEBmfikrJmjj+I4oz1q6ksaKZtLS0UrJDL2rlqqNDm7mi0OX
yM/94XVPovagyP3bh77dSiHY6dXg95iSeXP0pt2TVigIFCxa0yskTR9TiDm8vYg4cNTnUfon+8Cl
042h+U8Gouts8/NH7ZmW4BmqS68kCY4hUePX7aH5S5lxGBm1g9V6ja4GUaw7pbtIOL0eMWxOy+Ty
wYftaCKoNhvBCiwejMWD4FDHwSVUF0PSr2kQYlH1+wsM909PzJ7Pvk/u6VQDc6btJQk/AuiiUMkI
zMXbvUqC/7yQXB5u6pkXWj6eig1maEmP6AoqcdoYBcEX0FiWWfI+E9O5F3yYQ103hUnPf96sLEEo
4yD0Mzlh4Xn6QnuU/yiZha9dQWiSUNF1FglsVmUaTmnI1m6I20LXz6DsJOfHmE6Qa6BF6jSuG4Wf
oHCXw4wq3+uykPXJMIbOQ8XXn6rjrqRvMWM2hzVcEwuQ0vD2qk7UIqK43YgI03MLHE4wCbloTzm2
c6+3X76qgxyvXQlj9oMDoy1o7UMjOAL6uX5RwOk7MxuMKEXV64asjG1G0ZJxCwq+0hEwMpM7MQ2I
kYeqFpuaQP7aQzFfHGJZ8+Iu5L65vDeciZubHvYj7bQFoETU7EFw1AeIgcFPMG/K8ZofT8obsxv/
rcOb4scdYacDZRpLiRfplK1ZINki9FEoTS/eoCD4oThMU6dNerQanfaF4H/QACTWYTQ9sQdnSe58
KF2VUAD0WYM9pmjEtNwiQH7/ZIvY4agHSnC37ken5YF3pKI7Q3bI0Ga+bKaCslSmQBXQ53gXl7Wi
spp+aJ+yhDQ6cf6Las5xN4xunHdochM8ZVTHCoHylyhL4QMCsusgwPKUIzh1hYF8hyfMhNZYUzmo
vnXKJrbK8/JYVwFFNvF+sn8WuwHK5y+wDCad+H3RlyXgsp7k6x5d30r1m4B5emb5Ttws3mCIURPq
AXdZxjmR9INE22VoWfqOYfy0bwN+eMPqcE3mLSSLR195zpQcGriQEhdcNDgLOYQ3ftVSxJUwb5yY
/FQy3vJUc2QzYTB72DdY/xr/F+kHnugqHNV8jPU++1Q0ZOGjAX8VgQFLS3VCXiWwAd04xKNYclQ9
OF4fwFBw9rmlOeO6sFnGTsw1oAXf4Gg/t4go9Z+wFkekT5odT4qLBwK3PWpgJGeKrzTa2qyJTXoH
mZGXp2wQTb6Leg2QRstGcUTgiPtOG7ZVb0IaN0aZHZpyMKvUtAvKZdHfD4a0/mX72BTitARoqHA/
ArRpRY6jO6WVY7anjcXejdcjj7K45orhLe/3XQ24lzA9oSQi9vPGNyVH6j12ptpXtoFcpDpqTRuV
tC1N0WxJDuD7SR2GBlxUOeZpGEDRqReGOugvTLAOmahnD44goxl8PGc8+VXGgtU7BdnBdICankIP
wxrU6mqkhfytqz/dbYtOIMkEexWyxZN2xgqr2wYdpNby5pS8Z37Xi9ISQVg0yi+BnDVO9Ijfd2mb
zDaTqqwzANWG6UKLjSYb3BZbWu2u7d+dPYvdXO5OSAqY4a5dBv49LMLKeloG1rM3xbMGwBAz/5xm
QJkJcsLfdg7XmY/5vPBO0S5S5TLEMboHpCYVBpV5DhjdWLDsfCuAHzqcnTYYqzoQLqNu1QI3q8fQ
y1sRO9iqwUbLd377i6qjaKo44k/TAJipm6SohiZwQkJAjiFFKTGBNfL+khH8nkxVlsL6ZcOhyZB1
cFU9vBbv+xlcNJx1JrEkCJEBbF2JkPusnc8do1SHIWHowVOWZD3ZXXDVBu0gAGjcmXYzeFCG8M3T
NrET7GPUWw5KrhN5l5UqwELUputcsiLBpQfbNRmFd0PbDVnDr6EpGkbuakRSUV6X/UuTUuKFPnsX
b8aSs9cxB6JYcVLtfBAp7R1d81oxGcgm+HaHvAi6zqCOFo1c2PG6YwzcdIKqLi1HiCZOFRAZbWmg
JaP33ZEq8Gjk+tBFf6dnkqVqTWPU+PW0Jm+hNLKQb5hnV01hN6vUItJGow4qynHEQE3cjtSB284Z
2o1YR3iUweW6R9JscK+v4AtLemxSP2U1LqU3dJIxbBeb30M/NAuOm8/VOmtIoKvud+KZemS2IciL
+amTMu1z6sdKtHORrk0LE55R5VYMoLzldIK3VQ+oQX2lR2tBFKZNIpqMOBfCNT6XIt6q51oout+p
kszADKeXOO/PshjZEIpeLI7+qW+lWFik9+Iv0j4EcCqw18t0je88/LFZUxih6vx/KanowsSKjUOc
jdYY23UgtHiQFW+5eWEjYyNCVLCOuq3rc0jWgVtc6P2JVJVcvdx7cCZPzn1Pgcqe8YKfIH6M4gCe
mKMOTXPz5gkp9MJHj7w18GI1MBo62EPBEG4RJsncZL5XklumGXt0Ozl7ERKSeof4wDwweeRrJdi+
n/lfVKc/p1DxfpMSIeDb2Ke/2jw4XJ02M+fCuDO5vUiFwPb2/RKZmQBWtPvvG5WpyGTtvbMp90MR
EVzjX5NG7vw9poI3zZgG8TGzhFxdhvg7wiDgZ8wcSQlW6KeFekEyUXbN1yZEYHH8O6Lr18OJYosI
9EwE7Y6bLnVfoeXmjfGeCdXMiaO0QOor8z9eUG1WnbCLD5qnkUMOe6T9TRcjaezocKw0kc+BlgFt
kkdBkzNm2m6BGZ7+oWSl+KHgE3P/3uEwhB+xi7u0wh1rBMOm89gl2ObPUz7hv2T0nQepXjuJdzEb
K/XCfLh5+N26gPxvWt8AHK7AZ4VAOuz2Hmv6J6ntNqtt7InKBSLFtsbjdMvrtNL6m8LBsAzbhfmv
4u4vtiz09eq3LTHvQRUhzyKqbXrxoOp2oYSKMBToDFMe06RXa1WXB9T9xA3BkIY25eNmN47KbOQO
07kfM9ksqVpd3BWY+6o83vTgvvUSXYfsOmoQwsc93jlfQc4CnW2WlSF24FfM8IgNd3Anb4ldAVVl
pa0LOGE/7fhzbo0D98ewObw8WmwWE+90PbuSc+z8oiMn7ne5VcT/Wow0rXU7BiFTccHt+tRiMB+x
NOu+pjJwNLE9UKIS3lsiV4lnOkQZ0r5kp4AWXa4+pwjHHW1HhBgGJrfNtf5bnepHNejkYjmywEf1
erfljGGqWK4dXwfiZ68ayQCcil+1hRLtqZWBtmgDlMjRx+3bpumB/tVaeP2s0+5tUUJRVOH4SAQB
nWD7r84ClS8erb8E8105iFqQQVmyMc/bxJaShFTsBUlG7JUO0NDUZvemF8vnbtt8jP/k02flgylg
D9ItRZG+gkNYN+PVtA4LyGRYOU5VbUc9ID79mQ+dOQUyE2quZTQX3lW1joXtRxSlOcv4g/piRxGV
Np0ZB3L2kXrfBk2E8L/zuVicWJtNT46zIyUIcwlSq5m0BrnUNLkcQBEquPTlQlRo7H7jBUTHaq+n
meT/zEv6vVUj5X1DRckjr7AsU6DfYdHa2lWcET75Nh80a/omero9UUZPh8V3oN7ZC7JgzJU2NCUN
BLYXbGl2zXe4UBoNcvaKhW+nqnCyk3fgfFzXAUbwsiJHXiDolpsXEgd3/C2jxrn4xyfrjJC+w6OR
/b3o/Ehd8YHgfhijYLL+3n0730iwncfjjUNnYKmnWsBbmHkFN0UIxZKsRENJ0mTrNotkrBUoHMWg
aSuI+/x+PVkTE0rM1IaoL8cTzlgSxJM15+aXOWkqWz2nZXRpORwP7gINn9FwjQjZ+SANpqK0egCA
Haef+wLZsghvhv4m58MA/1fha0yTl92FvdkRNyXmsSWrhV9TAoKA7YsKWjl0e1cY1jLggQ2Vi21z
X1ml7qeCl6LxljOhSNO8Pr2WxrBqmLT+y7gxaiJ+ARel2ewqMeGqeacyhb5wvI5HvyPimuRh7/mX
TiE1gPwBmAh/AgWONDP3nEOKwsvObFKoIqHwlAJY6HdgswyuT9cegUp1KtbBtIJvdGXYknT/a+e4
/z9CNTO92BcXFlsc/B7jn2i2Hkbv93SVeEYBlbj6A9khkxzrCLoKdwPM0wrKN4HAineBSm62QOOA
rS6/TjXJapj/J/0BALPqiK7gK1eNW2H8EREQVbOO9A50Z83ni0Y45FH7jIG+7nllsT1qQuWg2uv6
tmvxz2dvlO9yNU4yNbuuSSCzqiM8crp3KOUsBURuo2x0ayTcTrUc4xi6+ft0p2n/GusD9oRmyY7B
UwhwX5Fhs/5iCKIrwYuSG48eB8Av4lQQ9eJN40k/PTC6FGzKi8BIbjGfMCaGZuldYrDkbypRx80u
1ZO4MehTI99he21Ow5IDGOOwDqDxIWm8WUG3qBQzXWUWkHUWZPxpVfep5hu8/A7kebJC06Wl/gY2
Hcow0x2xNZ8OFcj3DbtkV1LCLJWJAF4ZI7soX2UUnMhJeiIVqqyPsqxrjKt4t+/VUrafrFPAo7zo
yN9baRz8sDmcN0eOkaPMjTV9Y2Rh/wEGxrYBxVx2SUCmmfpa2fe3b8jkTA9uu3gKU45ROmex5Hll
m8MMMBb8di1X8+yntV4pLOadXHhcCK5yKH7rmrR3Ypd2EhsuMbODtcAv8o1y9RM14MKxHHuRARjS
TFfbQRJNx5TB6BYgrpHbVgMxSPVpgHWNWSTG2lsYUde1t0sVYblisWdhKYyXiDA8CwSyLSvksucL
tqaVw9arZjCfzUpFjVyExnq8iwyKt5RIIOup/8eXK19ucFOutsUc+Q2Lc5uEqP8yABPZoiBXU/MP
xK+9oWQ2DSzre1MZ7TR7uhYsn+XUeid1+hhZBf6qCH3+YXauM8XP5G64iwleCikkUbxqR/KDtx1h
CIH0suYwD0LqaCiTQrrvc5Mc4MvaTQay2LKQXp8iAmPl6q9VY5Wj0ApFnq7tNooq+hOYc7ZiqGYa
aeHZR2S6kq1YvAKGpY4Njeudg7IajYuGshEpi4Mj94GR48raVViQqfeCiEBuVJrqIbmAYJQ8GT90
27oAlLtclGXUrzNYmMCMRt/pjgvriLO+XXtKjd0frJJPfXjExxJC0/COT0SBhpF1XxC1ijeGVxMz
B+k3XMEjgrmf/u4ZpfhC33KNIR3HrIdO4/K1TxnZw0KrVHrVzsnVKHkcbqzrAqyvyj3dm8rLl/3R
3tQbpcupcsNqkDhrz+07csATeaMAeUT5+CQFy3JB8De/zp3XqBguDn2PVfI4LYQX7g4W9ttpZQCE
sx7Z24576635seMYc4Tndirw3K/gTa/BMEX4/hRpARz+PfkncE6miTG1/Uu0xhisk76l06Asw+2U
YOmUE4FGz/sSOQEH3VwWmme+f815HeRFliQs0uBCTIRMyA/6qcVPqraLN+9YQPEFkkQcZpqtUuk+
/IrnsdId69ToIM+OzpgHNe90NCajkW+uHzB8LJrwoJzN/RcsRK9S8DX+OjU+Kphr6b0FZhNKEe+S
RBKubrkCPAxOwoODn2ljPu+XLkYPEYz+14PSPbwUjUHH5Txt6Sw8o2pDpqM/q3UREcJ2oZ8BeOsM
4rXM7bdsxQBiyBOQ+5ETFf6bz8LOxcpvyes7RArN12WzKEMWJfLFkICj4LBB4pOIsbhKyiXGBq/2
sS263EM0nkclI+BuOa15BfPMi+xKze8t7Tdkdp4M++CtIH4RG+bA7mIX98YcprZf8fc4bJVTwFMd
iH4CBrIhhSDhhKHvM9OoVfr//fo1RoL/MjmqKYI/7HaK0i9DxZ+of8k78ljco9xlK29/t7EJ1ni2
BfhJOaJLeH2kbprG6RkmJsCdbvu8/8anJVTnWWOleD6NUNmyukJlnXf5aXYrLHdO755xxwoH6dnT
2k+K3UO8wIs8GrLA0M4igM3Ruy44XHHC60FHlA9kaHH9kPVZOi2PDTJs/z1TDQxhRlVOg+H658bE
jivDqMa2X4Jbtlk19Tsmghf+jKqlYNfT8slf45HkVPktTF/03qYaWzM30H0hUraheDQnHWdOu5hU
Bji4ib5SyLDhzCxRas6UQDOZ29gMeM9XPjwmlusMH9iHo/Yn3y8iiT23uSZzv8ifoa+KdFBR1Hi6
c0rq84YtxBEh1/xiiBJ7TQcsjd4MpBYVvQh7AIxWd+zmTd2Hdn8XdZVB4ctNqsCjC1J+E9ujlQFt
170IAngEJqggQXnj8TRqDP4VpPVISN4rdnfBXkpx5SKcrlDMp8dlN3T42wKZesUMe9r+J9BFac47
mnyHsX/pJIpyWUpPXz/UlDShB1OqQLMwPRavinCu/YPm6mU1F/PGuQPToANsMMW1M18WMNhg0YF8
a3h8gjoyx/MJR6VPXqCYZd0DKTcbXZNfMNSfxUXPArfnab0MPKTHRS9i86hTgST5nbDeUa8mPCdc
1uvdlWzNDBaYs93bAZ4DJwzIVJctKYdu9D83gHj/JsVyCSegUekha2nJAZFVtGlRo/j5dNBfWa7x
J7k0gnb3PPobtlC3JBbut3+qHt9JS5KuCl+okOWmb2sS7l+Jv7pbfpflc6f3PETt5emUxmndzH5O
OBe6r1LzkrtXUGy8SxlBkoVU3n1CMA7ATvr5vIj+IJX0BkEkFbuw9XFy3EFh1yrDbQfK5LEXeqj+
FXwWvWff0HD5Zhre6OGa/Wb4qF+7IMczTgnQi1nSuQv46VXqBXjts3hNcvsoDOuyEAh6gIQoFH5Y
vP8DdzG2oF8tnFQAeUzzgPP6PcpaNctfLUjIRAcNiGZZAv4l+jGUUXgF8Q7uJlYua4XjfmhrNLXS
s5yEylw6uIMbaAC0OacDLZxt3nFLB9dQ6xMquDmZrnBpFmIZRGD6A5INPBVrlMFPSUVd6XU8vfPN
14MjwW4kxEHKZfxfaz2o7+REu5mrwtVq9avn0BNMlbbCb3GHDPfdO0E3M76YXIUiknscE9xjzCsv
cEYSQuVihziYQOfC5qntnV/1QFHr06tlSE7JELWDXSvbuRU25dKrAOyFEz8R/el4aGm9Iy1Gwmg9
Su8C7QzxcgUe3gBLAtYtHSpASj5nnYNkxiBoMYVW2K9y9ixOoLvCILQ7fUKlICXSodYOPfC+vkDE
YKL5HN8rxN+B9wK/0BUeqtD+oEGNKvhEVplIqYsARCR+EbIQcM9MCsI1nqV3afjPxtyDut+1QJxK
LOuuRWSIiG2md6aurwj2xdPJiYt2RYUijGbdqtBq+DROIHLawZDzQpwI9iMwDDumMjSNUemDmbMj
sAUiMMRxBp/PUxEQusb9BysZLt4v7jSvpaE0zh231ub71yoUXbXYVF6c0XniyBYf5weo42pDg1Fx
72MWywyIonFEVczHbCq1Z4UFeBzS2teuLukJ04XvVb/6XDxdCyGZ88lHYTOfFaxFwxmrb0ZVcVyM
69agMXTXXL4CQlX2fjUXU3dbym2nZ8we0ebHpSOdyl7mEzAI8pgT2WI5cAN+m3eFwEKafClZGVDu
CVom+XtFc3ETy4ulNKzl/FCSY1rdckVhljLDsw0Oyzhp7cMHJ7UWCOg5gxC0Nl8r8LB/9449s21V
CSE68GYh5khemZlFyI085sWf3hOaClQWJ9EDzKqLwZb/G7DsJNp7ulwl1XS8RMqNZ4jmOYUCKvvt
0IcBHI99NcMeUox90BnacIlUmVXwz4wzZuMWI3ygQS9rtuF7esl2IWGPgCA0oB51LcbAdMVnDyPC
wBaIHm7679lh279TIIA8lTItVpj9fotsxXCLB4MrR1h3Op2ETR5dtUvwbM9VhK089NaH+Yw6qFqk
wE361ns91grIPHk2a7JsnyTe/OOh1VDKaQYI8BxB3eW0F3GTotYfV5hu4gbjcqI6V/a5Ebskw4Un
SWoBDEHxt+Egxvfv3oGrWy2X5otHZhvzl9jrcmz9LNaPMg+se+Mue+joXMNoWtg+RaTJU0E+q/2L
lwwsmaUO+KkO9mffPEmsACPM+gWIDvpLmwPKxDF6VH1zk5+5rqX78C9O0HZ0Wy0w/BLY3KOWmpzY
YLyPnb57oOIbFIg/cEQLpvn8jeCZekddk4dmR5bkIngAeC/7aG2Es6vTmUI4B6cjSHGvrx60GSwi
39qc7hBoZjGdunTxZP8puJabSDV4cS6sYsgn/bfTjbbLAJlunc88EPds8e1aYiD+SPAalrJQsVM3
3gOSA+GvnjSHykpQhLKh0HSNpq7NkrFeNT/aK/bhq7qo+W3zKojP4V7UXioBZOv7ZI8aF/WDFGPX
rYbF2gRA9Wa5gFX+EWnZgPAxoEWxTpZ/aBQIoSYjuJrvj5PY8jGah/zMi6Nco5OfJmIRtx95NnrI
vjjFfA8mA3VsKNCyiRq76+g98CpsvxwqPXR96JZwzTF0JR6iBjuydXOaJ3LICjuFt0YsF2P1u0HV
YObRdaJz2ylIOc5jq09d7UxSyL5nWR3/g4tY7Mt0yudlH+7wvWxiq1B+NYzWbiaPqnp6eBhNAB5+
YAH4JcWXi6m0ZNyeV7AEryTctYEo+bjZN/cBKGfUFxIw8Bgdrfliri4UVN9pLBRhjhEAbIvxqk5a
btYBNI5UVuKwZEE/TV8wKZtagnHcGFm3K8SrcdklRIaRp23myDIIdY0OjhXB4i95W0t4+wkODyKt
y6imVjTs2+DPBXf4PAwnGbE+1QWUnB9CiQBHgnwz8pxuHglm6K2OOIO+UXZkkEDJPJbZ73MnY8Qu
suX87BqtC4S3vncodpF0sXuxUUUkMpRcN6Aj/dJnJsRM26aOqD7zrntlC2W0T86/gOHZ/rQ6lXys
GUwNFva65h6LQ/Hm2OJsTCnWvAdHGlI/r+7jyYd++CZCMg9EoeEO3M6WjM4kLDsBGz3lmXYHCgN6
OqUr5m6e76X6ek/2ACuLS2uNumEwYdmCESwziOhtwnA+xsSJvEiDUbS3Mc8yKRFkd59WphEACoNJ
+sTQuPQp3UaYYEj91RyT+Fy57TWrkUq1nt9bvstu3QZtN687FKzREy/IbXRsa76K8Go1budzhdFH
Lvtlptb0kQsWyIqr0KAnrnl8GGw8be144Q0eFiqfa2S4Lkw8Cc6C4Eg0wjs91cUlg5pi8pvkwbXC
4DzVXHkrd4LPxnzWAQjrL9eujVbgt5C9lfZa00yychEERt+qWiOtblhFbwe7dWpUBnzaW2JZAXbO
LgAUFmCDGFyB7aJN3Rccg/yHEcBY12ps8gCBn56OqJDa6HsPiTe6XWuNPD8CMSnNvGg1LKvWfQ76
Z0v749UAKvkp/yba4n5RdG83hHUSdRxHhCxnk7cJxsUgdaKeG9M6+1XOFlHIsE6RcLtMeVvHfgZ3
52OOuWempEKIoEv3hVjzYm1KDPDO5ng0ryjY6GXkIucbTJutZqrOXFlpVqy1R5GM8Y69jsObYrC0
a9i5d8ZuBnWEt9HAb1f3BnPhIXtS0k2QHrN9fMrxjdil1IVgXsNfrBMtV5O676xN28t2qNVAHAts
kvEJzd7gwlzMwbK0omO3PsMOFVlj+asSVBfuYe442Crg+rUPahXdhRXqqCj/7fumUNBEZ4gaafgN
0vYKpmjAgTQhuS7q6ya4UBy38Oslw4GREAjGY4hMb6YcFWi9ZuzdcQNrc1JmcwELdMnsqHebciXF
ntzVlg0hP4Z4bGhNzxW8kvxHXUF0L6Qe3J9XqE9eUDSdnNpGq5bEfBBFSvO2MnIVl7jwatFDnS0f
xrATwgo0Nekwt8tQNMXusIyRUPIjST+Cp+IOpVreelpVi4roCkrH/s9YdVKdsIgx9HcEAg+hOE8l
IF8/8RJhbtlFjGkImEadXe6gX8GNJG2bnt3/vL79/TqNNzY9/QNbb8AgjXDhmrVs5DYxhVCp4xUG
Ot5xJOboO65Pr1vTakLiS+9z8WDLH9uGEVwttdoOsOJ1hsp7ZboH/VeUMq4VAOMfLPAh3gfI/Qe/
t+HIE9uYG4m+UR4tdtFn/0SVWO9mcNqhjz5WnGjhrnRg8Tgf8bW4ysZJhI5t6EOlzr+smxgEXHdf
ZGX1uWf3n+vI4tnPxwIZepsB46vKOP4CMyrHguvF1TI+Ke4pwIw50uA1w2gmukO8oRFpF/94UbAe
jVZJcI9H6IUOe4Eo1aqiIyxgREpdCo1aiHh377zOJg0eZnWAYoj7IR+X+Od1Ncznx67xp1zWjl9M
IzmdqNPbJcNQItODQ1fOr5dgFTYTl3czunQVLZDJsPCm3LyayjSN+57cB6D+L2D0DOX8Wz5X/LDZ
go68dFwNGrSkQy42cmOBaklOYjOxad9x7Wpy+qUBv5qQY+48MpN3+yWlaW3ewpPzCbtb//wMftqu
t3g3K9FCDLXXWU99o555DdJTlB3UEhwKtkpj1Yh+heFk9+M1PwCex/jY/knXrMbgxKM8JFg0ceUp
yMycXJbNurfEAJaKyDHHEyrh5r7xVUqOZoMKMgYJpZ7b9rDuRehJneVnpA6gj3WkUjbwYLTkeAUO
IUiVXXfG/k3QAVbk3ecqX8k9/uZ5MeFurMx42Pno/11vFCOgX2hh8ge8sMGWuzXixcTDLrZm3INY
aomzLGP8hLhAd+KeEqRH5nP0hwR9zZWjvAp82AUn9z6vWXBO0RlQc75wdFrA6aiHK6B8WFF7sVOK
VLMaDvO0U6cUPefdrANGzgMlIzgkJaYU2kCi4SrwLDtWgJ9rQRBXXoJB4I8pSgS5F3yXLRy1siom
G5/cbazlPkUo7ioLv3YovJQPC3jmQfowubZbVeHZO7XpYzprKrp/CtuNKsjirbOreeJJRavKwuTL
f1KkKNLqgW4gaoihm54cHN9bGYNjszf3snxptB69VXpP1WkCRD3NJUqrsHGmyVqMY4LVKlrGQ4Or
M6rXaTqEuKa/umdRr4yxD2pZYv4+avonWrvYrwfn8rrnMkoBkfoOpJc+Yw/vsB7CPvOd9R42tqo1
c/WtRAzPPSuYTanyZ4GPERec2J55EyMKHEcv7tsLmsQSYMCl9a98+bJZ0KJxWEVU7f8s6kUQukPs
ahfsUAaD5Vd6dtG/dV9kQdSGYReMBaI+jcdhN0P5C7fvTG7W3xUugI6R8hOoXsPB2kT4l22ggr7x
TRd1+YhDWWW6wKc+DsOHWXZUsp68pavkUwDaWfb/5Q5SsNyottIj9WJL3C2KIaFQ8DVsOruEtRci
VqzLk8ll756zuLnjlPHsrbhQUyepRRb9je8UTXby39C89gNG/ujmvxxg5VpZA+zo3OJpBM9SvMw1
wCkuLh2AVlTcLg9nR8qmrylthKwO1YqMLYSuvBIS9aXwcAJMGoTFgpywLb4p1XpCXzAExc36EsLL
+ZzcpEnG1FgqyzK1Yiu8tTMebjY065+EIv/9YfCJ6Agv836f6ufIWjXISvQ8Pl/gy4Cfu1kfqRYz
e46lJU9ozLehvWZM302OC8xiWeuR9XORVMbxIaC1NWFofd8DjTe4eUMen1rr5lAegSCAcFvIKJy0
FCo6QwVPcVG5AM3kPxyBOx+DQiCwnXRSieyqUJ/kgVOQLtDgQspm/M4WH8zlIMOObd7JoP3ZAzpP
cc5rGWjw0HhRbScs/07YgpEae/OwfaKG0ivA3ZuCea6kFrpGNnSVCsjAmWNFXjfuSvj2YOxP6S7F
S8G5kj3EfFwp9saLYESL2Mzc5zd6/lFBAZd+Pgk53oXERoB1RG1vaO2Q3SXsVpQmg/NWfYXH+8VR
xav0jt0LZdGUR5rjLAw5iU4OP5Roc2H3pTvAQz9W81t/VFGng4j2zprebdG/nvCwgITRDbo0ZXQI
LxkM5CM2R04cWFnt87kmHIDwSxT44+/Wz0j1YOb/FEbptXzO6MfES9zmPBvTG2YjR23DT4hIfKXD
8HE7GJf0yvw18xgVs2wJWsWPkSUdgsT1Hf9XPQUSHzDffK6YQXhiO4ZjYjYW0+8WaMMDZk+ZfpOU
xpWkCOan+4ksFPUZXxvcpO8Wt3WaJ8fsiss8RsQTFk5eWztA2GuHUZY3X51kjlHTVfhukn+LiiB7
mL2dZaBIcf179Nl8jDO5+c2jzqELm5V8kXc+J9K5ho99z2GNDINgclNG29ALBwBE6bOTQF5eLAcF
ISQR3ucGAj4MLiRd/H+QkeXHNrdf6K84+9TGsmUOPSR5GLAcph5uf3MuBo8+L5K66Fh07VVDqKWD
H0pJ7nusDh+wT4Z2aXwyttM8HR+FGmku8M+j/Op8Gh/EkQtDyj9LgLPle7c8PCWhx5RjZz0+ZpU9
3tUgEgxPS1N6mIvSM4unhCV7RXiO5bn+/0gUOMaVqawqmNyGMCDNcNvpwtBY1KEZyVZVHBOfzkRp
9CM10CMWZidhPoUcAXa03DEjume11qoljItDo6geNJOLTe+ZT/Eax6/mdov84wysHXdZhaErKB8E
eHxL1REfCF4OxsJ7+hBvezZ9U5AJ/dGeV4JHbiC4B5ilXBCqoqHvYoqS0ZfeA5imq6XXfD9xIBFO
GI9Zjdg7mG2sQlh8BDvIE9kax7eC5QqjEe+YpW+kyjOvY2BfGye8q5fYcW/+x2lLFcPzMqEaw0gr
toNNdERiRvEFnl7Tlr3D1Y82og/9zRzXWbod3KyOyE1YK24+mwiSW5T/k8PCIYUxLgfht5bN6LsR
mJWkX5OAgIVY5W3g5u8k4m34f9YT/KPlTUQWimq5CTa3KTpc89jNBhBgmYZO0C2WTcCDKJFvTvPV
leG88H2yI8ZQQT+lAfISTGO8ohmdddlXT2L6j940rH1aLmY9El8e+MWlMkf3B7HvBCiSZsCIl3Ei
ylIAjAznTxfAXu8wch+DTsUdoZissd+iCLMPyOZbPFcMC+WYCrUGLd3wFPP6AGS3xfc5U8gM9D1C
IxXqbL3TCRwRi6aZPh/ogyhWXqWJaZVhWWySK53IVv+6pEWOtOudLRxdwzbiKfBC6mmYfGluOQSr
FJse/ywwoAg5nbA+F+BZRPQzBXHIv+yU6aRIGlfmpmDJ+IDYSP3DStjFav2K+wHjcXgFFve+aqJB
A3BqbmaxEwaKhpIam5XaRJWkkFg0pIIr1LI2HqA6NN92jY5mf8zjjdBNcltTi2JUO4p+dsS0oVcm
oMahw+DrSGQhr+8iLdaRs2XdYoRVb8tngimd22MuRH/flwmde02rdqk77JBgEGUFfY3l2g8EYqPs
jgN7FejFCwBL9yFBMn33/w6zlZMqZqG4vBcpn11SRzc1PG41oOMHWJvDP7FBpYv4rWUbhxGNR95S
ABvkekYhcehM91UKwgX1/09is4K0Ue8bwoFWHAkw8rfWquVth1SAoyw2gF9ucDnoLLnEwwpQa/2M
N47iq4HXbI4ZJJ2ESqDS9LKaCEngG2ZOUrsiWH12xGbl+H5Nll3xxv+/Zo/bZOjnbRC+HS914P/D
U31FLKlVqjZMlicQEZ7xrmcQFKLtUhCm52TJ3P8efyR/bmWuYNjl6WvcWZpQXYZFmXOhtJ/wLnfD
A192nvGLTsetw6pYGWNYm1diMg9xsJcvtuSni1XxsjQ6Q99XXzb4XpsCDyTrLklraygoa6Fi/9Ge
DG+xe3fnFflOq0wOG5/DxYQh0BuO1Ic+zuO82Gg6duTdKArlpKlxES+CuZz0Ji4oK39twuHrS+ET
CccyynEg1zwRfb5oJekGs+d/vDYsY3CDKzKUYWmNNOofX34WXhX24MX16N7GuFKl28CVgkkUGKKh
Sa7QHK5rDgMWpWfkAqWDBuF4AFGr2XPrelV2gH15C6BUBjlXQjgd/PE9y9TbPHdjUougz5HiKA6D
EQWp75JZ/z1KtLMJn4RiyEK+X96lQzC8dmbxf8pzl3JAGGh7Wf7R1Co2OdtOkUg06h5EZinvrE9N
PGMoOUfpcClWkB0eKdBMJFUIhyxPfJWx4+eZNP2KQiFxXxFkqyQ8ROyhZ00aou2Hg1Mh0jRpAv3V
bO/6FHZTAk2Dd0PAf+XzTEhIOZklH2xEB5mvsFckGUq0z/KcZhREqA+JvktyRHCU0E/+QgoI0GgV
LtL+Jgl+AD9VCxlgKqfKqfq+uT7bWHwfcfquLhXf+michLl6wRkgP+9y45/faJT3LpP11PWNMfKa
3+6h8Yt3HZUxVpZBqEHoCr95oT+j1uRMIT6RAw905EYvUxAx1QjUC2eZJJcUxHNPJ3myQc1m/4BX
5jbgBwFjUwg2ghdOvQcmS0SSeSp5Vebe9KoeWFO/dEHnzrrwkHOrlwUo+cyxClgueyhuQUPlahOI
HEyzNnOuFqzoxwVaDr29DgZviAVK4jJko+5zQbwpZRYEDv/RkYh0zcKcCplsIuNe41YBrm8WPtip
ADdK8ArKUY8ebNBQXK8DiYd8oxG5++aJqUJI5iF3KNT4yJPiUT2NQ9YAfOZxOA5rm6QqwH7hnsTL
Robq8Yjm3ksI613aT8mvsvRt4VUQIkl1UXcGlayF8RjZGCcjJqBwungIiR3MjZxW9dxywNFa7dzj
NAQw+RcwZL8s5lkq+XtvietQp3IsZUu6BANNeNplCVvHK81DddaWmWhBVZ/dFqhZkuiYlMLaDskx
03xvBVBKsEciSPaflH3OOOPXMhSJRmqf+HhxDQwK12GuOMp58u3kTPHFkJUlS4MWhePbYkqBEwwg
iuWpBxBqfltTIgGOY922yxf8+NqdImqBtao0PuecN7G1JfXSTHCqoF54GCkPdI6AbWfFE53MyKjD
78dDS7USmgKFv6BiGXC9TvygaiqdmC2bSzGCCC5ccSp2SExX2zQFiOwLxgRzAv40gW9XHEKVNAHf
Qdnhmr6jCqz4L8nmpXld3JVcJNVYhHRyQK2Ljkq0C9R47xxEaPwvxb3ZPY+dpCrs0U0FbbizZocB
mfZqmIrjSNN4Rm3NokRNQDTgWjg9Z/Q+heq6yM5/QfnmfIdCfv87SBaTjKc2XOi92tgANuPwYvR7
HfzttYhFbsC/iRHbDtAalg7ypNmdlIsgSKRaAN+gIGa1zjznwhw1OHSsu07Kkgyn/O1d9HrV2Si1
62oc4fRdPI1TmqJ8sFR/5G9E3BwT+n967OSa0wZCu6Buy1b0qGhHAt6ToTmfXeEfRjzSn2Y/PX+9
ZtGj/92nSU61TbQRfFNEfBJDjEmYAvOuvJ5i3KUQ6jLGDpoMC2N3D0RGEgFUJWDArXIks/GNTq9S
74KsI25u9XfWpx86qSmQnC4g6bGEQoPhUnjEOwnRee+b/CuGCmqWcZil9L4gb5+Fg2d3sBboIjjN
Cn0gwn3wcHpRHmKpSFDn3hirl3YWnzypbLz0HFWUV8SxHM6xvs2qx1IcARtU7kC1G2o8LXlXc1i0
sacIy62IA98Bd7M/k2I8UDTP3k+UR09MNv/S+vBAWRjhEO0BQRCKydJ6GLGnefLS8mjTdlMQBeUV
EXxQ5pN+kz8CvjW/UpLyyXd+Ggp+KMy1nOhOB/YLo7K73t4r4AsTuAMB7q5fCInSY4nzC9E+szZC
9xzqzUR7K4wITK86fKWSgGIIIPclTtCSYNkmZkmuuvDuzzSdxu96cwGf62xlIV4ln5xp6KBMQEwZ
Vk6r1DsN0bgArQY7qeOrYukWGFOBg+dckDKNSD1y5yI9R2kxQOkYwkcC/UNGkpyIhtRK1i+0ledV
/4BAsqKXhP0e01Fo9HdfiKLFTihmxT8QdIkoCZVFYtm+TJUEs5UDhn4FzhyE7vrIk007oZlWrjhK
y6HAOLQfArfrfDkcQ4sgf96PzgwRMhuER50iQGpozewQCNV8GwT+EjT2TVrXG7TIQYCfWXM4wJ4Z
2A3a4sVRnmQn/FmXNWnP/Z7HQHY02yXJWFHss2210Te26AI8U/9cl2PkTB21Em4rbLVnw0t5rB7i
mNAcZOV4SaVTTQFmAmjRyOIYRb/lODiDGjoVHe35VdmY9sgtbCLopumNB/+9Z7M6ZvqKu78/1yZh
9BJiXOI2tnyY6O5ps0gskGybpdmFjcLKUuYcjSwGH8F/q+sVSf7AUTtigx5AMFgfs9J+g5yOCVMR
dK2J1MYK3TO+oTFrTeY0DeNQlkZcD8qz1sI8joa4Oc7pIS6RuA5L/P8kDNPmTrGqlM3SYQUOc/UU
eBSss/C91JZKBfZZJc+P1qBw6t7/Eh13RPDdpN+A8FXx4eCsHETpxWMVyh4uMsF/gTDMBpUg/VhT
8zmwBrq/8cF4cFsBLHlskPK8emqhZbgSVC+EcE4GvpCrDYF4sznW2spKvamCANWe0lTnrmy9lvpg
HKn+ejdplAsu4XOtQ4RczL6v4qd3mJlRVZI8Qz/oCpz2oFLT9z7G22rfeUW29yC7f5ziZWzawIZI
xLXzgSrjb/YK13CbYw1r0vTYgSTjvYPnDCsbM39j5M5pNOlhMbd4M4JVyPLjI/Zo7q1WMhbcJU1N
9NLmlYxCmNTEGlCFNA72I5Xm6m/RaaDcmKTtbhQIu2UxDXOIvFy5vlmQtW9KcqZbJkaqxH16V2KP
wQJ9kpGwgRlZWFN5koCb19FRsnznq6TbBg1QdfzBazIhIGvaBLzJosVI1Iz+v4hakLunW/CwbxUp
nafZXHyfClDQ2MhcKSAeQYS0kvz1bfQ7Eevswr1+LvVr1KkxHyGxhQ8QeUvg9/+j1hLQEf720fAE
a3zRonnNugEJYMxjoqmhl5GAz4W6SBGvibzyrd/anPigL2BA+Eo9rmiiwAPXCHQACh2AeQXGbloq
zn50YalFPtHauJDv+etDuofG45a6UgNEFkOpn1j4cFxqMcu68xX0MyVLZvSJmTVEcAi0xE1Xbdkc
4rnj1VlP9pFWlToy8kZu2owpZIMZR/bGGW3fHCZSu1fyvvsIXuzICedoS6sxDrwXe6EgcdAc5ShA
0QH1bPE0p69rvbbjU3ybDokw82QD3LShnaqT4eAd3/HV4ZHi/vDWhIPU9aISun13h84vWEhA7me6
RzNHoim0J3EgIaWcWrJmCikqwWyvMJ65kBGn4ujxFEwn92bgvwlbLphIOwK36TFaFaVUXMuCIS12
E8m6bUmMODeyq9yZTiubBINUShFSF5ZEN6cr89c4TyVr3uYvuYvNDy72cMA58VqtTVG1XsjjhjBJ
8sdrVQnuzipde+G5TX1XXgnL2wk+QPnLEGm7nuarL6MdIlmbjPItCSS0p1wakvqebwIFom6Mxy08
lTc9QXrDYKTOYa/kqr08JSnLGeFhMLXCqxg8pWR/Wft9ppwXNFH6kWZy+3q11r/U8/7vfQCL+wYp
LFvqWOE91/eQFq8w+AD0eDEnczIKbIfme5yuPLxs0+PrVEs4ZpnEiOPF1A7sSTX9jFaOZsn3LVkR
w9Rce8K07+pUnIJlBoR5fy9GornT3I01JlLYhlLacudCRYXSmk1/uoF/wnHdLW/bep13D5pLBY70
bqGBSbiow3NvntKU154jS0fmnET6eXlD8sz/kWFK1mohu/P9qfRxJwTumtUIYGAIVeG/CcOyH0S2
w0a6v0Yysi8AxT6ewL8WaDOStfcU2cNwg54UReWwDxB8vDnpsC7ZUW6BSC1Fdi8s8kacB0QRLRZZ
0u1dUPDfH4RvM9p8+9DuSAfJdtsjUwSr7+zIS925mab8c9VTJ1AQhkt5p0ti0uDZQfLiEyBmL88z
S9rSu5fQCMg161NoK0FNgZeBFRpLrjR7o3lZFs+V04yv8IanbJyDaZy/sJdpdpL1scXoCRAbUpv9
QqeIr7EFvLi2ooXLk1/NFJeNY6RbWOe4HhXEIByN4pM0dXZqwzFH+d5mEEZjEK1zGjsSRHDqWNy5
Ja22kaMlcB/nhp6CQIwpcpwrZeSAZY/VHnEFze3iGSXWtF6HjM+o/sIgyuCrKyqo7TnKXOC/7iJb
FUdOlbI9se8nRRe26nosJ5XjyYN2Negd1yuP1Fj2V8RvOo0Yt9O8ZFKI97vi+vhlKkV89yo9wipg
/NFY6cUrkFIH4TR1PVXYhxpjH57UNVJjAyvkxy3iDNv5/4yMwnuSomlMPt59PbOeIsecyeqV4D4F
QLapUMC0as+c/CTey7kNqcub0VVMHsHM90kG4F8HP1QC+/RLFn9qV0gfo+0Hu1LK2P4n2mk6FyUN
r7iBBJ1keL2wk5OX3ultQ3J22exdoaJ6Vo3Slisuqkk9Ncc/p2ocf8wUu9Bch3OirT/+YqxoPJiC
gnw7YTdh5sPrSQ+wRfKsW5nE6E9PlQFhkLAdzB0ZMMexGMu43G1twZ6iWA7DGd/t0cMpC/uL9p4n
KSCZTpstCD8x8/7y2Qqc2wy7pf824Uy9txWaZ+jisK4z/UuE1QBcqH61ZpSK0ECbw+j6uXimRNLl
d1hiCRlpo75Vu33/hPFyGQobG1BNGsNQfFeR8fRL0Ee+5j7t/CWXU1Advk08lSb2YVswvfiXUnWO
IVKIUrlHlgh/Wp2dyZLXSKhyDHNaQ4G0GybYlHJS0iw00SXRgPotyoi2OK5dPPPqOqWPFAOQM1rJ
DO+ZgUnEDBm0/86YkZ7V67QkeijssttJ1hgdDAvWNsGWOV1naBJL44hrUBODUUizcmnYctsgriQU
BoWDz60nUIQC6iVfsmzxF/Hr+3RM2axt3bK/lUkeUW3dut7qzq4izU0eqPv/ryQRWJekfafwhQVr
kW5bLvqVGHwyobzleF5JnbRRLG7zaT3TYzOGayt7h2knisG/QmS04QFWpNg9RwbBVyaKqanCeG8T
3TZzh9vw9GDtiSr5lm2intlg6veRgYw2EJvip2s/SJ0fa1MEhdkzsMGb3JjZNXoqWBsIKJszGTzT
VHoq8DIMCkFOcfMAM6vSJIVxTcNmKQJG75OATGFjRTrhU3JjeucgDcSgMwOvWpXmSXJRjqsMJVS9
7YOtcPJpEEWx3BHVtfqxWFUqWIvmoxsH7qAC5DahVbF3U5gjfddE91smQBD3hA2QgBK1WDEwlPow
Llse8napitfHq4U3X/gUQSOD+rvdUfc35dTW9kZgjdn26uoIMSKIarXiqaa2vzQ3cDZVKuR3EJww
Nx9gH42y+e+Cg8b6AALzJkpIuNZN5e/p6OwCwhwBeu1PygqmW65qLWBKOa17KYnBwmmKtsshvzwO
isxp+a8U7NA0ZFmNoI1nMmhlMNaNpJjDeKpGzLd8FHyAYApZEjsxWYuKejCTrH9B70pYtVPKkQEm
PMHJhA3Yw/mf507mgwLtnDrOa+KNn/vsxEjv1sj4rPUC+mIqFVW1sBA4JWVe6iSatx4zj+GYYWNx
TdMYQl1oj5dLmF4jL5BuRSgx6vsaBScueCyOwAXnN2DPCLxJWZfmvDZEOxZlYlw16ObSD2vmCusN
lugCH1iTzu7ByduLqcTdDCmpY28UMz5xoUvSzsxaoMSOGozVCUapRkPcEEMeiiI4LQkUuWpLCOuq
ZbaRQeoxRy9oJziq4R5TiCBOq7+SGJM4+yk4503jFtmWpgorSNPOz5fa9WtVAEfjwa2zjgsu9LkI
wBJpeZmsML0yr6MTfyrPFEXWK8BSVmWpmfPqruSkBA87HrCJ7x/J8KJI+0mjRSnh7UuH9LGKkp9w
JPGIhPCSS/a/+EBR9bN4FyuseFc2vhpmAz06YVOebb9byT6fwlYcugRjQkgQhfAOBEUOaW2StVBi
RXQhBwWaMbtOzcY2ja7R/9iwH1BFA2QU41IGrr9gK4jmWMqFENa8bjDo3dSX9QDHUp+l5yyqCqQM
6D/0x9Vdi6MM7nkFn6e5S7HMUd1PjlPfEq4qemzGHGMS3Jf3uszxgPwELCrwf35ku+eDP/PLgzIk
gLmwhDQK59bXvrodvIdwhTCBNoaKFOVXn3g1ctvqd5mbgbTxMkK72ywClVKuwlpmtfilVXUOX09k
dO3lU6FzbbhpDBcITKsp9JP66dDFQToxOAznjFdIXyafW/LhVT/j+iIQH41hUPRfOjffTuNv1D4+
uPFRjVNudClpMtYgR+6dzgIwylQM0cnl6V8/i1QmJ7nw3BoeTwdqXQqGBF+ss5w4MNIRV/k+OHR6
wR7m/9zl5mPu6+dpSOi8Sz1ZQodsfHSdZ5adtkKoPN1UAK+YJkENwrJ4et7lT03wSt9vygA/b9Tz
R7kqNwxF8EP3O5J6x5GvHCSlB2tzX00PiUT+r0Gkege1HfM3hEa8CtLlz7UITCxFrAJqpwR+Qtt3
BULIEO0f9FjjRZNriBLcu2qacOZwhCXOKYo2cVSX6XOuLgLBJYrx3w47zwSxOEkOBNcTqCnprUJk
A1/recBiH5sSqtbr1+Cw7PN4V4nFRv3PJ8iC8A/iX9P12YYulciuGQQeem4MWZfTilCgoKJ6TOiQ
rpA0A8yvQQsGPCjdT2EasN60HEYKwqaACSc52HHYljn6m2kf4R6ZlSOxn2UZB96CNiTV2x2MfSB4
hmXS9xCFEiAWVNEkxDDyekdHSKtVjcVjYODjM7MTYmYEWsYW1Jd/0Os6t/ga1N2VYHucahsX3OQ2
KuAMU0UkV5m0H62+js3JHKBYaOZ0HPy06Sc89YbTFjBR3nmj4BmJbN36USOj1k30xVorBw/olNmf
qIh0mZRSZeBaSR2jeqLxVVh6K2Btg/RccP3xjlb4Oac1zliwho6GFwTYW+4Ai/dGYtNryPuYtTvO
hVNoBdTaB/wKbk8migi+WiEp35T6wQhvN6o4foGhVLMj/mrg+JkOYWV9TErNZ6fzSnf1zq32xmzZ
9tPS/BtVTpCMtB4jYzqQl6AgDCcBPyEIFacrphdogEiXJX2lkkisIsoKsmB6WXzsre466WAxoay9
sXxH75sq++zHaTMprdB9tmOOBPFpA4/ealp04sflzMP6mn+UyR5gQrRXFwLZqN5PEC3kZNypSXJs
S/nw1zLXnmV87FKKxV9YUKqyn0MRmi0cOSJRXjDF24OoadAtVxTggm4gemVW4eAEvmfleA98QkX3
yr9lqfiftjxk6wc6UdQPP4NljXlMtcwBB57YgiIn6nidgS1mEELauQPO1gLETR9/Y4LYIkTlmdvO
PIqYGt2vXrcfqGdKOeyMVNrMoSNad0mo5G9uogd+gA+LmjNXbKZUjlqyPWkrKDZkggCeYrigETez
74SP/3+DXUGC5loLvzNqeXkPCE8bqZ476/n/kmGHRtkkqg2+VFxlDg1KRxDf7M2oyajcllqdskMX
BUdZj+RuFa+g/qG1a8Z3cZLoMRO3jwbqXLIh7jKtc/MlfqHOohwEp+nfRTAB2ArApqXvsDcAy6zM
UEUvn03LT5d6KMYzmeYl5y84oQPdYICRLO/OErHGVA9L6q8W1pYgG5ach9EGU+6XqfbdwIPwwR9U
ZRlBB7qKv314jQYuiIL9dh2jR/8AebvrGH7f7Z9rSeLkBpnKlh4RS/Eo/hJLL+UYHbPZoVGG12WJ
wLBqfV5n/Tb2StaFsHV13KVEE3flgTLEedM+e6wugvDUv5rirtcbLj8fNlcih7KmlgMBLTo6GA0T
Wydn26kkKj+ZBOjHpUd7KPc8jvloAniyPKE7fNLLnJSivkRFcAJLQn3IXMTKDdCQw3Lgk3N0X/sv
kZt8XgQiWx4I5GuQSTKDhu+tgDra7HZe1Rm3HpwAXULyQvltpnplo/iGhzgLZBDj7YTWamD2ZyA/
xwVIx6H/SHwL5A+/7csDOyFp+7p92LbZaaV223Vt8Px+kv1xDYwzI1S0xEeibtPp4w3quOM+ZoJ4
IbEDC2m0ZlGZ9cnsi68ayQBfAIVJ5+w1nu4J0huKbUEZIVwgvtSjkjtalu5Akzr8W009ZFEcjAjy
vJYOXJIrbyoQ04MXr/CplQUecpX8v5xRTsWfS+LWm2fi+KmfKsWCBCMiKFacq5lpXdLeTkGZyuHM
ME6C70IjXSJFUVG/K+060zwOHXw+eDeFtH9zwvLJZ2oA9hPxB0/gsUSkCKw8xR5QgEFaO/noE2IN
Ar+rgVyOoPPrc3VcCGerphqf80zUaAZL2XX/hCa1pJIZFKXYbk997VlAkWeSnvsXU766NdziTCGa
7gZIN+ZkGxLHEsW7vk52L5cn3mVnBiQCogswBq9Vos8+6omBA8I0dAwMn3x6kpFNNCP4S5uUO3DW
sH/64mCv5jTKhFdV8Ee0KDzTxLQezJZ6XF7eZ7O+LgczzFH7Nzoh6a5ggML/0mgA6UQPkQ3pw7zt
mhcPoX/+sVh7pOZ6rs+51RJHb6ULbSX5CJQ6beDupVsZAkOUG6wLsSj+ldK2lgj6MpWZg6OY+yqn
N0vxr/H/nGC/1dfpj2hIGP/A5WdtNNfHFyXlq2ChY0W0qmLbocdAg2f8MijwpzfwxePzIU99IUdM
DqTdn5nHL8lPaMpZF88ow3cgAjyGD6a5KLMrmyRXdW8tAwrN2J30lzY3wfafG1ajc258Tr6INLaR
C9fUJgsK0jMIU2rGNJD0pf2nNpCAupknbT1X6KdKwPk/I8UXEhxmMlO/bMoQ7ZadYFML0u8hQbpQ
9n6hrJT7pvcF6vpW2nEg4y2DVJnhDu/sOj5/+tSmhMjScLetSWNiykoEpR6HbGhcmkFH3GCA9yPq
jAWfk6a7bQALIIiEyVMEiAHBLdcLrijkaxpWuhHoALLjvpi+6tZu2rFHeCGR6whlppxCHs7AbpDQ
aIzNYWoRtffYePu2zYRoaodD6cA2gA0NPWg5OOo8dkvzzYZqWX/ePzK/j8pdufZsjggOF5cFcRzq
QFl0iH686hMbHakhBSHMijHwiKEYGYOpKCIkeEF7V9OaUQSVZCyZFIATWm23xBbq+WdRFLc/vsZ4
sjrzIE2tR+v0Sx5HV7Fv2678J+kqdrmaH2mZlXYHXgPs8TjSfWyoL95H3YmS60mEA7fc7eZUDVoE
Cve+gySEFoH4ZhCt8NiM7K5mdigOhPROkrqNDlUwzdrsqfhrfakCeJMvKJyLmYKpbGJg1HX/Ux4M
28u0Z7Hl6xO0/GWgcKxKCrqgGTqCn+5nAHJiCCH02DK2+6WdwpWgLG/SZw0S4zYPom1swOs6mOpb
FsVat9Z3SV4zSu3MMHvaWps1//85J1XZ83uyl6syEiA3KcFKO0Zr0sUl78A0E8v+DcwZQ40NKIyB
PEXWRDhwTbotoM0f28A3e7UVwhUf4tgzNejEsl15MNk2qJp49xd5Ges9YcHnu1a44ML6ISkzfzGO
dxdmenFA7MHSiFh6+UBUtYPOicisxxCSm9hDY+N9bsRy1PCXVaJgn4XMUWVRladxFTWx9UtZmhBX
i3DGN1w5aEOqrJV0idOChF1vd995Kj/vuQROjqMg2owmsy4vD1ZWpe2yMfLvJs2xR4bhcrBrUY79
KUtpUYaE16AhPNwAtcnNTJCFCiA0WH6ApOJ+I2DcemY6tpD0105H6c82WRodPij/9kLnQy/dodnt
T7ISEy6sImP/wVDPRdHWyhF2D0vIiZId5BY1HNgSzNTmXCFPsn763+tPKchhgeC7xS0IRLlpUPdp
IC3AhQRR7wJhuRnFBljNaRAytvgHqh/hMhUV10FvG6T2UfAZLoE0CLcDqgaY4Wfh+144oaSASQcF
dK90YUnf+3tKr4TBK+nvaaPOnZ80AmlfYsnakEinOawPTHLuljaKugdIdQlF7t74/G07Cufjnihg
xWRMZl14FzHc97livuA5tT5aGsBjBpsIemNBY/bAdz66wOzeoHfuHpW2rGNSMfZjv8HC3dykrvyf
mk7uaQwQf9FOFuqtptuaFQkAXsptxgz6PpiA+qLL5VSeIi6Gc90xjRgrhcDxoYx2gDuO+NEaDkLd
EsuDhyamqnMFCSB351xe2nvN4W5lB2o4/sbVtRVqLlVl+5v6hdA2H1zbwFxmiXo7or20GES2y5rV
1mDa6KIMNKxXz6+G32kjP0Ol6eYG/YDsqJx8Xgd1jmOsqSHBWRJel5ndKgDjjg11GyWkYuoFsG+L
6q792QSjQhP6Z+XXB+hkiJ/gexP5ZxM2L4x8y7fuXUL7eFrhYnbg0SzjuslwG3Ob7vwvQ4F6oBHw
7t0/rDS57fWjkrdYooT60Pl9AjV+/rkVJrSUmP5O39Ocs0HDDjd0P64zmLzT43b+HaKrY8IvyQIV
pbyxYjeXFvCgnltpKRJDmEJtAWtE+fo6bmM0LieGlekQC0N/GDXsW9//yyS1MfMaibd2QK0+Kpfh
oBd04OMJwNgd7T0zVrO3Q0jlOgZzcPkT1tUXyX0gxyTDttpZuCKIgucXzK/y6sxJBpSuwleVX8e9
Zpi1gVcHmEJhWvxKCfYgWjR0KqfHir73qjX26F/uyjhPie3CiBs1bmAP9XZ91tbuJjJzdlLCwWLe
1XseQf+Wel29qPqxle8LOVvUu5B+0QDNCoqKvkwPd/O6cxk08f6Jj/atdy5L16iwmVE6eImNqnlM
ueigcnYfXwT5PyN/oslPrLSPwNnxa6PUF8Z1oPgoQG0jJiCsQK8wz+UgUzO7sLtnKoZDLTrxAAuR
KwKbeEby4c98ck4L4AVGsPSTw7aglb4YSCplmk7Fi2KvoymbQULakHVF0+p02AD5XNPS+/REICeb
2TiSF+jQYpBFhMe9iSdThCu+n1nW3KWNp59MJa95EMOa05H5/hiJpxBRlY6vmjvxhKZzRRRRO+Z6
Qg/0GeRny0Dg9CP76o4EZe0XQq9vrbo+lQgEI0N9IYM1nW4fRKgxUK/h3AyAIYj94FfNvhFgwgsm
x0OcD9H+iZydV8cpSPFwa3ohLHe9Q/Kv27/vPewzCYYLQXIsoh6eKq4v+CwGLBYmO1Xfofdhwdel
sF82vnNsMTsz0hLNwBpRtsdLUNMzwVGJoazSEkZm3m/pSlF5k8EbX94bK6pO+wKSLR/FwvofS7i6
bf2chpKFbZx9MOUB6wxwSqM5luRYOfQVHIlYxrxKHxZMPU9uUZ42LqxRdKQNLkiNbLdGiHUqLiMv
/4MIl9FNKdMeQBEW4EgxVXCsfCowZs9CdmDO83v1uk/A8ALOeoVGpz8dW7wXAxpaUREjYygCeq71
aHHTSuJaFQ/DYa6n81OYm2QQ09MpxxrqLbYKrCdyhnG6bCnuBGDHEBd3GWUCOD7GvSlk71VWlGhW
8vr9TvarV2pjOjaT3MGedmW7d8y6DuAAFKFvTkk+F4ltVDlUPAE2xxO+weBTet0fwCkWHUWMQWsp
g1EFrjB+T45I6sMTgLhtckXuzGeAOEs8NOeF70qzFmhWuFeCjroxz1xztwVcNBErl9sFsOpSSRLE
h+22jzjCITcfPQy68B+BHl2oTngYBkrt/8KT3Kfmd8lNqaMlVozY6p2nmxYzCgCDdDPoOYfT1FN/
QQe0aVV28ri6NrqdZa0dSK1+Lc5AP/vaL+ouVWQZg54UWvQMrVrGX1y2VS71cvjPhJBydvsEglap
ozSYo9c2H463FOdcwYPiE7bzeODbsg7vJk7sn3eTja8U1XDNJge+jFe6P2RAX1AiV/xfbfaoxN97
gav/uOZ2mTXJViTKO/gBJtCz44qCNSt3uyabiokSWnDBoUIN9mzHc0cMAzTtiFXuzDyv0Z5afkyH
WmsiaVvBrNJ7fa/L8NuhfRg1mBFDqP/HsmNc3JLk0AvrxpvYndrTv01tyQXn2IrdXV3iqgAGOSVh
d109PJ9hH0Duxse+2OE9UN4ZIhlO3akbYYWWhof3da1NuP91BoTOnrrEnd2vsTMR6gaSgOF+HwzS
YoxzMVPcFDa/ecCA0DKT9sndcgBCJtCaWq+wQfNCICXTc+SoIvHvB8qrQfLKfg88FFq+bAVFK4gI
k92xHyGI0TKnPE/FHo/q+375myQffFxZeIOljWzD0SH5g5brwIrse2X9hxTIJKyGd22WqjZZhi61
a0P4GYflUDNdgihgWs7g2WrXt5fGSpRpWdd7+em0knUaojgEd5ykSH6jvpKxMVAmkGZ3ZBTGFaUz
10BQgQO9LB6MnVW/T/UGrYBcwymHHmV0pt/w4VAlB/NEuqzHs1ECn4FArDZhvQv7nwA0yg50yFyB
IPG5yQ/wlSSdV8Lw5+ZPihMzit7QHp6XGEhZFSpSPPgCgaxGpLXFG6oqmyk/3AkcFcv9uV0ldId9
cJ+jYqaCoU/ETvKCJQ4DlG/RHe4v9OIL8BmacEj9ABcBVPhudwKnryMXI5+usa6r1T6HPRjpydUO
Mm4iMU75sT2lm4XjyDMNqMJ+M/QJxpVidXJvBLD9/Z1JyeYUoUem8lJEp0HxKmmJFjdUVQraFvrP
3jt6ukltqHOjBZhK+NbZsrv7KlFFS6FuUCq6k9BnJ6hyRN1APp24jMHfM7evqicvc/5ouJ9RN5FZ
YR9UnZHjRXgjbhHqGFRjBsd5GiG9u8ycsWeaTEikw7MEbouBZ8Px5CSKu6Pv0b0nbY8REr4/DIlJ
mvqgPKPwzDy+5VDs2qg1n23mHL5WUDhrra9bli2KSBiR1g2NQ8tsM7hGpnP4ycOKjnd5o/3mm0J4
ANTQy8H94S2pKOMJEUMAdtr6OpjqXsJ9ryf3yBybKVF+yt51dtxZ/fjP4xXTtNalnmfQk76H66RL
RRT/WRiy3/9Q4hen7NlMF1uxg6d4LMS5/cHWlKEjtAJe735QBIDjD/y/UDnav4ozjnD87ZEdrZdo
97XTY45Ffs8lueA4kY+IAJj9n6pXrMikeM3BdVqMe9nmJaSSFzGFjlPN5SdaTEumh8NFldLyEhn8
wLHN9XSQ1aTaqX4Ta0JnZptcM5X2HwrCKs+yUDemxx84DvK8RQKAJcQCvtpRWrTAcAyvgiMO0xk0
uZpK9oK4QCVUKyNYTpF8ll6j4uuDxPxqbozTKkceA2gSojTGbmRLHpd7NbU149CrBUUfBAl4cv3e
uh65Qn2YEnnB4IlIc/wPwb/4MHFAglbkUbiTS4SjjW5jh8FU2HGYqVA2hSXC7zyvm0rnAxjCmJqb
P62Vun4vglG0T/3vQPDQ4C0ha9piofaAE6NTBVS2qX/hH2jVOWSnCJPspf7NpFWd2gBSYfGJHXOP
X8OlqAVy0C/qdByrwCHTPZQUQUBtUBO+h2A8zIZ8G0asxhOiBsWsyznd1d90nBsC/lum3mwWSbmk
0v1+4aFO6p+u9CVqD71MXOEKsOza6HYw7Vqxhwfw32Zw6y3KEZYIULWJn06asFq1bwmLzOjq2mzz
qoI+lsKeSb/X54E/xojGR05OR3z22WrqZ5SCRcCD2OqG+qUHf9oiL2WD/zBlNnrHoxRBPubQkqZM
HLCZX6+FEPp33XiBsddz4bTjdY7vvM0ds/G+/VPsDUmWU4KujrD0ohNzpdDKyCBlE32VPibk9R0K
yKg+4Bt1KYRUEvCBvqooa9ZDnOis+KGbiFvy12rI8en6LtJFyieh22UA456q9Cx36DUGrDcKC2BU
4hsTZZr9F/2O2hAqQFmDvtLeP6+rt2tNXXWJJ6IR6St9zDRBl9zpk4AH0WonGNp5JjXApFANVkzZ
kVp5XKtJnVBrW/aM0b9tspzutJzwVVVs4PZJUBIoHO2S5Vw6ZompRv5PLb65wz1ZsywNr/dObk/+
UTMGqK952vgUMoGBltroGzFRrJOxiSDz+IWdXphDnWEvsk3+9HAddOXKwmx9VlztDExjYo7S/pPu
Hf47XNIE+WZ7NRr/5o6AlwSWsAtiLyO7fX+2VzeO6xuHBxwIiNwk3NnIxdCtRBij12S5ddj8yghF
ZBGTSM0N4pJJxSlBvQLnneZSKF66Jc/zq77kFS335CMktHG1+NhVjPncdrSgsFe4qzQriNf5O4KK
uayBC0gBPlQHpB5tBdsv8LDseBwQ4Qrt3U/tP84XvMwJO4imjvlCvcnqGPIQudGK06gVAy912/WP
EY6mI28mYPe42+Rrq78rBFhCmC/v4zVF8EKudNz4x1YTwSho+MTmyjB68dhzkBwSXMQ5eFzlZXmu
BDj+ug0G/4fwdLeiML/N/xe7aU06/xR6P7UL/DB8byDkjiPRqaX8inAvYhsWjGmqhX0qdtj9ZwTt
KiS3l8hRCja/JwGDtP1rz9nU453Flztbovq0+NGyhbD5os1PiCBiqws9a+sOhEHsX5X335TIyJIu
Y46/T0qSKfkc9BcWGFQUU38fVBaIaiG/C9Ugye8IdIjSOJEfWapGCD0Uu+5wmD28tLmOv6v7+3Zf
mRvNAmFhGMaw7ePq85aY7N0LY05e258Z4HVV3WU1EqXkhvNEQ2p8sEofyb+EhA3x1K7LTBLgcDKm
Whrb1qUVz0kNivWfj1VGQ97BkPw+fkfBYzpQE0DLo1c1l2IBDMXTPlnVXPiywd1z1Upw1A5SdUh/
aWc6dxYxs3UEnMHsBBkN5v8IVUO1js2CZWY5NjEktdIUUwF5dxAOugBuf9fz4ad4lH6ltqY+Tcjy
g36ukjxZZvpT5oH5oB4c0WXZVtpd4jQu2OUCTM9j4cFj4w6nbC0TCQvMpJbNGzk+9SwSmMRnYORO
dEaZa5f7w4IWUy78Q2OtYyEDRcxkZzq3hpzagtYShteDKUjjJ6bBiGCzGZbJ9feNi7M0f3f2COZD
mKcwseZSF6AP2/X8AsddykE1qL1uBFOdcNIo2bH95gKNLZcKDQ5gFHRq27KOJVaHoJsr9fV+ATNQ
870WAmnq4KemVLlLLR+a8iQEPl/khDfMyxB1+xqoZ9PkPZrCFy2BlQfxOjecM7ff29sQ/PQoC9K0
OYGb+fXJtt74Vn+ds9XcWr3bD0W5/s+7Kw1Cm93kHrKtkt4OqIbLwHqvpcpBR07RMnWcX4FRbU1t
OWmlqUwBJAOo64b6eQIdNiEzzLTcbNUNZiVndhEKUhqGk99oOHKzNKYY0IgzVRwkp6aHj/C/Xgtw
ZiyUG3bqhYDXXtVdi7bsd75joxKjQ7WQ934XPpHm4bVAE05K+8LdUzpOOMsywnY6XeZbL6S0cvUg
kdqd/9FK3IIvaAqN9N8JUrRfr43Au5yxUrenoAzA5XFJBoEkAWmd9Ke5kXVvkZP/7tbLBRfEf438
9ALaeVeSRIl9NutJVCSBNEyDm5VqCEQfEmszA6u9rZdnoC8sFjzaSn+HJSTKdMibtzsuSSGd3L0U
LHBWfI/Sj6ivJVsgNMPZwP9gavLtOCQyFOvLtfaAc2Nf+HikDUcI1BBXPAvqsk1WXpwgGT+elegG
HzVAq9g8Sqkrtd+fSssq7xhClwlzgQYRj+C1AIYT0nXRyXM7Sp5lRfUZApjWYikLcU0clwfd3PYo
H7SKSYrxzLR1E8SGdKSFgBkDHuPq9cjy/4bWrk+wC+dj8DTMaEHvbQBpg/NPMobnn+8cgwFeb7zt
zSzGQBKs8fdS9Wlf5FOVS0g73dnzyyGj71Ke8uRaBwwnNST/lB+T5yif6P3M4M8JOUa7q0NESW+B
k8pWgbTRkBJhSfdXC05akciEUKoqFg2gaVwQDjhYAzwxLbVOLhC7tooXCyT3C5d43zzVt94YeB8X
yrUeS8aDVMDtEDScLOjXTU/9+erD25g04EDf53pj9Mg2c9EBi5NDjLKbHHPb0X1ZOzCkpjQz64eE
uGK6Y5WXGVfLB07MOpLVCikDO9VmK+pmNUy6rC5zd5sjF8zQnsKq8xW7GsP53wLD5HlxRfkmNC2T
ZB6+RBqT4VXFAj6Kd5nIlmy3+Iq6eU11XTbyhrmiElbWtuEnrXxDhlNCXKlFxL8wN01jluAo6421
qlcUuaGJB33+DdbhILO1diJ3vqSgV0iqp1tpQtEy8Jzs6TdC+yVNR77/epNE1/E3WRJ/n4HM5VgX
kYPDQtdSJCRI9Wmuw+VewLDQPzlcq9wl7gGHXFH1NJLcb+5jszU505hGANHbXRGHUfIRRQNRuwm0
BFpUU5yTJdJRPf/ORw/YPhtWkdnn4Nyz0M1Q2sRQQrn9dIYPSR1lVprFdU7vzroF0OqYNg4dhLxn
30EBjsDoFmK9lIyvnRwnB2bnC5NbqOY7KyvUygmpo3jx5gy18JF8hscXoQ4gOIWa8sT23b6i0WyN
EZh7wB9/vh0cjFCSiN8QEyONmXHztqU/nimqBVhLQ7CBFPH4COroOjP4md8IRJsZkJgly5jVs73Y
/3jtFnrFyYS7diF8/x1gn8vT+mbRbezVxTJaOK0SnnPiOuxszGsK2vyPl33AogwBKmDVurnvt4XN
OUWOYIvn+D5GOmd/vJtoEEvgKMb54GYa8g+EPAwU0zttZdoSir6KAc+9WEBF2QUIu24EW56Rc1ZM
zn5ZCdKAEXQE8tRkJk9O0CYIAw27g1OW3uH2Se2/ZEyhlwBLMha45dexKDp+MDxWV/+u2UczExMw
HJR+N8a8MAhGKEq8xciY3/z9apvdvDRc7R5YJupD1f58SsEfMu3vOjygC5tTmSTIRkYSlI9yftOX
TlUgtoP2YxVK6Qq7orETvF8c7/vnAKlc+xg+dKF+pcwiyKYE3baXRBVk/PdMCHgoF2Qh1RXvvIJs
IP3hzPehP4Aiatfd7kFKrcRHqJZi21T3JPBXZWCqVu9YzkO1Mq7DwXaFtplBbS7LkxF1vMV0OBlG
4Wee91XPPbOTlWmQ3aOKVQnACCRd/qa8LdnfivwlF3yunmwfE1qXr1tA7Siq/gKv22hADIV5Lie7
rTp7EQ2wTpdTnhrkhE2UIxKhBF/dZj25jkoHsr/Q/ta3kC68DI8MBK/CwxctDueWh8kPkgOz8XuS
J10tKTZNcVJJ8isPQL0AXTG0+J44FrOSJ+djzrpPuevB7eChf5zCT2s0bWSMPATR7q1AcBqYdLBD
FSzL9kyXx0qCqq2Jg1drt9bfr6OEXGZAFELMr/qcieeNg1QzsP5uTGmVRsvdrhgGkODEWfbxlxcS
r+j9Zoh4xnsJk4K2S/v+TkkF5NvI5ubWwTx5ssh9HepACwatFLDJsIHpCMd2OcLekgKYwd1Td9bu
rjyfbs8k5D5UIAEpeel6gENFK+DlGRevThKHRpl8pkIaFYlp0wDox7wJo+rxiUNZ7yLjgnPVIPf+
y1Nn31q0as99mTxK5pdc6pUgEDLkNyrIAVAh/H/aW0+FXUDhos2q2NdD9I5TwpeE72f7cejxN/wo
ggGQ71y14K4vvwITrT5bRCZR11KAYAI/dse9XdTt5ueSm2gbbCM8fPmp+xL7DkcxeEwgq4Q+3XCj
TBK9V6t5FPsAl9Au+Jwu7VcPry5Y8X+KIHBevqCGHuZhzV8qOosCcvJsClepxfnN0P20zRrhxLFA
m6h/HnMz1eZGdE/mPAY8sbF8GS3d5cjZ9gnqvC8KLavnibxTYw7vS6Gl3jpnoLbO70MVIiVIk2JZ
eLYHATKqUGMEalWBrXxXbuzqfMbVijKGI4pAXzDaPqbEe7ijA1l8WBvqfzqe/jmCpJyBVEMNUQ4b
gqPXplTTv1CDi/JwkoXzks3oj+/Hx9KuTlBHXiA/YHPnpY3r4/yyoyTNkQwkcrXcoLbFWgYHlce3
OMO7tbdRCnoH+61ra/61+wBJ7Vrqw7IpCuaf5n1sDAP5m5TZ7HKkdDdgieIThY+fnX7/kyL4pQ1Y
5w5dztcO0Y+iWsF95rNoum/2bgojF9mTuD4iM46iXwPD3nYjrrEaT/4+kayHouqqPG09tHM8AuyN
bLZ4+Q29JWaArj3Q+N5fUb9L4SKlVZDB7H3z84sn7JTWKniMw8yiaBh/u5bvqczin+KiWCrIoVJP
3KS2XxPy2qmBXqNQTSv8SZn7YLHEGAz99bnHAtD/u0CWnIBP1nPKPB9hRr4B2fEecOXoF/YnJsx7
DxsCmSYjk6kkUUoh53b3/6eZEMiWaoWHzHtXCOEZUILNt1cF2Cj4da1vvk1N4MazlYCB4n2njDGE
VsElSy8/N7CfLgWyTD+y9qcpH5+5xoO5D1GaIspFiWb6jn/54DK9D4RON6WyHznJZda1zWF/dAiw
oEdcTALCZmWZS69uoA/9ri1cvQwNXB9KRKSSbJeoXulSMKsvUEkKhx0WoD+QsKe1XluM/8Kax3GP
luDLGXlj8/98FgXbhSt1w28PZm25K8UV6sO9nSTfuM9fAzjusKIa3hbfwOa8i+gRQkhy0pbCDLlB
E3N/h+gdBVvOLrJhttI3Zma/pb80J4Ue9wuLQS30z5t6vtK3/UeM1cWazzJj7A+iKwBNrQZ3XkcE
ugDh05zQ0WIEeV4BKOLfdh/B1gh3CEA20XHPGQTk5XGkDUgQPTq/QJxtc4eG/7tMh8Z34D4+swnV
+gDITtjrb799IGC1CPZ9TddvZTvE2GQhv1Bz4TnBT73IxgE2hqQWvnT+ZfEt1EV2qEUTW13HMQ7s
chG/5rUhOJrYd8hV6gwJR68u806SoZ2yqZK8PY+7SKdJTimyybkitjM3Yty2hV3Pkl3aeypsW+e9
LaXfBmsczvPJJXrSOngDwbfQ6PiNb+4uVlIJ4aBnelobWJRJQC/ZPQy9ydzrEqUnIs7tlpwcWB5h
riMeIJo8G4mad592ZIe9Xv/dD4xHSRIjKoxLeS1KuPTyUghLx67+ZwGxohjuo9ySRaSBV/NoqYRO
6wMUd+O4V8tO64/iiwIvCjym6AdXWPJn54IuUlITjU1C59m5NlPiv9G1fwEEtftR75T4iNVWG2TN
gYAqMpYgB1WafhU2LojTxPa3NpQg4R8xxGSnXSXdgqKxa4DurRqUvQuUh2mzw/cOmLdJX51Ju16x
mnEOWN9SiCrWqpUmwJwcv2Ld/SBOTSOMbl4A/iFkYg70qMF6grDf3G0bxN8JpNlAk2Ckat6fZ85J
vBae77yuJZ05disr3gY3hiAdverz/5/tYcbVhhNjrWTtnRY3rbaMmXz6KM1oLLuLO6jZw1l8d08w
qa2386HaDC0AyLO4LP433REnlmlAGToIwOxbZM4NhT4GEbV8YgEODnmoMd0uDbQ2CKcz+9jRaLDn
EYcOtSg1biq3N5JtTXAG3OXjN+JK1JUr2mnEhJjBHztpPp6j5PvUaA6j91n8mUypDtwAAus4Uz06
5YgLFUjryvteaHfFBFGT0yrWs9YQOYC1xD9THciNjY1zRQkoZtt8LLvBXskCL70EQTZK7J1QDXjd
YFWfSxvvwLD05I/l1JrJN2vue4WKweganAlUNnug9poLiDtojT/JZAnvoiqLPaNMAf7ewlh3Lff0
O30oSzpQxEuj9UIT85SiUxenrfgMcv5xxPVyPLVwyRsjiMrzNRE/dAyu05vboKlwEZtgXVeaYbRp
3OzqAp1fmSj7dxkz74dNWBRTxC1SqKihF/7dFDj0+veWYhNZAIKLGwwfST+SojPDgYlTqZHiHhjR
GV7JsBY6DiWkRHo+BDyjd2344sVJ60fqIBfPkhbXOerFuOZRqBdhb8KKILYOJoa81NroIG3uwEg+
ueetcbpisbBxtZe9XmMWONaGuO7X3CkEMq8nNqf0qIsf8Vy6PmDET9xw33R8Qom1WHRxy4tbsCj+
5tuVlmFf5fzZ8cb+KA/tBooz/lRr+KRa9CdCQARCtAZZW4n3/MEimmLg/+djaJ44PvtM0Zfo95rP
H7EN8eDRawlqguyt2ApsV4Zf9r50fde/UMQkPKD4+zMKPQ4jCGapkq0Rj0qxrq0GsRHa0xV7pBqo
1Ijhnaj6/jYvnqVRKSxliAhxd7Ar+QKQGV2E0e/wQMnpKVHnsVqwZo9xOid4t50C+p0bQM/Re4a9
VsCjg12+yVYJC/hjZLzbBD7C7dmYhQ4ULA1R6SKl6x2+vUUhiME1s4SSS1P/xqk5bRxjGrMjEfaJ
CbuowsdfFi7KQv7z+wZ0ny5Lud4Z/bNOefb6Udlw9AqkDrwrTOVI4yBVAU52XX+ciXcWnJS9/Ue8
Dtc1wpKq7Ehi6W1L30q/5ATG0RTroKu2GnuAHpBrcd3f1ckUxWeC+iCeDUfr+7sFaec5//TayNuk
wrKtqju2EXYiraCrliuNOPHFDGqfhg6sJsR0TGTaQwszFjBA1weFa1zLURu2sr3hlD+YntHs32SE
iUnsSW4V003DmqjoTHzhaXij5dFr8jDsBjsp8FOZlIMAZrZbuutRLqqcipkQHIeeXSQvdp2NPmqJ
pnVFQLF+rFXHz5Jt8CsTDk1l4vGBJslTTA9eCDay/veAKn4ArKo5oobPNdrhFjV9JQ5oI3jbdmxS
SlzeEcMqxA/PEvtd+WRqtMLBu78dGjIXLe0odG/IgBICDKpDQUvR5Pg2/OxazsznEpTDI6Zu4uqR
5C0XLU35WQjBm6+U6ifiU5ui6CX8gTa+8ngGPtoPcF3Nb+Lljda9UWxrsUlY+U9AhfAeqe2sFscs
5E/Lbz2mc4az7RCsc05dDhaLvk3tImofZdgTrMADxulQyBERjBrtbWW81+pmOnUMHW/78/z9/rYr
3b1wuIe2SmSuvQJUcEkm5DFk59tEVoO2s8egFmRRHMaXXCIwFqoLsIZKGsdRHfWHhOwJDEUloyzk
HohSagjhYrDRlycYTQTPsWO6hS4hujhALwx3rKur8hGqMKO5qd2iOd0gB/br6cSRxnzsbzWcFzkC
B6NjX4M+XSOdnclYYWjNzCdMq+XhltUbgbORGCMEJqvY012VUczzI1UySCIft8zPBcxIJKXagIIj
ccbWDVq1cD3qUT15VsjSSDmFOsTLL1lOSV5hrgTY7vLG+bkUa3n3sIF/Grxe3Ws/CXJQMDwNyLfJ
vqsxMGkhaGXFSLUJXWc+XdCwQT6nhmM6gc+vo6wwwyLqo2HMl/KFGnKkyG3uGnEU9ntLbLmEezzN
atUnF5mTEVwm7gXbsU8yPLBPb2sGO50jdaQzDJUTWeqimUa7QRJEvkZvQQQC9jJLGH4uiCnTwzFg
XcLMoJ2CkO3dsyC1X/3BoI63QRwxOaIamo2IZdnPnX0BW5KYVi7Hucrl+q+jCnHSefdA3aGdEI/A
EEQVmqJU5BVj9+jJC5fiy1ndI3WIWbKIZn1f5rRFnBdWl4YjyeFULmHx+yB7i7kf8x0A7PZ7treh
vJO/lJGPPxg8RqBM4zV7uOlTuZ9Y/pMp5kuj+ANN+EUaqh7QVJXzYsJek+2W724JfiTfxaSMwCYm
8FdIktUT0tZlQ8LmPxBF9ErQ+mQGllj7CZUB24PwnpAhF5OUeKCnV9CF0rCDMECE5jEGCXj11d9d
1CKswIEH8h2mg13SIJs0EL5u+3o8iadxu79IMxEhBSqsV6WKPHZUfBAcN6MjfQnamMZ34W4rCS3t
BDiNtEQ/DCRWplykTeGb4vJQ9JVNad5w9X6olPuK3tAv0hebZVOMD3ZtxS4qQLXebecFUKt7pU0N
C4+1UnjAMcUJYnwU7Z3ovpHxks5OcmzRtmbbyCK4K8keURoC9v/8f1Jc9LNRwIJmlFs7ldt0tWbw
yYMMouZdrfYCRDmPxCT96q/ezcKZfdVnYqC23FBBerrfPYSD3ETMqkJCv2RliXnCR/4X6dT7Vaxz
D+xj57F3k+Oabc+33KYOsFT4ZkCjRJuTs/jrEumzGXOL2LI4ykqCscViqqjv//DnR/6QrQEJjUBg
+lluijwNgFXzwnH4SZKZoUcNrymRVpm+D8SFFBRbaTJgb4nBPEj70hFV3u7gayYw7AzGNYSWEf8A
qlo52h9qcxTW797L1ERM4M4VKodeVcvvnC6OaBG1xy0ifeq8BmQ5+lVChwmsdQilu917Ap2EulO1
7I0yppXdZ9dj6T9KhyBEtqcEAVWDd4dSy+NGCiFTMQT30DzAcrsELy5ARs37+4m5DFTBWWjeGJO7
i/XRHyALnDyxAKOyrNoLBUCjnYajmMvQTbUH4IG0XG7J6hyVI7MQbjxzkzIhYdkR+8zB0Bnph4JW
Ta7hSaCvSrJuMJEvYh0FdrrqdTY4P6EEp4orHaqqj/2aoxdKjFQvk430b+3m778O/Hn5ETEunmZA
TZ8z4lkMwy0PN//CG6BBCMZKp00F3OPN1fpHWqv6pZ2m3B58D6RsZebLOKOqyrAMcH0MwMmfopvv
bv3CvLxuWdb4BlQdJa6aSE3wnMOb/ZgkIm+mZ5CSuJUw/ltJH7ScM+VRIITRIv+8NkfT3tEIvWK5
OkIkj+wuPWgv3iKmwy8+MbpGJ7JtwyHxpcObe50sBg58KgQSdpXvWoX0/WGhrJ7sLnlNNK9w74U1
aVGYhzIoSmQKb+8KklYAyKM++2w/f1B95eS3/QQ7gJnGqx/+O9cIKWA9tfRw5j2MgFI84pGPMnJK
3DJk6q1VV0R+9gRni+kZKc7iN13FmEoH+Lg7JWDmNXbKeTf0R2Yv5pgWephehV5UKVeFzPcq/CJZ
auTRSefcrNAH1a8hKz3G0eLy5DzELJDrl1LaRxQAr2GqIHTuRWPFic38KB4qUJgGegzVugfwEMyE
j4Syy9ajd7DD5j3v2yDYvy7pibIBZDwRY4tNk30Nzz9KbxJxF0n3CVDfh5xxpnRfeUYeVmnOiO/t
TOMIsPilCbBqar3HzLOwI0rc7fonWOIwiX7adCnP9w3NwegO0rd+W0zumBmBTRdf1YDZaLI+moho
8dPClJULsMvLG3nAEgApm3JKx/UUsiHdcNb8NnCd6CMxE4/YqoNi9NV7KWTvd+4fOvjUrGPDKU+V
hesCyhfHa6Ke/JDSenPyF9Tn3E+q2QXrjYtVnkedOveJL+iZ6dvyjFj/zsaLgNUzqdkljoO0UkpX
Vz6IiXqfh1nL6Dz2e4r7XOgVZ19QKxRwVs9QQ4/g+6FCQoIuSc32Gu2Ud81YckI9/A970AJ4jGec
0enYqtXVCQTX6TP1Ds6t8VlHtz7HjYxF5u7QgjZV0MvVOS3jMKUAtiMFkmpN8Ei8dzyjDYlGL2ut
3OW3BHideGIYVFFHAp0tzEqIlAsr+9UAVjVx0Cx4i+lKAJ3L/fd9CLMUE+J7xlzrmYZUP/3zvbO+
HRqa2vueF/mDKShYH54Z5f/jUSZZjGv00+2tOJAcIRrs71D9fUJ9HeHsgddWibZJH3dXBqr1PWoM
9oC41IGBNPiAvWXvbLDCsk/X/bZfS3ZQrM1ftWZGDSw1O+oqvt4fXsIaI71sm0OS1MfPS4Nvmxzy
PufrfFvRd2ry9jmUV2+AvGxgXw6fVYi/i+jh9S6J72MB0pk//6BL2aKSc2SLf0vcWjokM1SJJKUj
TQkkLEIcIAzOPe4ix3dFCAeQl+Aq8ijK73FZjRJZLR2tEsGNyYXKUL13H3V6xa3YFw7s2J1sBJNt
odu4K6uZlTgHwnDO2zWdByQ4sPRB7MtFTkzGep/GRcGjAEJFUZC4YruK6HgxHiiMmlYZkB5SQZWL
m+RQ9CPunHLlqQtc60smtfUmy5OLHwzM17dGv+bHEDIM/jzL85eLz4NmlUwCkXqKugp+7qFN3STX
wimmQCDUMsiYBhlLegJvjHR7reE3NY5kLIi7R9pKTV8tRiBSsn5A2Y6c1KbDxbi/ZtNlXpYjhFW1
e620jXKw7PPVYUgI99PzDUXYopORnw1XcHohyuYUTQMfFP3AjkjBoHi/vwDcRCZoOXZOUgse9/Yk
p/1MtZ9prvCxrDgnomC37u2gkTTL9Lg0GLvCbViQtDBLQqpWBTIfg/I8Y4ZzD8X7pWK8L3FXhCFB
fs/H/8QtO0c6omGgECEh0N5pj3+kEwxDNRCq1jN03/axJo3CIZ2xpx9abUIjKfoiJvHeZBLV8jcz
pFSkmBKmgsnT2JUyW23oKf4yj8LMM2pSKQyT9xl2WZmgJXNu3lY4Glfo7pdJ8/ZB9i6z1kdLpLA2
0VTLksUl7rL8GAJTT9yKgW+HWlDQz8n2Zzw9h5/j0j3smPcStj/oZPYudfLM9RRfeHgAgWVPDvba
6aUlr+1kWXvmR8EocbdLVeiog3RLwFiOVx3D2JKhHoVmKQySQzndulJCfIo5Orr/5u6KLJo+UEyW
iHYWd30SvSS71z+PyAf+WvqlCcpnsZ0fsE/VzKWvm/eYaNC9BzMEu2FHbhyNdRQ94XUiGyRCx4Lq
1L72quNEfK00gt6/I8vcGE1YutLIHam32yYuLL8yReYy8RgLmI5M2qaObakd1zuviU6R67VUpq22
b32kBEXXKiWx4aJyi6mvH9D7FiPHZZaRF3SeeDzAPKipEX9raSq/YWp5vldSFyGiG3EA7urzB40h
3IOz3Zgf3EOyOGJGAAKQVNiwB2HLC0T/KaWRCsZabJEU7EqFWsghuVCj/1p5ADHIGcqWgeTUswpz
S5PaUEhD1b08P7HB7d/QtLsfDDnzrNgp+JWaG9MFW/Z8O5CuF/mJeudxin2hlPCURmNWHWd5Fe1o
P3SQw57F7GTgxiKaFsaoJiISGLJ/9jOkOcMqns18E0Gzmk1lKXVYgPm7ORZHI9rC3564/zvRyrkF
2sEfqN9ci6hXyVZTsHjn3WkdhkZ8m+j+nBVi1uuIXo+787U1VgsY3breal3LDe5v0uc6Y0rNNgt5
E1B1Mj8N2i3b4cNnhfKX3EIsYmhpsLAyCfAdSfOSXVT+gFp4M+xxCXvFdzF6DLEvDYPjL5vxqLaU
lfPAvBeHOlSstCr5bM/bhRCm56ZMy86v8E+VYYAeamoZ3lxUk/pjbzqZv7m0x3qWYxvzACgqtLNB
jQLKLg69efyWDHxEoCW2t61HxWVMGgyr391aotH6BglceC+X70iJ+QeH9rYHuQHUTaCld11k5CvU
/47ljcK+CR/ZSV4tuWolk1jGy5JGyxh6/8hpJPwveRoe9/A26qP8e4v+ADue7zNcCwObgwVYZlqG
6CYhqgslMkuqdpl7pF4nmlJ+OK8o0wmJ6B3mR2pznPwZCgWKaHsRP2ZJD6LCJdjDF39heaXnU/2j
C/Ouzqh19M+FqyY13PG8WCXssMI7/LnCQc3xs6HkHXFMWuIkYOeAStq78UfG89IGlto4u+QyK7U3
0IEovEJfsxMaJg+17N1NJ3f+v5ws0+kb0Awrr4W6xkKsBHvjHNanbpV1vy170uUHI7nZOskMD8R+
nQ9CFU1NK2GVM/PovOJJ+ZqFOM5UBNxGV3JXycAspdIRA6WKyAi0CfDU5/WsxGyXWMYWfiusPSUG
XX37DccOlbkQOuLRX9tiugN2UXN7KLWk2JX5wHL9+YvXKMWV7FchQH71nbkiylyaSJcBfyKC2ras
EfHq+GkP4w6CEELfmcRN5/RMFM9zFwNrssm8xBBQnMk7NFraluTHXmZmIVROkG3v5OMXQxix8QJ5
aMlk490Euzl0Y9ImNlgWe2XbGmICbumFmdmcXdGWE5VWgm8+r81MblChnm3BohtQok4aR1zgyK9b
Uvowt4TpL/JQBXpT1vKpACfkJ3nFawTg52ttV6GZQbWdmxY3ffLbr8oR72E8qeYutTeNMjNcvbCz
WKidZAQ/d8RHKDE61pU/yBXEpn9xJooDNszxRJEZfidh4SPv7uGfzsDmZED/4Iyf4EQjTiZOxKSU
YmimRxmvc/Vb+7c4PZeogUMgCAHJuxF/N4GrZalD+kvLKQOLQNLDVpCSkDG36N4ZsPwvJ7qUPCdA
3WomMY5L7xHq81b6mB5mifn9Dqu2I0zfPhWRubLIcr3UK/2PM83ciHw/E+FaMsOlv8hjoAbJLewq
ntQkuhJCP+h/a1G18nS1Lh9MW6euK90iltvzqkH1l30kq3WEDsiVZHDGpG9Hrl9IzZb9WjRxX5dY
re2uQBnboZfJEYW6dPXnQI6eWAuz7tFjmEziclZZmTlJckKE3uB1cQlM/z43XcjQy+DfiLkxHFaB
u/DpwWmFB7/lecet0TG9j5Dl+kIzn9TnWkKm2ALFpxZQjiz9qavzRHZSHupu1sOs4JwbxkZrwOgC
n8rCscrI/TBQS4jW15blpLJVsork+omB/ai9drz1VlkeNcaZdEmo21AsU9EhlPAQThfHslagz6WQ
oK3QlUj60AEGkxyRifBd1g4nYNcN2qBx87/EbAG51vGUER65IJo2eQfFsvpis4fQ3pdi0s5q+83r
h5CCw9W1lbkLt2XzAd45i5oThwB4zHYwxnf2pfm4PY4fHF/16RBwuTWHuYF+4fKpgvcWZ+ZJejae
JSCVbJWPs4zDbQWCy9GpwJTvAETFxMv4D7bj0lEV0u2zMwKlo3ewM9ho8pOe4x9vlQsbpNut62Kh
7WIZo/9sorgHsBBQIxCHk86WXeE0kRahd/IpP5TUQI383KsBJgy+tOSLSIyxyHEon6AiuxbPdShJ
udzAAxiCaaj+vn/jZUuZTokpJAQGbFKpJTZubDeKN66MkEIsZVoNEgAU2tNykWRvUwkQe7C8baMn
LNacqqZscwjkDQY1hxqotbOnioN4SfF/Wrjsmb+7GvuakFVSBjewhjYnBq5LbRA6tdVd3j2zIcsA
XqZPmIu6MmLNhTr5pO8UpynkC1Xfdn+iRry6J7nvZBbBSK3de4HPirBPaBsjKycOMzIjF2UPhOxU
s2zyjm8jENvxRWIPdcy2+/bqM5eV3lDk9nPxJjfMenctyttQAXAYTUAG22xPSTLdauNjE5GufyhM
THV138rpwnJibQaaWL7nqv6B9tJVQVYSmk3jmb2WUdTFWcm/WKeva1eIup3CHJvH/QueT/4HcJjQ
i+6e1MR0db6pEUSRPriWYW7VNLx1N6MgbhnnFbfI8UZlMJtV+2RMV3rmiYFmuKKKxEF7R3itpSoN
lBDUKaFlbT/8u2DvQ9s1TSxUhs4U+EMqYLexvB73J/jHJVT2Lx9p51pgxSloNgbUTeQvLTFs1+Mo
tgUtQWnbin0TLe97jPx30uKVSkpAw/+Yi5iV6VcDZZmHTcXtz47aRgMZVAhqZdv/BHQqD49qnBUW
/C2+e959yebsc+W3UseIPgHO9YR7DHYfEDR4Mvh/DDdtFsocPUvlrtJU2EskzBPFfWZ/pEddOVDH
bQ0Kv3CVvOaNXw2ZO/4c6EUJfvKrVUqxEJ37EBBBIbVlTKmYJTJeiTdS6YebFd/fqp7an9a2R6/o
NVmfxyiSIlsTs/sNr99ZNRD5OIK9RH7LvPl2Tk41cqgZnpJmT2Nqj0Q6eoFLvCipzbxC1FuQ0gt+
t1a7Xdi9C8915xCxs3uo9JxfQQeJ9EeI0/wHQw0kbupLMg1j1fG8Vrc8zjdWpBSLUUUmZzqtfVH2
Oc1UOWRNJbwQ547s7VSLmIDVBkw95nXryo5HSSVeNBwhdWPPCAr7OHnSFwgKncC39FKjpssNwFox
IdP9vVFB6A8uaX5SPPq0prMnlEmjWcwxUU3J0yDoWOZEbzS/nbvNiJuBwFkvcgv5cpDATq7QZW3S
wzLyNPaj9nnB9qPfJYJQuDOLhG4m5a4RDt6qchGjmJ1W4n1iVKSWWv+aXWnN18pov1J8suLo6PqS
o8a/Pys0sfeDiFIicCXlVi/v8RvazO7W21gL3xerSjGX+xq6FzdZAUSoetEbLiSca6UfYAsuRr69
EECSXjjq3MzSObFxJsnTgIg3marzO6H6N0xu8AS4miO8B6B66XYIwrmUG5JDUVTzwa360skHftoq
4ux05FCX8g0enNP0iIzEYLK/nndDiat97q5O+2SqPcRItsGGrbgbfxbzELIpOx55tR0pSAH9p8i4
wY/WdchzkbWO+/vAYtr7tGROe+w45RmnlS4U/EE2l/yXHzG5P3BIiQYNvizp+lQbwZLrX6iU3XJN
Tb4RwKWtjuImJ2zQIFYPzUbgyAHyfTMIZQRAFh3XYRWa6cuAHVk5iGuJtRA/aPLy+bmCM7Uu6VGI
1VXs+IusxRYmc6o+PXIdsF09Wr8hR2Kn77nK8pN7H2LqTnTuLj9nU/jMLOR33GgL7TqDn8LzW6Ga
fU6PLKY0DkzPuvohYu0oWCMyHni1Poh7kLZk7n2bX8Jsq3Jc2UwduJHIv4CbtQnT9T1nnwidl93X
nSumfbYcwEj/5PsY5BTniepT4HqaDzq/cinXkaTAWyDZO51sCihVyitpfskYYbUGZXWksNZ4GZGL
JaMS3ji9kIsEwBWUCcloMI9s2g78dbiCtYs4aOgPlzmKRHgLKsGwys1EiFq8iHslu5MVd/mu4WZ9
sXbbQcOpTLLb8XVRgHLJol6BYWDeOtRZuHamg1xv4Ln85bzID6hkhYjvfmvVyxCLbDPmUYyq6iTp
dKmWFDlAGpS/qTcZSwfufToJwZa7fq6gXhiWE929yss32nvpxazBweLi0Lv/DoTu2LxKWwuM7VpX
tRworjkhd/TL58PGFC6e6DG7WsbU13oW657qgBzNA55MsWlPXh5dOId9XwUo+B2CbUY9tzFz7SSW
aBulPpAUKaUl8bIFSn3e4xoqWqThs5bSmBjdl4BnseH94J2v7TCY21hyrTZrWVkKeMJgXam7mro+
hagkR6I4ucXDSaYF8ZVhUew+TIE2BkggIJOFEHen41MulYeqw0Q9djYzmDizd3vH3+ooH5kV4hlV
h0Og1lR5iJJUL7ZFX8k6irLzObQ9EiBWoNGlZ2YVgOMzPB1gBUI3DhLTrSOA9NU4kYo+ATwZ7VAL
m/eK3xA8cYM8lgsTc099OTPUjdN/4gPrE+uWhgUe7RXDv8MH1ct5Gos05eKAohs1w7Va145F7VBM
EQazEEKbAJdAKWPdbr/4EJwxiJWDhMCmaiKOVbRD4XAhqbrGINxitkYtNH7a2HsRgpoMul0/pbek
LTb80nS5gALTWEhgkFq3+M37/SNDxBEvtc8XWPk/oLa8Y4ndWKOl9ky4Rsd3RIo/nDHMy9Vaobs2
xiYDHsk+lp1+hzDUbBurMdrXQm1anNosd1pd9bheYmszhf6qb0TtKdz7d2XXJvsMdNvkrIFkvLj2
wFLQsLFQotNL1hiPBvpwMN3G60aUZegRFMf/HfaeF21dY4+8EcBUphhTSvJjcZnQ+cekJZVKM6LK
binPw+C+6H/gY7ueHMCQgXnptIBVBdkemJv90VMzqPot7sIPhN8Pg8t50yme+5rNL/OJUHU0J5lH
Nxdj5BvTxVNm2NbNUOm1LWZ+18oyzavRhf+NAb/NQ3/ZCSHDKwJGPsugQCQeFdS9Hragkq14bOii
PH7NaT703vWv2EpsB288VOOCapTjAdFZmp24jNzIw4kdz2U7bdZ3V8OzjGkUo/ZVlf1NYHOXn+jE
cbwbo0FwmA3A26cTo9H7mGk7aoixcyUE5MJlklA3EMeip91O9zkgHkCd0hdXSi4ppJN4758If2DC
yqDPjVzxk0YPEznZjH6SNMkfAwgy32jPOOd+e/m82msCSFVOvcTGeU0lPVqvU95VRq76jnf9Gaq/
7FCLtpmGd1JKK2lv7N6JIKKw0ELwCyVqPRqwJgzowG0IzfNbtzcliBMfZ8cgFCIY8Ev7PX2slj3e
JUC5b4HIejOiWP3cdHJ8HBqm+MLLPjmCiJqXnuCJXnQ1ZB+7eEpB4dcaWvHYbRKJUgTLyjZguZTu
KRI4EvQLJYDdXUasghb7fdAHdrM775chzkgaMo+ftc5ZlWTF97hSH5Rry4Rt0ajYRij2od2IRu80
iPkaishxzdBQoIZ9/N1DPkgP72GskZltQERPXoFklQ1No3xEFDFyXnQcmUv3CJEX8DaOWZKgaEcM
NwmaG1ePfuBDWW9urT22hnjit3UA7eD/KIV173TBOSepBSvS1fSXSMMYeB4VovUSAljEWL3HSlkz
1qRoKX9B0NIqLm60A00tHUtG4+5GPF24NDG1b5k83oLNobCh23GB65/cl3lkwX7yh8czfW6TkC58
XEkCClop2KNb5d7cYMxnWnRschYEy82oef8I9sD3NJqMwb79tnR2FI8LGPJPmVV/Nj9RHfbOEqbx
Sz0TXjmLpApVlm9MacOFEyH5TknG34+X+QS2pcRbdBCNvVVi2wBxPajquo9hFSw5eipoHljI6NRL
YHqLhF32z4TiaBHAR+LVOODIczZqdahUk2TYODj+AECJqqIsSOcWRljjLZuUoXh1cyknz/tyUBVi
a4cmzlKiHk9cHPCE4KkW38jXexh7U2kR3S2MD8x8/GrJCIjNCFINycnMwlbUc3cxETvv5oolaOuT
e5qL0z0K753n9MQcgLqL2ICwcG8v7+fBs/rQPGJdl8A5ldPPxyA2DqgChSVO9rpYzcM9Ux0WVoCU
pv7/lIfCjZamC6ujanhezFRV2YSEoWh86CbRQGz8zFVMVI2syLdtZDOyj/TZ0VM6hIHbIE8MyvbY
fspQdyyZxmKHx1NF0hpqrBNbql1aT7ac39IsgYmCpCVikDqMn6dknNDnp9nHKGiH75j38J3AuSEE
Sdl3fjNDfcCiYMTZuzT1qwsON6Gk/hhLfAvq0tUE6dtogdOjGS3NNLCfpmhiJ3ldoEcmnRm60aOL
aG9/VTceWrs92QOC3VlWlMASJuOrToOlFBHCTfGasmN+sqKhhsXbb/ntSo150u4MmxRXOeq8xKuG
3UeEARgZZOi+ufHSvbdg+2No4H9y6M3Mfj4SgichY7upIYrL9xHb4RYlfxv+8FtoxwLu2Z86/e2f
uCiGt3NxipCbISaf1Vo0DcC4S697jhrQvs/DAcrt9oEFTVxkXKXEYTlxkmoWGD9uBWlwHGm/+W6y
fTCuKCGCDhttvJqAZByzduOGqts4DFVN0wgqD24m9zpDIFYjftRgAIQ5n8q49rw7UrGYEi8cwtt0
VgZD2yAfbTDVnNZyo+eotP4fvM8atkGA/Giq3r5yNMfJsB/xEOqfyjYZkqlwbhSfuotreAcGZf0o
mJnbLUicqB3qblLc3fE3Pcj2BIi4XCs1d7Pg0xIlv2LnWrwYNYd/gB29abFLXdlZTiRFpCeCAyd+
vfonW/TlCMgwQUNN5+o4fuYpoiuzSoUBxn7qv5hX9GEcaEnKq4uyCnoWpxj/3GuV7EJG273UQbdY
gPVRlONuww/hBWdkN9aOJp8Oe6lOZnVmY5V2VEZ6lYrcUPUCS/aFHsPt65BMcmIUKDGCpSkCqHll
85mdJFbqvQEPKyic63iJjI3UphOkNBtxNav5QNXSEF7vs3ir9b97Bbh9xP+O1UPBOW8tjY8c7Eq5
XyVaueIST8TfcY/fy2PbJxIvmnGbRjcdzcms2O/i2IsLFQxm7qrAQ+Xc1j7RswcxmcLTRWvr1vKl
vM4xleKJU/D4Uh7rTEdnHl2fzfE8DxbSiCfxdtLlhq2isQy74Fd8a91Ywv3RPlejeNwG9Cmh1LOj
WstrSkaWS9eQJU28Tno7y08CjFWYvP0RPQuvKgH2Kp70Gxsq7NcsdKHr4JeIgoc3cQPDI3lJBrxi
3eI6xNaNVMoKScrLn1helw4JLg3rCO455NvnCOGuP6zpzeHMIti5CiHaVH9j/afzYWUa2Dnd0cmK
5AL37ejCNYc3IyHdNAIoSdzQ+4YDnbgu22PnDc5Y4lr5JNBFxuk/Ay6nRKg/er39Ql1bmBj+iLx6
6VpuUkj2kTPXEFQH+SMOuFtZ9WFZ0Hjcx3muG5Jd72mp/83YWNLoEoTAQXUta9Trp1bSJM3sgc0A
Z8TnUdNOkW6Lfx7gZu8BA7iWlkhstAL5abQttaPhoYhwF84MwDrnegtVFcD09ojG3Haq9cUeib8n
HM6GeSO+lqjyD05fRju0U/QBD+2Z3XBKh9SokH7GkC/m+Rn2tcaEqQaWK3Oiu1jUXUWozhor3twB
rRcbeHP+3Zq5kfdiVPORxCEFeCfGAvlDMpLRaodrBfeCVM/osVUU6S9sEDUmI2Rt6UMnEyRSpxz0
X4SDID8MZgW24Zlf4mZNRjDAt+1wm9yelFeTkGlMj0+Bsqtsy8hT4IT9r2IQtcv9wC1JgsurJGpP
h/AtAikALTDdfpeJYIMvo2+NxyEQ9RZ3308uO2Uwp/XsT/R/NkFIbIMQ7ql+6hUGVkDhvrHpX3XZ
263enz3zxtaI8JlGOJNUKMXIfAOehzyE0mR+6zc8/pP/2knXCFFXadZkfqHCP2boDeHmluvIk/uF
U4SbOFexUReENor6mq2tU8428eVQ1PT3hUTLb6rKSKli0Bn+Bnm+yRJyi4+IAtlDL7WPFKyi+lp3
NljjacL1yv8YxViSpFcbfvMFWwoXU8i5bEkg//7u0GZGSPKaZaeBrKUKOxlkfDo2FGb9eCd8h2IZ
qfvydv5+HBmDTlD3RkWX/bn0AC3yXLFZhOKf88j71zsTUyifsm3SU9y/f3kr8WBtP17a/AOy9ct1
SZ9LPxOdovMW9x+61MiCAT3FDBhA7lYx4Y8U5Uk3WXQuaa3J/Ks2J1DwwVDMS0MQZ7dO5j71qkqr
ccgQGNZcdPzw8VmG4A8jmcoej2z2WROPgPu62nBGitSNCv6gp57vpz7Qsx5y6TTCpOk2880e4kHa
BpCnZMxwLtd1linoEz924cdl6BBcSiA71WbDSOzfOk1+zj6uTiaXRWetylyXmO563YojGU/H3u6e
3zLdpRWZ4UaF5sm93XZOe9T2/p37fffUiVZ7ueFZJa6ssKkQT+/qWAgxhcVshLj/nkxMM7VZpseW
NOyeh23w1KyZLrJ/k+zQwEibynI+N/u5sgmDyt3Cpc8j1B0pfuFqfUET2RF1Y5C/8PtD1Z4+8EeL
LX5bEOqWMWJfV9Cz5ZCYaS5/lGeXhCtJovMkA2JeP0LVsaoo0tCnIjRaf1xqKddzkQYYELxuLMTF
2E4+VvDWLDV/SfxOU+kdqIAR+PtTvLaX5vE0sRhSllu49CaPTdbdOLuSxkswB3nakC0Ya/fSJuei
JF0PMf49CA+FJUp2jAiHrma17WSSLYGswT25zH6Bn7z6ju9RzUKIhKNEhkAiZAOr0kpuoSQVVtKX
2JZ+dNFI/Mv5OVpL9JUGIswl9xIWDgYIVCj+38aGQZj9EhtoDLhyyVp60lStjm2kCeNUEHdYpmUe
AmNV7Mw0h6Izd+PcWgkDzLufh633OiE2lJWzDiS+FDVgAd8oGqbQO1qIB5/loHMZl/YEW96Q9SU5
DsPXKP7EP4pRP9PsHjYb31MOOtDtdt5p5KmG549rUojMjGo1CIX+z1o7cck6lIjrMXhPfTp582GJ
xoz1TAa80HMAkHl6iV1yDXW0nTWgKtzOwP50mkF9nA3fM8kGRYrm68SjSN4wjL/2x7Tw10rntgxJ
YymwycPyj6RfzM7iTD3B5ExWcWcX5BVeldvjvxEFaja8l1YFYfbOKHTc72tGuQWIFjJs+RoWMnkO
x0tekOQBUv1fQcFXhXuFkz0APuaNytlvhuPrLyJUOQU/jotconKvTanLKeN4nNWFAVPvxJI1WZva
G8IZqlNGKZmQFBl1ReZ7c/g3lNaUUxtr61n0L/uLyLns+HQevOQEiR6TPPdOLrK+RTqSv5gC8ufX
hCDbjs8jHgU/aoOBgeDAzcdf+I5LP6LV0mYpy6lJiaA7hqL9yYncxz5jz9R/FPVW0+EUNrDFZNzx
22v/kQuGiB/adlGHArCQEZ56wghLky75ykWSLy7jXkO3ggzL4M4VUHwHNFcLhukYITS9+kKIZ6uN
KHg5q6lklAC7f69LhCI9ELfCx26zBo+b7zN1SPJrnLuNpWxmIX86SuznsFkhRnzEkjbMAexSnlnz
oQ4vkgkNhpGvH2M3k4lshNuOB3sTVBGcrvynQsGp+v85S1ChEyNSekTdwGODJbdagljgf5TLSc2h
nXvOoZXq3tp+D5u0evwVK7mYKuQfb4FP1zG0oqhZiRfNGR4rC3JL9Wzw2HhjJ3chxFSylVBwpkE+
USYL83zF1X/zf+MRL0ZIhxzyg3WeHVH7P9VzjI7WHw5OuM10JWxvCO2O6Iv4MEYBqlfJFjDLVtA7
s7gTZ+SUwoES6ol6WFTo2o61DnetycpT3U8sqRrZiqt2oDm4hwhQQ0RFxjc+1rWUrWHQoh/bbgoH
KsWlYlhsSW8/BKh3yx17y2K6JGlPGNT2fTuMLMm1IbR+QEnZaoUdOL2PDDryaWBOYGIimxyWMhr7
1Mb6zcxbwh7TAtV7bZ0xJK2Iu+tzM235Y47js2HqeY1KvRhZJ49YjUuXuku3Fo16mltNVPFdPWGB
JPdvgbvM0QcCMrftvpKJM9ei5J7REal05EcRKffZPfx/WC2B0SMYwNmlp3UKPRuKnrrAkOMbrsOG
+5XkpNgEIR740KVXoTIRnqR1/9/wKPQ7MP0MPOyW2mC/lmu8xGObIRxZodpSRDy5RtlUhFnWjs0D
+TVOXh+1G8Y6XHkFhuoaii1eEdnwZMf3SAFifOk4rAn4ff6XTFBZY8XmDajd9HvdEUhvkSV78TNs
it/q+z3S+ajYVV+6rLNTq7grjeEXx/mmX1yopI9R3tEbEZMXMUNBGIm0qYRuucShMvcOgFhJazf6
JADG1wuMzrDJuCWCb0jhHQjN5tJHFOxUCZDeAU17Y7C2ML+k4GDflugz1V868a8z9PItcnkmFqwU
drpQecTMzMmDWFiGB/+UGQCKT8rjE7t6qriZeB3qaTN9GfKNnXo0kNZdB9XyDEvcQST65UQmP9AO
/9VF25VeQtNl5TVz8kkqLDMdSUnKOAXrZQgMHajNr/nJJwB96EjU+JlJTqtuCvE8Bk8SuHcS5MC0
puelrYNCg6LQnyHIkq9A6xIxkBr1VVx1/TNHrpFibVkBJCqsQL3+bpFCZYP+bQhg9ifoox2U+W+U
WPWq4XIX7Z0ib8qPNyuvso40BpcNpGT3vqIyJ/uHr5io626evSoLOWkRqUluB3DHbZgLWcdSRXE/
zpcl5vDTIP/RGBsXPoqetdd5RfnwTYvyKWaVjzeBglBJ6HEthANY6Cd0sJLk3pZc6xKHgHMPGXWr
zJTKR3eLr9tiOKUOtlKN2QdK4xi8DebIbkVw1cyfd+dnriVy6np9Qkqzs6PYy9vBYfgO4zPPkMer
pnQEZ0UYm8H5Tj16D6XGIEfuGFWfgODOVaxn5ihnWlqNcwdpjO7JE44gbIvZWYKIsc0CbWUn5pAi
m8B97mGILohrZNsVLypVnvmv2qczPZxQRGHn/axx1T2zcgOHq+T85sTtt9nW/NqSQmFLBVIgA4PE
U4QgfciNvUfrt8/CzL0yTiu6MMLSUzUQ+C9r92WAQcSmZ6+otrZevWFqkjMYq2iEGL8fV/O3m79l
RGCrxS27UUyW6xo6LqEK3KD8f7QyocspL7d0Etog8dkjMi1ULlyQC1IrZc5qYPbSQpKFNWkqUKIR
6wkVDU8FjwjqbygT4tiKeK1dvKtcK5vQsXSKU+dh4kU2KzwmE5GDYnLq/MGOlg6oGeU7qEnPDPqh
LugT6Lr7t/9dsLTtVBDj9xVrMM2kdalZ1GF5aolQA7S9JmPPcJ66iqSEJz6lvF4wVye3Kz4usl77
o/uOhGuRwp35ddJgQoHdH7l6ASIjRyHtAuVGLGRp+Y9ZcrijFwhyuJKOMjLuJkvI5iowT0+zuP9K
t0+yHJoxaYObeBnvmmJdhsPABwDpKHyZhOnMJnvtzOu3OENtfs+mVsp+BSBUzWTJSJemhl2uiuqy
CTPm0f2L7/q9hL7p5DXe6/4IbnhQR3ndeYEM1VFi2dPb68szuarnFjOhmC5KCn2AnlkdS2+SaqbW
TPhZ7KT0TKLfh/Zdg+DLMwtMb406SDbW9hbk/QxfhVMhCPZcExUs/SGBH8ID5gpPnsWKmcRD424Z
yoFglpfZGfjxmEFKlVwkNEdrFTr/bBPjjniohgDOiQ0cJVXAL+/3bVrQkpotwYKL2SKpvkY+0MO4
VMBMtbbihRgJ1Ew3vy4Ebeo6Om7bipPFKtlTKRGATLymP7+Y8EdhiBZ05q1bEj1cXpmQDmLe8ENG
MerXE1yQ9SAZhySj/vBSkFnrztg203tkstUL3FVTkh6U5zbrSMBndcAhSNlY9IpeEMn5883ecABb
rE4EKgQoPXQwMHI92R/FJ1pxpgkLjQBjlW8gaRvrgjODYTrZRV0uXgNPQC/VlFNyEa+PXEvqO2Sf
OEpxnMKtjnI4QbkqVnvd8ecQAo1Gi11FwPWVDACIv3VHyICXv3NwlKPJFxcqebBT1Hx5TcfPcv3u
5od3lXD9iFJQHdWK/nVtVTEsGVB10Hqx5eJL1ZhfU9jgmq0jmAoqtZITfzXX2ZyodKji2NfotXOf
cm1utXqZ2cu6fDhNCFNU0YpPtSjEwiwg6mGPOtzCim2C5szpcKAE9Lr0zi5zNvTCDgOKB5QBsNvr
UQ/fRHzjZJeDhDfaOab7MifOK5j6Q0UJrsjM4mbumNdu7AygBWqm+VQbx6aLGfpNQGBk1OqceCRr
GiqXX04/jVsYeiDmO7ID9w0oNgM/7gOrmz2E1nI9eGVQp3GcUupBOXXq+TrvB1rJemcMZsihzzJx
MOdbjMK9jOosb3pJgARWOnC7hdzU9TX53I9x0SrWJ/AA2U6upPWgO60oWjAbKYSpd+r8hTG2lIOD
LLLYbqrMpRYndw6bL7Sg746VoweIRcCUUoCiGNNu/q6D/WRxpepf+qm1F/aYpxZBNJn52fszreMf
ZbOsEy5+XLVoudspl3GyCNxDb+ug7x/LGeOSG0D8zCEY+DRjHtJ4pnBiiekia7ix397vGFej71wU
o7g9Q30V8WlCjc51218hkCyBY7wLfsOo9Ms7vla03YwLMmbZF92spPeuhBQW00k+hZaLliID2LTM
6lum3O8Pl8ZJYS1xDnTbIhCrdUO1+ydD/RuGjAVQzmzTdU2oIL3KBPl8So7gL7NFBdLdkqkB0wzq
DETjei04o7vWRKVUDTzzPn9GhOdPPA8GkRFWXtxu9y9UgDk19Z1K/0jjhoB8Uv0xCu1Ef82e+kEX
PkZB28Y0t9xET45gZlqwNGBQqA7NIXNW3KljeUGkh32r32oaStRCfUHYqJzpDCFPwGc9n0N0rsd9
sh+RhzlzmTV/LsI8Ls7311IP8mzGzYK4OiNt9ckpNFvQM33mfzzxeoebQI3Mzw3+bqq9J9aUjs2Q
iYI7/rEl16j23nUQquSG3o7NVeBZxcDAwlurBYzkLfnzSXLK5n4zBsIELbO3TufMqRROsvnfQu2y
Wf5jQaW6woBPgtRfgu5BiMQorM99PE8Mq5u6ssqoa2Wfsh5yuksQko4hxQT2aKMjHK/1jKGmCgBG
ANdMaRCm8V8eFTaxqkLNPt4AHYcOTxxapBxzuMLRTBW9EtD1XZ0e6XuSQU8IyUWbAGyNesfYnKz6
hekkO2RcJTUQK7Y2r2sFM8OXOYoIKvhPqB+MXWbnRfwZceipI+7dagRQHgLz5nzKgXyg/4TKDOK7
PPcXChfA+lifL1aBkWjuJiCsucLvSy8mIKzBrXjGtwOpI3L5Mz+tvL5+AhfzyzJ0EYqPB0qJoflo
z9qbNgptLX4v7a4sajT1m6PrumfuI1MzZSmZVHSDftpgiwtq1JpEQC0P5MtzJ8EbmSmZAdQ6v61E
+9TkPBWOaFXzKlSZrszWuNbP1+NI7iy5bQTaCy+64IY/Z8XWceMZpN4Fn1sxblPQ40xEz/BVTUnc
8NGbePCPPwPxwSLhEBSztBq4Fy0Yc0KnJjxoCLgycI0lGxMvFqb8uleu0+5ylf2x8kKDWGBhLaRT
Kk/7fMUxNXVuIY7MPHV3+XJ1iNsMuGumgW3+1GYJBi+SvRBj6Ka9JEr1ZXuiPf603RyGh+chZlct
4Yg19n8OyR788N93b2FkXklFldGKyYjEENpDpuypJah1Kc8/KgglJCIvYZxcEhAor06bryxKSolY
TaiX3mjDM5qaBWVytB1WxeUh7VoIskTYXXDo/M/o7zQeDBJLCVcZU0ptkbyW7wno4kp94O9IxvT8
SttSZfgof3DhQt80REAf1qhuqYc781FjKtKzRkTfimWc5xtoEurv6zOFgWqKrNVwt9Om7bdSS5lm
XG6eGq5iGLQGHBx2jYFFbH9lZwYTVn+YbYKiFXcsjEgKigDX5Z6sJtzUIr/Wjt2QScbZ9fLr6BJo
BXP/Dkk1ffh283z3de0MtKgf8DwoDPexOQbzlOUYcS6FhV3udx7FEfAi7yd00WzPyB/1grf9sXGy
QqdNe5IpJZ1PsJDWaOrdJyDksbAMvx6vzyitPKGHs+mJxx6TZbiHwhLU3ecOqvcZjey+2YXArsEs
x9Ph6WHlrHmepZObPLzRjS20oW7pWX/uV8PMv0Wjvcl25M8yUjvx+uqvpL7iTD8E2ehP3ucR7mqv
apbYmTM1YuPHzpqlakbweOBkP805HevIJpMv510HFG4OA4oWNVsnvZeodFkDIe2oQIcyhvP+AX9Q
bLbsXTQN9GjTx2/jbyVHfunSFAtD1ouwxTIaPzSTGusJEZWiqbz3FXJCFxCaKefYQ74ONq6mJZUp
lSZQpJHYDzvhxy6HtG+p0gRy9NzcsyOOZyQagp53bh65hGXGZG1zDn71Sr5TVm3jiYe98OLJo015
tI9NnSynVYDJMBjyubacykvqQAt6W6LgszgBZ1Jri1A8S7X3oS62GLVs0jCmJ82A0Uy9cAN7mi7U
uTmMLarBdyI6YLbTW+jDKGgxKfdHdc6ZSIUpeQw8CPrt3bLh92vLLWWutqKaRPG4r0HFkeR66PFS
bxGhk0REub18BkXfkgHjHUp3AO2tu3etyOaGOB2b3mob+QOwZTIHNvlvtrCGtV4XZPNJHo6FFI3O
V6JwuUMZqNWxJ9eZ3xW+vAy3kexwaBhgGO9/Hnym4HP+N2JRxcQmVpksSDl5Wpd+4uMaws6hJ6ZP
vDX15v+xtGZDXLWU8U2/89FFB2KC4AU4FWJE8WoUQOiLIMOyLugNeOsmjpnsB6GUy78WdBYqYCrk
OznbEcPRtnuZD6Lj5K7RWmuZoUYJFM0WCDVYKYTpOYLgDn7//oIpQiNGmILf9zpCcHOY//RTZJAI
Y+X524T5YdUxXdjeBKuYUHVVGdl9Zs/yLPLc8ZHaYoheiRcVCLVJOy3TaPlm0EPK22J5nuKGKLDX
1SdhDbkGtdDFBpo75GKCPwdzQtcupcNjrOhzqll7HFcGMZglV4mfddxhKJ2ofRqIV8mwFQcIWWUT
BAFzN1yQTSgJ1fFeS39wgH4lAm5+aq3ujD4lgJa1l4dSBCPL5pmbizvEYPlovz3+jDJ/ofacEui/
mimWLf5x9Wpb6wuG1itv6Afm+dyADbYHm5kzW0vJWfcyovLK3Oqu/BvgCqRIh/VtoYOOVUExkHuz
nibm9w7JPHxR8cMvaFBgijtj9pH0zL0KtNpNbxw24GcmapX3WO9Bt8pBeNx9pQrbzr1KH398GaHt
vq2bM8SXBNfgeUjjXOnfXnYIHpb7QMwOcxIcjNGRe1xIrWmGVGoqWLZOpdf0WeUpNESsvU/dfkpW
NjjICkJgrqgG2nV5L9jnHQLj/ahA9syknUxi2db7XT6qLn7XQ7Fe4QTwuixeJjmM7AAEBVkaP2p/
C2ZAEqYWTRhQ3Z2UTlH6+vTY1/FLOqhG+ukiSjru5PXVLQ2etcxS19f5x28U79OGAiXu5UNJNi3W
heckItG2q9VSHwl4uVe4iq6GMtdkus8gmfgOBMXLfjETFZ55AYJ5CnqeUjyicGxF9w+i80Tgl/ok
ckuPlnB1WgeQ5253GfwePgVyguGNjX84aSMJPkRhVluW1KX+chLYrkAcmn1ZBRWXezb9T5Cnqi26
05kXSe0j+r8v29unyP54QOfWrIjZWyqyzCojqNq2qpCR0T6NY2zOBmUeBKfnd4tt5FQAB/V5zcET
aKiOAqsRh6fYZLyUlcGOJGY1mkmSeHU0mtwBWI0UKFJ5hNNGe0HiAztRrr9GJAU5JXUMIbyyLSvd
lmTKmM2TBOBtuAajTgSNwLeAozH/exij+QADFkl1f7yTzbpFJlOJ9g0xxgxmSRnsV4mDUrrmLpME
xsHMSKTCcQeJC1YUCa6HHUjBqanqtNNr8O9tEUZm8vfZSHtikbO6m54+AQAg987GpHKr+3Vh80EQ
QrtCRGdOs6+RPbpuwPQOiQ3bLH9wXy2i31qwhOiHm7q3CmaBDf5frUoqbh68H/b2U7IU4bbAxTbD
IV6+SLqf1c6LmXm6C0yr4N03fYAbfjhMXZKfHpHOlN+591MLYlWDV064dOMKyaqc9fB714K/zY1y
boXjh0wy4IaGujlL2bKjjgP+R9UzwvVbmuw0W+eh/jkDJ4aaSQp4YUCSYCDWi2ahLbzaUWxv4DEM
NXJ/ckFOJRCnwsA9Sqj0fkE89sta7Ho0muBTFtQj4TG+KTKOpSCFccDJk0uHK611+g9ZfB17Xg/4
Ce95/Lh+1nSVjwrRegnMz9dYP7IunH04PXWs0Ym09DROYXdgvpO7RdcBlvzAzeuKiin5Sw+JnoSJ
aVllJ8oOY2h5qKUrh+hZG9mYlUQUwaQwA+Wktu0j3U9kWXTESIEOlhvSSVCFWGwXPkM2151TFAe9
Ksts4wguUEGzwtDHtiGL1PlSYlW9y0+Wty4ezGyFoq4yD7I17qjFxLbWiGipzBpR39rzPkIjdZaW
5k4i9c7p4JAc5QMkg8tJAhpHRJbdIOVQkGXIv/oAhk7Mn9eO1/X16FW3uIc9Y6UBWXzf5Op+4yLB
Pbuu7WHSq4UQcjBIGECTnVFIzzksU5qoe4tJcYMvsO2uC2opcbxZ07sf+Y0kRkpQj7WEGnFgIsbJ
IEI6F/I9jmF1pBRs0tEF5MkXO6/NC035WjLtR9kuv0zsau2rOOItaGcb2BSwMiwsgAjjqZWetc34
Ulps9gGbkLGkN/G/l80HVvb2/ectMYiVxgkWnAR+9yuKEPaTrYKejZBrEpR64x6S2CuM8J58lBSM
m5a7c1GoVH3Z6Xdjt9DnDp2Xwv6T07tQiy0Z9XWAxdRuMlBpeecKQytj792kw3Hiz/n2mTzk0i9l
/XTRUmGkA3ZQCRoozMGK0WU+o8kz+HyuabffQiyTIRw7IyLRD4EgtkcFjz+lBQOmsy8KV2uX4lhO
guyDnaUEDQ6Yv4bP5nMQh15dE2vbriqxdpZxJVTEWixZgDX7YB/7M/3ScqCoGLF67fGUxMD3yik+
J+YnaKJaIpcpLLDYDMooCLFafgl0st7H3jxZ2wqSwdxgfHJCifpLhlqCr9BPZQHiIXaI89pSwuPn
T5ktawecob0L01FvmauMhS2q4CT9+OVSqV4GkCck2YI3WcLWNhxcEsCPHmHAht/vV6NRZJhTgF7e
HfHBEFQKtuWzJ34JBTk5TplPdISuGMei/g7iGf5r2P0wLkDane1eacKfYVx8sgffXJQbgTp3zSm7
Scc7e7lhUx490BwNRRoVJS1qnXtUuufWdew1hNYNGCe15fzwq21psDxv3FbCV2Yq5XfdHG5xwgGZ
WIJcBh1Bt2njDrlxEF9r8vVsK9H4iX93NNNQyqv6GKRd4FExHJqMV97qE93RaxG4f0rJcbTEXBaY
SvUAKs2MI8mXJPky6k+3z04KLhdmvLs1bxG4R7dgndfthJWIBI7RPkbNdfWqNuzC1AoVcUQOFKBY
gXDUIdAD5rj6hwWD7ZePNCJxvEJJ9trMelM2XpmJZ1wEsr2xQL1bsd9u2HqC2iSwGHroLYIdRZDf
AJcayzfAbl92qOXbRmzFyFlovAm8aKOFQKji7mWSN+h7I2KNcK9XlNvpH00p4dgbiBMd0ADulyQi
j/NKWyIpyCpUOMTZ0dslwl/IPBUKbjDN6XLGgOglEN6CkZa8KfRjvJ2mRfd4KUuh22H4HNO6y2m9
P0bGGDUleUbWPFvA3Zo+J6T/v61jqKDXCTuPqRvyu9BElFKOh63b13oXjNVEVKLJF2e0fZtItkRo
LBd/cj0Rh/nnoja1LN0MjByD2WNJ0l7STsoghiSKgyXlVF6PTKaqtnVZXVzBcyRKDSEkHNJR+NIx
ypppavq5pT6UNeDLxo5b6G66DvyoUvdyK4AKm4bmtdFDyAAYBdjv2xozTmin/609l/hZgjQkkY9y
M2hBKHL7IU+AT9GJ2AlmaEkaiVTJpzCLMDRzCJfoW6nENolgC6LboQZSLUumPTJVb2y9hADDrEVW
BXXyEuRRoucBG+Y/FjyYQgcGyA9PMCNRDEl3c+O5yZVDsh5qVC654HlG6GAKivct/JqJl5HhyI8G
Hsy4j10s6PHCruh/68EStVA2T2ZQJobEgWm+PgBBVhwNIAMI2loQibXh2XAIwCCCJf/1MqtUJW3B
xzkNxIZMsMfNDjR5qnv/Ce5Rf+JEJ6pvTcQMBdkomy9FXtb8ikjhkBuqB0NZnkU8ePyaUWMcnm6u
XudUZb6Ol3LfR8CktCgPzuGfCbDhgchZ1mWCo26xTQlufD7e53nBHx4qfmSxTIzPWS98EBY6tSrw
dmodmmE5GjfcZHH+w5/VRv5lkJYsWaWL8CBFkIUhkxBHyF1xQrN9+DcWr5x7QB/JOAU+ARIL/3J+
CSHSyJE4Awj5LcikAANnwetcRtJIEhIaHt4RXXziUjlPt9wpOBlU6U7BcIKFdbYJXkotf3sQ/8l/
Kf1t7V5D/HmlZHPHGRYdk5RWbOhLz8BJHvdY7WPJbwiXvZFBqP1HmDTrQ+zlENAE9lm3ot3sRnTI
RYZatYNKYLay+3wNkzIoKSP0p+OjbBJQcJA4JNrDAUHKFfV2ZH6/3Vwqzb6JSDtHZm1/rOH6OBxk
ppX7HIydtQseGqAFI3QRGhszF74G4gSvcf5CdHiGzZON9qxvP2oxQ8V8aQC/82ds/deSJObTcy5d
/XgSeA870VjZdYNu6Gb81XXSe6v3zt987T11i4IgWjdrENZYA25WWdLNl61sZbvRQmL37QSAJi17
BkNzqiu2EU8W1PjedAsG8juY/Bdk3zU1Zj2mVu2LE9v0zzk2LCIOtc3MWGMq7KcC9KzzHpN9wDVb
2qDocvMYYNEIfjG3vwzEYIj0Xmh59PmguM6qeQ9EuNAAY3hhErEfiR6CwvAFp4imEsvwphkuLCBE
1JHyEjJzbXLTOb7VfNX8kwlNc9Q8DhUK0DXBF/GGqzR8UY3zLOxZIRhwotVm5QtGDnoFf3UKxgYx
GrOr2056CJTbQGyc+IU5TbNG47gFuSZ4VS9+qGpxVVWOcd1YM9edrTe64lSWyZR2nhCKh53Gvjz9
Z0yogMb966A8l7c6bEZXmkJ0iPoG/Mf0YvQeUN74lMBiw6rwLoqLs34NUkI0rGzTDjpo6jrEbfMZ
D3vdqwo6+jSRFOslZOCdzs6uOKTN+OgySObYgYIKDBQ+u54dFGET58Wi5FARNLB+Yg8hrl78iMxT
VfM0d62koXhf/FLot2eowCB29QgQEmu/XmWCvTI+rpoo0fIZEmN7k7T/SKExxn/o7+POa517MCHC
ooHoUUrBXEHpX51KYLSLpZ7Pw+Uq/HzJ4tfMWBo2vpKOgcyK8s3JGi9fSNwUwayO+xQJZRFnULnG
J4kVjE7Yy5C7OQCpeCSmyzMerOmtDIgeVkkcZp2TyeINrJ8ORIBJiQ+T4fUF1mxKjIvfXC8Scs0Q
BZM1pcwNVSDnnle2JOsYNatqu3OTWM9UJzG5hez+Ps29im3PS9hXnimFDzFXDKWpQdoj2cVgTcUR
eATM3UCvmvor3uCR7PplKauQvJqt1HvI26CFXfvgvDkbGvCDUI37uAxFEZFpXhOLtM9cDon/nfHg
amjMBHNLm5rIBUFOaj3sBeSM9I1tHrb6IgdyKQKW0UEPbFwqU0gYdSgk0VOfECEgz8vV1hLUsf3a
ZRIj0kJc4ra2efUr97b3/n2/IPuhctLuSeMuLEY7hsJGU1v1LPlvPmtuf+7dZBBUwZsEaQ68dUHH
0nNhmoWY233anyE9Jz5ijmEuoL3Syn3c/eZnxPxnU7NYHmjwVR27u93vlWRwdcvOV/wxsnM8qoXa
UY8YWB22QpP3Oa/Xq9mmqjATjb4bN6ERzY/Wa3w138aF8XUPAPnbYyWyv8FPopRjyIW81ldMGibh
pyBU1ottphEPv20ut5VQCCJ9DDFnz+roHSlcynMQVK9ssXo6QLDyhq9bFwfWCNWKRTF629o4VxBO
tN8YoqVKY1XQUBaOlh3Sq8aBHk3l0itch6azpmgEziFJ0Fs8tCN2aeQ5cpPpTCztEdqI3pmKO6Yz
1r2eU7Lh1ZKe7KT9Fub6T9RT+k7w8YdhmkEKt3bsAL2NOFsAbglTbcuMDGZx4TRQExKUlUnGhq3S
ETgH9pKm/xhMRXtO1/jRNg0hkBU7dhbr81rOPSqepdtnUo1g3p7du9TlvS11QS7zVN4/d101g66h
1oX7lfI25yCQNBuMkMz7QPlNbfvDsWVO2tgDONcqaYRdsXlYQ4l2I4uyaRVf5f/IJZDyUL/JhsZD
67f0mr2nr51xlu28d0p6hahI/ro0i86AS7okHss7FZf430pJ7v90hZivFodS0ZYD5lZ/SGA2qjGO
xR5VGdz0T4EZGkajL/TjQ18GN2yJ2nUwts+M8tGumCBzOnlWMgLxlwDRiYRfvAo7pdfzJBG5pfv4
FT9zCz5GiDaARz74AdtlRqH14ACYP/rXzzZ7ABrt3Jb7eKkTpnxj1SP2sbtsF2UBB8kinTMTT15T
h9p1n1Dfi+0AWIjtnYa0B0vC3KEPP2n6CtRbYyawsy3YAPANFepvrQMO2Bk1wGOcs3uJFjqpYp8B
Tds+ohb0o+WRw7z6ZXBYt8JjJA9zQzy/L0rVh7/ZBjt2lKP4eSQxPgIpoBEeT0sSburcWZvUlIY3
5XRsLt3toyCp8dECKLz6vVw/KUC4l9exOata34+Roq2PfR1w314LFNKCzJ/4uCgPyOgB0j1s7gqH
YzTvBYrpIajfDkBtfqf2TR/PNfIbmGnhFgJkBOcYqfWWOnc4WrPSYLonyMYiQ5Nf6uxeHOVVAXOb
eEQvik/ApHCEkOp8cfLCbvwQPQ6988QjohGiSD6LjBKZKRm/XAXHsAmcrMCcPJU3JC2w2PeaFVME
J14YCe6Ll31B7CfWPmWV6MQ1Sd+A31TAm27DnMeUi5frepAe0nA0NWPUtrNaoPffwfnfFb6pBasC
IT34vK7j7b+U+td6RSSXnyVduSc3IKkP9th1gtZLy7ejHwN/JeyI6wiaRsayaP2dvZlcXcrqF/Et
twOFsM2Z5f4OZ7+8BUd5OocJAFNfMIayHclboqHk8a/hTxZ7QkcdC49bsdBAVHH51mIbpAaUjjvk
GoYGRMrrIaWy2dmtNxt212mKdq8zFCqct92wsFV0YBSGgKNO8dz5QCRzYQOhIs6GO1jOcTG3t0/F
DV3+qxROppkIZs5mXo9Mb40/kEoD9LHqkkVqCbT+70BZK2TSr6YA4PtExncn0zqNtuVYkLurEDXn
rtCRvnMFfWx6/o3fwn+n7Fgvhu7VEO/O+o93g++4mko+0Va58RLUILQXY266OqRrhS0GFVaNJWgf
plx5HcJbZBkLV5Gq5ZuMdXKFhMqalmbq8rFRgfNHolYWrUoR6Hud3LvyFVZQgb2I6jzO3+NkVXWF
r/4mY8XCCtO89ZKO6FiHiHja3xB3Hp95ojWuCklgzf2wEfLAuE79aPvVeb/LuJKiIRbhM9FbsLio
/jtTXyba2G0r1JR1BM5BtkZzwovq7rvcAHKMs1uiirE9Nne9eYwdhW5FafeYhZhGOlGRgDBcL2YI
DxnoxLZP9FGmWy7dzTBqDfPd6HDjAT/YlygLVznhEfH37tFRoUg1SjWsapVJoXscnyftmljQdwUU
71e3INzAsxlQOrgpga+NvSMlVvJqorLPxaK7QhHqy2RG7fQ2aXmCYAMoXJuW6MaK1l3SUEDNQ4+L
xTU8pFa+8U8fluaR9OtlFB2JGzRWrNnmVjUQciKzNUUjxfcDyrWQJRVuOmWCeIBlkhgViG2pUZCq
erPs9p0Iy2y5iwNNFRcX2EW1xSc0bkfNWstd7x9f2SwokEiC3kLGv8EJidj2PcdKrRTHZ0zGvuiP
GsAqqZjiRyOVRY+Fh2x877aMZGLrnzQgHU84879oG4MevmZpaTeYzOnV6XtYtT+miwRFgRtQsqPP
KEgfUz9pdaXMifxrfGfOLHsOLT3bz3kgM4eBPfahOuoJszzzhXOH1vvGbFncks+1RAyXMylPfQRv
VknHnGG5NOuXaRvqJTPREBb/hzbzK+rBji5XkWVe7qvmg7ZAotlBRKiHooouqQjxdk85Dibbq1PY
lGw87O7PsbHO7umFeohkdzwTnpCcIxL/Oa2ITLaK0u14/sk0pYs2M7WYOiIYMjIbYvnIjaFvJLYp
U76ML6dHBg/8LyFnlDT+sisw/Be/iYGKH/H06MmA3VV41QiRYzW4mLkam2SHOyrGY+VBjobrf35Y
qIlMjcTEijzYfpatn1NUMU5LGZU6DO+ZdnXgZGRNR9z6+fhfBFuhYDXW12nmPumbxSEZjr3b34tc
Rho7vWhACc5LcUl/j5+jE8/wS0s/J3FC7jnsPjxoFScNrFypJlfgqzucr3sE6Eg46T3b2uEUAIpM
n+lSbBb77wPmVB/U7U2LRhH5Nq95z/C6YebDSTL4o7pia4PfTcEAV202vi1fKk9/wSy8o51aVZZ8
uzh1pMuDTGU/WiM0bUf4cjYosykubEpbmC4d69unULYLXWixYa+sJ2Xxrz5wVbo7mjz2Ots7X1AB
g0SmQ0PewvolBvlvxGArxgygWQkhT5raSd61XInxdVNQiXeQCmTX9JCxHD/ukXZLoQqhVDlOtsyi
QsalwDbyJXwnXH3GpWA9brb4SU5WfqBvAwIsi2E15hHJNPpY7iHepaIVaovqu5m2g8LcuDx7oMU3
haRPP0DfX1bmqLEHu6uenmfu46M11pSrDpYoWbeHxOgoEWZ0bacrMwMWy3VxRUQpsYkjsK6LIDaO
2CtTUfx6fWIWHdfhYubpIPSjHZX6yN6ntv/5MSFoDQ17UMH9+qCZGMJY1NW7tkmt/tXT69nW/TmP
cMCoe6fNfwotG+tS3HUyWkl/hXc111zH+B7564Zd2+Tu8DlRFYNGgCn1DxokAJxCOpd1ScvRegbh
3UCKWgYc9kvpjOjmrd5TjhBXWdRmyV9UpwnGalF5O+4lxUZTL2GILjpEYCJmdIDb8GEVxH3h7ezL
cEUovLTzoxE5UQIghaK16o3wtIakQGHKkzLFTWDbGyKE7wKsyd2H83uEKKyApT5ii4DHeYZWUBXJ
9WHZFWDNOl+GLgULbFpHzz4DtSucRCstXBAznji2UEzUNcKyun8q4Sd5mh9UCeiABZiMuTcaiIg1
SLpCuUvGvwNz+dfmtz/cpW2HxgISCp7cgrc57BF4GcSfsJW1Um+fxk3T6Q2JfRlZr08ripybUT1I
BL0ypT5vvLICI9H1ySedr0qsELxbF8FoczWFD6BOr3lIsNn7pn+VCAazt0bdPrAfBF9tAyD1Zlvx
VuDnTBpaUFkFO96dgF0WMmP9z2T/dJvbgXHSoc0oPPHX7J9ZTPNcFWHdWDaooXmBn1lgMPqyB/6+
04eTM9SRyXOV2uclodnx/1A2D1Jb/FMWm/yPqSqi1/9nUtJhREjCZys2CTtITrDc7y7atwgZ1M22
v3fJiKxA83C+Ri435iX9NWHuGE7BXLnacxtGtMnHH700id4n8q0033rsTX2FcxsQIwC6RLzN7Mua
HSfsOMwp5L/8oIX5CoWh/uyh3/7RwA8/sQzJjGQjRXBzJAIREOM+wqtgkv2negaVLpzPMNTyYsGD
wUA2ECk8OXGTnDfXe/GSWEEhYAkDT/tx3TlfehvX7eWlIZUcSVJOnnRa+d3AadX6SB4F7h3DcLUr
8e8iNuucRlt4+yyybYnxnEaW5IQbKRkuc/mHnhE/wHvSwZ6dCZF2xe/V9ISTrg/mZOOBp8S01nBv
Vsl3cRrW0aSPUz8vZTOKUwgIjOvpxRcvuLd11Lf3Ljwi96V7Smw9NlcRwYziQ+89BG1OAw0LNoQa
WvNIJp8DErPnKgARSmJtXf04yfndW5CFMw7I9w/5kDa82K8h+wBACRydBuW6Lj0JmWFMD0DG90Pk
YYWQgxjeToQDygcbKdEU49TKaIoiJUeXXJBGWbcXF8F31yWdQNIJ00ECoYFWrJWbR+/PB5xFDRfc
wqQ0qluINrbilbaz+3MFaqqFWeUWkIVVatHhZdCb/l65gQJs+U81nAdUfMdzUAm6R7P+GxhBhV3J
5nrhGjfdRCXwZLQ22dHpnsZROsfFcWSowMKUzpXnIb0FWPpXuvXpMAk1yW9MWfrYew+kdVGYuElv
ky1YHyuQQuoQPwSKkRsAaoRuf4bUdwn7nXmzGJLE6FS56vCYJElhRGMUAjHZtGp9PjkSolx2v+gd
fRyXhXkasWFOc1Jex+2mbzoplzQ5Jv/roB6CFLyDn+OzySQ9LPjJCHVk5pA3H3b9GQOoiwUYu7S8
Qrje48XsDyUEeESBi7IfvdXe1HWdzksrsIlfKuSPwLIGc3QCu76sVuCreLylCggXhmSSkjaeCttf
LHbcLyIerxzdnkOmsBlRJX9cZ1G5ILhds+WJeYH156Qqw9/hZZ2eqmtkxnWhS0FakmuzJOztBFGO
2HSvcLRxehLaaw0wse0PhCsMrJEtFpIyvpll5H70XPj0r/BLB4dfeGIoApMlk+ZANajyAveRPEGv
aqZJpgdumSqXp1R9HjbR7aVRblNmN/gXuEYlSKahbyDaSDjEo/wdWunqDERDg61YM1F9JJ+zaVTf
wYxa+AXhqWEKyGTpZ7SvBjFwzqZixg7qrDB9RcIQHJyElQYxPqUwkjjMKumpC/dixCVH4Bz3xp3T
4NaiGV8bw3YFBaWBC4WWdlN2VfrviHaTosuKi53pYLmvrfMfoi4YDFKDiMflGskCqwGG3N4IgYXo
ax05ZpJ8ob548KRMwve5tO6DTlnVpY8VJVVEEVZPWLyT6rtIj8GXHZDKNFQlJDZv82SruGMKWNNC
EbvaKEJZADQ8sQ2fa+owdQX+Gz+5JjNnfhu21WCgtbcj4W5o12sQC3V0VIJglH10PKsfWVGhTGXA
qbZGjTwSd9zW6U/GVQC5koTL9WeDdttkA5bcYUqw1J/6HM77dgmIG711SiNC3eub6dsuiBpAjiiy
MAgLyJMuOllmBS75bnS79CrdaDxlQuxXezo9oxZMbEXKTFH6sntHE/x7FEh6hGI6LOrhzpNIjaFP
8OU+tBFbQFe15Vf/IVvd9wy73HZev2RHRi9gKZTaOc46SGEptYj2KLCzfz1hriimGb/N662zqWde
jcLPUsPLPQ8bq/jDCM6B6TQSo7uKROUwOlFm907EJWXHW1xUOfFNVIqXtm0h2AmVTl6mGk2esKMo
yzDMhYVzuZzH9prGM/CzpdyjuBMsqdhnGF8w5Pso2UORasmHmeBbiM/9fcIDF1n2wKryRiXDwOqj
kki8ygF5rNeSE7MvOX92FNvjUbY9kU27dIXyILWY3srL5ArjrGt74oCf9NzDwQFC3QoXHGhUjATi
H25WQYyOsSYAh3ZiVX/xV9VB8EYGMKnuZt2XGBL3H9o8v1yLy4g02s9RE2HbfEJFs0WOUln+t/vO
AcGpzxqEfPRABr21agiZXdVz+aDQaLin8KXs0FY4/znRIzGyIiWWeVaNJktg0+4hoPBdEU7AlYkg
H341aQiVu8RDinjMmUVqyS7N8meUCiRU6IJ+tRrlXUsHnDQF1+V+ySEpRprMb/wHcu+Dym+wVDah
HJzBJJN7j5Zm9ZTTLFykrzgYTIXXtAgFoiP8W8NSMPIKNMbRO6Ap3ZrTmDjCn+DmE5qaWL228DzJ
+GofSUoLlYNk1dsLE5oJv1RninCJ740t/FYv59Xg6A2DRsPr+5usQh0ylAEw+/PDWpYH06LgFX5w
1ip55mfMfcNsZO0tD9DER0SPa/6bCR+3JQBu/geczwrh1Gfq1GCGY8IIF+aiJFb7sc+6VVKDcfCP
/FjSAuib9LJO2EXVOLp1YfapUK2i85Juj1Z2XnEALF8RKAfeygAM5SnSW7xLUNruilQmLdvslcyQ
qDfbsWvt6Y6Xa65YCuOM4E9G2j6fUjcj19HVR6onip+eDkAni/kzXH4y6lCF0obimPWoN6m+aG/C
sHHsGNWm95KDkWE7eaup7YJ42wt83QfmNSGw/lnZZ+M/4nplyrdmPf5EpCyIVftep9u1HLTPwA9Y
hM40m5xj0gF3baOpZZ2sNLV/45sghg1zCGt+wyHnL7/WTXMl54Mxk9uwQTD4rmMKUXDb+3fMf54y
O81xTKOQBWuKazWpm0v/Jph9vyEP/WueWQwch/twiYvjV/I3GcFD9lAdoDZPX6T7D3IJi2H02rf7
+k5RvDXPitXe5bSXQThd1jrnCWr8UnQT0POkCfMZEraikjiFxjPPVMhXIiJli6MePIA6QVYypP62
6j22jFpbTxuklDVVUCI1dBxGhSdf28XxUtnKzJq4otKS6X9XlpYBJE7pZRIWGMUQX1xXTYtUTk94
lPNFUVelmt3QD81WU940RwaSA9cxyG7dYffZIYelHWDj2EXwZIf8pTT5DQ7SFxvSl40Jebm9LqrL
IBh7roodskOjcY4WbygKu5JyyBoUcJeAPyLxutlPHJ9Y8gE+RejTOLFHBhC4GjHoIMAZwRYVzEkX
tDAoGkso+LmDF8tHh00We1j08wRvj8eAyqxz/g4udgiROf/CpT+Qqwhuv45PGn9CI3NZi7UiflOT
mN6WiqjMT3nVcGhcVFgugr0YoGRN1INUnSsaWVpmdXdNXfPtvmQSEkJ1sUNqqsr/cJel/Omn4SUU
7JZuufcGx7n10mNJBCEaQZ4+g/ruwHj7uhshfzT4h0TGZ4uYElOejdJNz+pCFrirxKAQi5S44zin
m5/q0Ehrc6VFlCld1ayNvBjkAXW57Ee5z9ity6JaS1+1Mw4RItWS2wrY+krgf49RAA155sz04ZJh
bLpUOOcIgpUwINCTvAuueYWaxXvqLHzADHRzNiTj4T76pyqeIWgP4t9Sc77evqL8L/yk93OMdLYF
s243EkLJKC7DhFJgbImdYAN6arf2MbkVj9yFSjX8uXAGBh93QgtIU50otbPjpp5iEitHka0WxXId
1Phlk7a5Rt19PHEUbM6YMPtHc77k2q0WL35FrhVZI9p0ji++D8sgNkZ3Oo1R9tdJGhT80UTBw1Iv
70b8sNAeZXsxMJTwy3LV+LdPDkqWJu63H6js9Axi81dSLwVZbI62Lm+zas70drYC8+7pZX4PboGN
J+YIzGiI1ICno0xjlWgXRCYXRq29hY8ShIOHcBEsDZYgViHvwllb159HBX3CtFHyYrBnLwJK/Iw/
gftPpHj3CsRX19AYRcELwIAarPATJTnINpSZq8OSIdfhWkCmyNLcThixIwBQEgd+lEbNaTVaBiqW
8Fs/HkH712YGDbr+sJpXYJCt39UEqDl54rJxsa6q72Be5nTFFDM/BRtnUr/oXp+8npOP07EAHGVc
or/qN/8mMrDzKYsJx5UvDsapVfRmBBnMaiuH5DJu79BRC9VxhMeYfvoh9PoPONGquPrUWNprGiCJ
+DaMetPb+DbjfSEF57mdKOduiU7ED44zraQrzg8ceztaYgHGl6e0m9p1F3QK/9gzpeyA3HjysuN3
Dz5rjH58Ka1FenZHF4iEe749L+Iip6XfDrzfh5j8KKqSJL4GwmFGXeBrjhLD+IbX1fjFYUVQm2es
KesrGjWZ4u+QzUl7U1sFhEZg9c3VIIWZtiWG10aF8uILXra4b1LRtc3SzjTzaNMAZQoovVQyC4Mn
vm8EEmmGxaABsP2WnoiroOSOwoXcaXQzM8KvPQll4ZyJhoiRfmAJC20ug6fSJh8U2XYcQ/aGLKMv
q+IF24iXouopE6ESe8BMnAG3CATxZX7xq4OHT6E06ANlzsjY/S8+ULsoByk5i+Ts2TICnoX0lPqV
dZ0fMZPjwpfmpwWFHX8i7ibpGOSfWDlVcqfZzYjowrY6dQrK0wGnyE6uprfEMxk95Q1oNZ6rd0bK
olIaBWrxzO5RtMZog50d0R96ExTbCN0WmPBBsWLlsevI5YMJ9B/cDV6e9hKhHjw0lP1hEhXerICx
1i0YWXg6aF8J4DI08XF8r54YjJS48sZiYyDEwBYkF9ZTJvBfYemNNnBcX/U5NupmzHog7R8N8mLj
QoArmLc9vxWGKRWVuVuwIUiCLAV98tV6fvAGozJMXZRwd3njyEmr2zReL1uVlwp4b9bPpyrMZv3Z
iB2+/8cmWs5IEgJB9W4UMXUedzO+hDVIn1NhuK9sUhFhptKNfjDrPDCGt1pZpGujHskHziwD4Qw8
0QMwGJjdiCPl7D98aPpMNOgFxAjYx2QDzVBydOZT/ZvuyZMP1MEoGYpXN1aryu+JLbBYz4+vPmu0
i2CgpQYzzu/zUYf+Q4+XLE8QRGtVO1lsPGTKmZYHZXLc06eq6Bedr5zPBazbkr/GBh5HSAMEwS/I
P/Eqkh6fgH63QhkCRmkaaa56BRSkqTlEQRcjxTbz6xEl+AQpBZwx43C7JXi7ybQmvBrvLibLHiNK
siGUnx+6vYJEqnanCH+iY76B1W2ve8gZtZYDoFcawrmjPkcc2UedWhiAuXK/4ev6YMP2b2n6CWAY
11uS1g4J+WxLDew2J/kXgVz1qQDvAolIvyN4fxB5Skmf6Y8X25XHXWxKZhOQbJEkeNIJQ8xAHVX8
Ba14udIqb3+jRsikR3XFNTqEpqaaAQASs58Ag2RYtqth7rrgh7aAqtrlbSHOtw8ZlkMTcMtoxVEH
2Vkw/eydC6f6OaAW++JimmdHy7AmErrkWsbSfT2WW/QOtYRJ1rrSXUxUlpeI+2SIeZr0XArPuhAG
mtoYBPzygWePhamx8z3lVYEhROfp/CNEWaKj8TGDe9ZmvTrppTV9lKyZQPp5SieegnvJCRJnXnCM
hrB/ygURteoRBxeOhvll97lQfK6uMRMWufOUrW9O7+a4oZX2fzOGru62aX57bEvlPScSOMCGneOt
QHd4BtgsgKg6chSVdAs/uSwj4W8ytwD9TljiAIvg3qhke3wcdGo40lIuiW/WMiRCSvDtanltJk7+
e2zmdLUMSPHmqgO1XJNkBd+F25snhkftXfeb0vJRL3zOWKfsbQ0o+o8fka7FuEwXibGbtspzlnYG
WNRzVDivaZeh413QT+5TwEDa/CR9ZYCBHKP5MCnLmWlGjMLLuzOXgrlwn+kpoz7OABDWvd6FirZB
ub/HVZ5MeCcYfYT/UIYSOSke/9cVY+EFN50QHwrWDL5trGv9Cabq9gp0IqzdtpbPXBTY13r4EIVT
IUE74ih95Kr4ldHq8otL22TzTTD7FbnIfuwjXzHdDk6pYWicGBLx1R09Ecdim78YeRH709DCDjMn
rsPS7E1acoRvT0/ateXrPMNOZJqan8eyWGtrPLQdY0FzIXDUjnxStE9JUjYQRqe6/B19YftsX5WT
q8iYzRya2rt3OpCw/ErSx3Bl6GOE7XpHuWbI/a0tn8C7pOghdYmeCxdR+tkc5MN0bjQF9dxOr7t+
x12OFrtPZSnD8xv442schR9kg9vsTsGMPJU2QhtrH6S3eKja5d1xsGEnzUP5OVDbpcQ6TMjk3Oaw
D45xEYu4brJNm7NCXrTI39IZFdJbeBidoyhOw65Pq6vvwHfElfoxL2C/7NjLQu9FP9XU9BjVIUII
OaWIRQVaAIkLuNiCKk9USyGcW/vI3NJxTC0RFsKFpyJxSbE8zWpF/FXX/Xsj2LUC4rt18OK4rzlg
MEHNrA8Wdr0/EU6sMsVVou+L+XDibzshNP9p+7ecRzTDX12AHVYbPaCY8nFt3azLc4MqSid9Hulu
sto1D9PS3r/+i1pFyKmvD6qtdCqYZIqnIS9OcbHw20GyB2Wt+77XJ9BJTmwdwDsAWuOFRG/c0z1F
AF+ZA7nuZhCYaY0NnhE1KIPlSERwS9JbbCYmOcubUq5TS9dM6C4eZfY0a3TFx2Pc/EkgEusiX9tp
3skISIdhq0owC2S19ba0egb4IH8mQ5SZ5i7ahcBcgX6qrAUyXJ6Bldes3DDnf6Fkqr9VoXnRFF8A
VY3ksgt8DqHkUtCY1VXLzaohxpkPILx0A6f6Jc7dUx48kLVdvNFVdEBzMg8y6yrBZ63jH/pD7HlG
yG2RCdtjdLtdqDAxRN1VglpPaGFE2ZUB6yAv+S+OU005YRYFWZW5/KTkoFIh8irRy99lHT4IC6et
AqNph67Rx/C4VdgtwcwJzbgPtRZox5vbzOcU/XQCPZbNcI4+LigqCVVd9alVrd3IW1aMzBVOBhqq
a6xWA/gMXrZvllXB7yadGMHGchMGpIvOaTDb3jNcH11pR2I+HfFMB4uBmJuRTTKGDZiAIzv8Pjcu
YU0AgS5fiqMYI7xpP3HzgLz76/ve5gW1YDzihObWg7kGPdus/PaiboxiJyaDI1x86XZyW3/lklUu
dzmCdjWjVqTwvH7nsx/dqwnkelLp0UqFe6FzVrxNqsmw1V1w79seupn0U35fnVOKYakl6XZ0+fso
OPdUae8Ug1d2vwlvTpBksqhpM7p0zssgxRcCoZ7Y0lELSLrj+Q+JgacRJnJKye/tfzIKbz0lq/xk
jwQxg5EyjdeSeRLbbqagy1vWoPYyosg6rN8DxmOGkrBrGydXh4XdRaUiKL60zMgdCHfXz/iAnAn1
0/+mGJcOAHV9KZfj2QEsqXWGBGkwsC6LJ2rvyMdXruP8ELH4zS2zQL/1VvVfjFf7lX/wVJ7Jtp/4
VxcOlc+lZE/07FlQ+puuRa9DmtIUdTKOpnU6JiPU6t1tFfJpdq5xZoBOw1XnrFu+SBFaHeaVVogL
ed7DO406WChUy9rRCKypqDo4qO1EifBiODauax0W6VSJ0GHlgPU//7uz5BOEzbxEE4Ze1LXshms4
0liIU4JnSULD422ZpC34by3/yikHmnZxr4Z4X62AzwR/iWjgKe+3aS6n8wMG0P9Jf6xlDejftV+L
GHtlJ69xesxUeD7GTMv5Vaxji0AFDTm1/0i0KoALIQx+ZioC+k5ZrNjvstIA6D7/p13aRx8mDelb
+Zto6twQf0HirGj2qI6iiWARMsAhCXcJfB5ISt53Cuwy06r0J6hLQ9xRhha9bzsA7HUBQv4yTQiX
NMcK0BuV/sCPe8jLg78zkczZSaLlMF7Ah5uGd8NKfgBXYRrESZU65LyI38tam2dlQlroTRIkU44v
OUAloORrTUt2WL+BdIKeUAkyfzaG6LWGNwfH2VpWUm4fJB3RbbC9U4CrmSrA4+gOpzwwq5p8yMLv
0DJBJbOy+RIRZo2jfnJpD3OAlOU2uL0WLNeJHsMHCdxNPfuDs1osM83eBCnVV0dKIdJR2NZsuHhA
tF1OrKyZyZHyS0I7p21Wxt/hSqgFu1O4dH2QfyeGU55uDG+YQW92yDgN8YKntnpMgouuWq2CZg97
BEOsJvspStVJsyTSKKJ0JT4gaJTxBu0LZW8ALz5FGl9QbV9dDCFl8pW8A2MK9qCtrnXKpFi+AX2u
WXiCDPlYYXUZFeHiTiDo3syVZ70TxqCloLsMVAtOysLodPhroCF/ZZJr19GFa3Ho6hGsIoJakFmT
iMGvfd4FOubR/QTAOPCXXxHKs2+TE7TtIxTkqh03SHqctBMRdJgef8XR84wjGoigJlirwhphCDnr
od/JuTWFVzqh8d/m5x6M0DcNC9ruo6wJblZC1/g1OxyYw7Oc/vbEae9X5QQEbiXu+zTPf2AR2oQT
G/uaDFfk7uQtXyMEj987vS0G0y/nlQ23KinN+JJjgdBdxqXRc12DZgsaAvrY9b+jBAqkt8kOtBM5
G45/m9IeqmQm3Ifg+DyV9yzaVTUvRpormOMgeFGq29C2Fc6R1Cz9lujNHru51M4vIiBuqkNJ6qGb
uWL8xsIBI1xizNOyurp86weqcNYzB4sFxGFb2WJSrl4oJAzD5HjBdxylkGDuJjv6i5F1U4YChJXH
vO1e9+PJRrK3gyweyrMSYfnesDwQG5Up2JTcPC2pqtLL9q2y+QqJzR6gNpI44eYHHXByxQMfkaqc
MTmi/NU2hjMBISaR2QVMkf1U0bG3RkecumPyYhKbTfLi9YLDsBMQgVW0Ls9RMtwhpwmwO/lWlZdI
EpFDu2nKKW//1v9jnkTjIVLFUDRpW+0IJelS5H46RT/IXl/Q0WsGd0gQ4uo7rGEtwv7pA4v5I/P4
oEaMa+IY9BcCgEcD95kAdceXtRHd2Up7XIaAh5Li8XrfY8YAIs5gerc2rzuQA4JW9ohzKWLW8L2l
5C5tOhHQkgWCFMcnOat6t9wSDXI4d6H8eUsNA5MqzeEfG7LM4L5R0Az33zwbn6rMZ1zIYZx0L+E6
3FcywQOEPSbEEsFXQMzGTPAej4X8itN+XEkRrBWgf80XFlUgQWdNsoiQm9dG3YnnyNYguLWWBDaQ
kAFMXUFnkPpJufzv+ZVtNXxLXFA9A5Pu5yjm/8UbWEfwFLe4j+t7RmbxELSZHIYzAtjrE+C+atZB
N2+XpK8/K/n+kJ23si27L/LKRqROTKVkecol4F0CH4//HSSRR8SVj5m0ua9rdC7qz0PXQh2uFmiX
4RLwP2ZHFRyLax8GNoO9DsbyR1hrZ7HNsTjOTvGQVTwcZFNzArC7lvVdA1HMx2+ZzhPfoYvHncab
DkSft43JxUJy/blsmebaJEdDgUSAxeN/hDZHqztA19yyyV4HJTHAD+Ets9Jsj1E49HsAZaFt3B8v
PAkMfDW2rEcew4CmtDQ5D2inaNF7DuF8FJTDrBIWhFmaun3pg58y+wZAB3RLo56tSzjNwZT1LoDY
SiS02LOMLkGUr1pjpgjEGmN8RAYzbLFlP2qef2PW0YudLnlxN+D29pKV0TyYBxzWaU2Tu0SZMi70
D2vIRBYucvHkYQ7Bj9abur4EXvB4OJy3+dzG5N0pIIy9u6rDYD5EVP85phNBagnQ/w7qrzBnTOBD
3SSPhlQXYGo9HUkHeSaE5B38gtN5AfqTodYmPhdy6VCN+Wlc3uju//cZXhGg1vxRI7/3Ovo+BKTv
JO9UFtuv0o9XLOZtVl5Wvt/JeqgXUK6H6z/dqZcut1g/tzZapo8gZ+sL1MrznxCTt04+zKjRo79I
9M99zFJwmSf2xQ579FfhwhAYL9DYrnQb65SwKuq9KDBhHAykPI72du9rKC2gG/SDdWleCfjQIM5S
dYuo+b2jlJzrtvuMrjaw3gnotqtRroVW+++oQrHBrg8RZitfPisw7L/jv+EdoNZgVoonBXNc5hPI
0YMsrSXmzuDAW5tkb6wY0iSOlVSb4Rk3FxhjX7RpAY2RSMIcHk0lPCmb/i++nhwBuk08O3dpg5Tu
f/gGLlWD0EBCR3D3cgwbPB93CouFRJgwgb/Um2JX6GfJB94s9YwZe1CdzR7GU5kwuaLQgEThyfIT
sgZ5bE1HQL/zUb2ahOE3tm+crDAvhwB0LfXK8GU7be0HE7hOdRKVgJyKslqQIc517YeslDjxcsqT
3TwJeC0OFHN53vVN8J8Nq9+b8UDWfLDxi4bFRdUlEypqcATUfyExt8SzsmLVkOX3qFlsf4xzjFqY
aOaPanxqnKXW0fWTpqv4jiD9uj5JfA8yZBmDUvWX4BWII9d8BL2onOQZXKe97BPujY/3jRk3/3sA
SDzg5BnbVpAqljzDvnKVmCXPBDtFt1qBrskve+U6UWhAKljqbuJrO4sLLLzLfTXG/vBJ4GAeAwpU
aDKpUUS2yngJubaHqmwBr8d03/yseVaQrAD144GLHZ/e0IDDTe3rj6ISkHqRcFxaLIKhGqfrtZsM
jQ/9F/sSiSEs+slcx397RcIQRfJY2vpKRVbLdn8Ed+IL09phq94qX9ZeA4sLrYlQsBIanAEIIHfg
4hoIM4KajHL9zoDZstlJaBZNkY8mYgr47km901Xvh94Xb82zuEfJB5Uc9e6+sXRihhwHwpvyNDGx
6euKt8T/612bdcmZvEqUhRR5nNBRxzlrSvmIw242xmTQNcIvqaVrCaFO6m1m1hz43EO9n5L4JyLf
JIHrq968f8ueTCfRBNRSG1cLzt0hA2kD2VU+dsTCDr7vFScCtB0pi13oF1DXWuKHO7N6hJ0GN3WH
f73bAPs4Tg69tKk0yVkKy3WPoRVLKVKNJYKfpFH0gysuMEm53pxifbqjGaJK/V4/MhUSZMq396CJ
795E/FdHsVI3lfdBA4N3Qw/2ILiM8rZNw5CgzNH21PSyNKo1xKt6rkOZg1hxO3sf2t/0gCgn8SW5
ZBfwk0/N+6jqDBvFwmJ40S95L1wkn1JhT6Gs2eSaBtpQQpO22o+1VG3kLCgw/D+nWXSrkOTpnmk1
rVf0S3wxcattUFE02qJvO1fRRLmkASvjTsku+83VkAGz8zqhnJO4xad9oR3dySyyp80W5+62hON0
exk2j7kXFEbd2qmKjlKMD1YqYuHIfIQk7PmS/9Fi3Schb8weV1JFx72qY106lPEWazYeb0jmvqnn
dI61LpS4Fi1HmOfIw/E3Bf+aGQdo8jigj1PoD+BWzf3g44tg3y0fMwgdU5VJBsh2vucaNsQpWQ+J
50OzfXxisIOT+HSIfCFJkKuoWTbr86csuSsxpSsMryi/LEhb5m7uNJzxkrXcltybT1E29eUxVLjW
Rkkvo20qBpImrWQ9SYHuSzJ3CdKrtRgAcI4/+C+DyGSr7O6D7/aoSlkhY6lRgJ0g2sKycjJTIDC7
W4iD4oBYtd1xCrRwKSZ6BzxJM4sqj96x1nzDNoPm9Tm+5oL3cZYy5s3NkGKcsd3VrNDxMDWayhBD
7+2r6X0FllkgUMvnvEekvpMXbk5O4O0vbyNuGLr0Y3CkrOmCcUtC1DmY7vWVifEA97la2BmXyxZO
GaJlqsKa+bf5JZ9uVjX3lgRBUOkTcZ7/J4KVcLWgrimrldrNHR9k1z4FcTY9RJFqVNDZbvUjCdbK
dxm9Xu5nwsVI746nvDhWTP0k4ZfcnhV/+9+sz0t3z0oVTzemp/no8N63kn1Xl4f9gN+ycjQGPUad
nlNgUL10q4/4vBPhEvpjnSBP92+NsXs8qPuOwY/rroFayGZdDQdF/J7cY1vMIiRSTQdEv1+0StY/
YvIqW4dw6JD5xQPcPaFZjYeOoBe8k5Qv3SXrF2x/7f2PsE+I991bN7zn0v4vHCpnCMubEen70Ldv
N75Iem2FY+JULKAnJceFbV2LBNWMgyGpAbfQKgkoaGO2oIZ30BPM/RXinz+6KlRNvEBI6ZUQkdHQ
yNZMJzmB2OTfjOCPOU1VD8dfmEiYblsfEn6MlKBQ3M3epN4uTTIFfbxsSR88DNsJBS2gfHjix/Tt
XZqhtYKfGUVDapsoO0NkqFGv0qDge15hV/Ziiwxj3Jvjo6rarbEEFFkW+42Esbxw9kDBO0kNk+7f
zhdFpoQz92eJvLa24B16id+56O94Hmy4WsF/tta90AuP/BCgJaVIefNNFbcPsqNIGfpmXtnAqwkH
CSPmAalIIOjOBjwbZB3RS2fvEfed4e36BIYQi7lttECiwYd77dv2ttHDN9ztfJrBsnylZq8gMLXq
q04ig5IQY5ItAmQuaNECt5bUOqHJmk40B9KgHB5YfJ0Ba0k1AExD9mW00+yqwoApiayc11QNa6Tx
+cVp7AgW5vfGKhGKbUSKYHxzT+8YrtK4RkF+3uN0Guac7SQidGFXbe7sGpMo5jZOcmcBTt/eL3xb
7bBRoSYDaE7HbuLmZKXxj11Kv8+kaxok0FF4ZGrnBIdzzkHYqj+Wa77gYFuvECVhklwmJkkV3sQe
Nhdl0f5bhuyE+l9MEwrfCCFYyhyQX8DlztlTO7UyS9uRo8CyydWG4IJzUrn+2wm+2lGTc72ux2ju
kTb4ex2+ygqJtHdDVDp/jHDBNEbkx+UFmLmd7lSMWa0+a+UlWfdjoPqca1luccUdhFNRP/G8zbLy
DkFUco5Qn4WYbtNTPKZPcueshISAGCHU0p0uzdXGCMUNPUPI1sNdIruVOuKuxkYK6xzgnGqnXkoZ
VYNgTZydKuB0yU0iQVE1TJpavPODa6HIQQ0iyxeCJfVO8LgpaG+5MRzW5OlWwJ2b2Df2jbogXN9Z
B2r0H8HEbND14r6LuZqTklIAVdtvjjqa//fE39vJM031tAW2oosnMdabSiSViEbV23t1HrwOvQ3y
OgrBwbhnSp4Pq2Pu6uUn8mT9xE9sN1eJrruG2YoM9TiV0UBzBp9ppMszhjIJW+AeeZCyU0vrcMrp
jQopeL7uZlG7UZXyYemzBIeODiObMD8IbNXG5mKZFP4v+5mxNbrVcH9VA3q93ub8AW+scdPQKckP
WA+A0edrinyxIqJxdClL8pNsSaTHfBqqm0FhQhlfAKkxCIKSaBF7VHMhedz4sjh91jgFEOd8R7W2
MOw//OLN+/PjnUpY3Zt0lJSUJLGMaACq+6C6qgiTa3LCSqIm2QQOPmbwLUy5lMwwrYsGZgFOUCak
PqI6X8aR5vDhqoYNZNDR4yhRdpXWXe0fBceBnh7PRyxI8mmRIrxCLgV5sIi9yfzlkH2dxzimQcsG
exRyfCRmMsawaj8Q7cJiWeZmvheIWFM7gvg/sDqnM1xCn7O7/YsH+ozjd9XUuygE+CzLr0Q3uMnU
KEyFoZT9y9Hkx+BdEXFyYoKt3fieKsXbCvHfhFEMJvDVXYZlEThDSDJqorYHUeCaqriG5Dn3s9Bd
T5bYeaEsJWvo7Ua2zxvhQRhoIMysu2luRkPo8oMC0DjAGb10Y2v2vlGTFdIf6HTfO8tutrF7l22o
T6xhIrx3CT9+ZDwHMaseBRcm+JBWiRnxq5SBps7bikiNorppO9LzVUWsZoAPTMuBEEbV62KvkMsk
kzSkEVfPo33FGjedk2fsrsWYmDigbwJne+3nuHki94U0s7ls/DsUmFBA3iC+DkUj1m7Cb35fMaEt
kH2Gg8ixkTWuNYTGMuIwMuPz5XlhRdRX0U+gzcPziWXs7roqVd8ohqFy9J2+2ihZWsvPEF/Leatk
SQvemYvQUpeTuhazEGQ9gbll0JKA5QxRs4XmeRA3wpdj0SSY59PfLxFALmRdHYuBFzBNpq5PHA2G
JeJl1Da1C9s5cYlXVs3aPa6S/IIPBaO/qd3menJseL8pxjT9nzpo3qp0OKbc3U4jqei9GZjRdQAw
blKZT1v3c5vHAOIPT3VwHrPVWfdK2BwKyOI+yoChzatNZ5lbKNu7sUnSQ3uRR+1TChKu7xAkgleL
exsuQjXMQ5NTcS1N0IOPME46IutV4KuVwBWZUpBTKmlRkeR6vJD2xBj7SkbESzB/CSdIPk0N8Lml
AcKXx737Zz76ggTexLo0AdbBVLPSThYIhQD6OfR90ZuwJra1GgRvvGkP46hELfIyhA5ZuTb19ypg
8ZlAipPxzrEs5Av63Epm8kBajGODCT75V6gw7SWquZ6y4xjGpe0o/38qI4yyH7I4lSJti6PLX+mZ
JvCJNZyfBqkyPfPU6fz11NHuekeBmjXF6dXh3FKFB2UKUsln4114ZCpVt0gptP7ZkTUhy2dWslCW
ObX1c7c+rjqA91tFi8X/Pwps/FpFx4XV2GkWL+gjeaR1dIwTlyQt0YIl+xs+5W/DZ8J6FjvNhOR4
JYMxkZvcp7BlQeLf89yBIcRzZmzxCDiahDRGpjbgXRrspUOezAaffOMrI9xfNFbc/yskdDciM3jg
5YT5utmuVySh3Uz8R7hN/ZXDdUlnr78AOWxF+KIAdT6jevP8qVKdLXSxw/ZlrzcScvb8uEjBe4Io
M8jxBx94tPUUS0x5mpjVJjIq+pO3UlzXJA8KKEOQL5SbnNmDjn+2P/ldg1D8a2xjmldEGyu7TFPa
+ZnCiAscVHDokZNEIL+5lV+Ex0abqDzH9ueUS3Wm2A7OaJwU2QrAHqxxV6ZISJW8orVSbNEtznTj
wIiRg87/22czsw+/1ZGH7ZGjKoBDSl9xjs6VJ2yUA7Mua+2MHFYMiRjexZ9b/AHZJD8aC8P+lZlh
J9TsCppt49unIrPLzJIAq+lIg2uAVJT+AIBUNEMTWTQuUKotBLoUAN2R3ZGxGbK2Bigz/9CJByom
inioNLfk4ZURC+nQ5MAao43hwps/qJr8xNK+fSe5qHzNsNjR3lwbPGrBOsRjG8Zzfo1FEUwN5BhK
5TxkuAPqDgzApVgnlk5fBHWcsDZ7zyP8rcUNQa+g6MCWChQp4vy8JOxj1FiSbOJa7iBCqHD/RWBd
AJKUJPjt14GXrum7pCtHc1w7bIICs2BBMaz4c4YG4B3a0roxFZuZiTLYe6MvurSyI9GBGI/xT5Fq
fM/jxPpW8G/+g4txAxSMELekIzrYiQV+P0VDlTLZoVdt3TLHnB6u64sq9zzNyvCSwzZqpinuafu1
a1gaaF9sLUrJWlvJ+xN394P0UplhtibT74NIcRq0XUBx503b7N/HvVWhV6wZHXDiqKyB3KXOeoXK
RZGwvoN7X983L5p00uvExvL5/l/5Y9l4kAvPtan3WsGcZ4ReJQbcS/O4p0wTHmhBpsjzZTyVSKWN
/x42+hdYkVxsC4s9uqZm6mzbJJbNkQINf5i+gH7yZK/bBoBc6Q/+3SXqHKviPw6UO15a6bqrciO/
vaZIbJeRhI49Ti1Rj3JmELB0OHb9Gq0liY5Dhss50Un30ajtreg03Iu6eeIUj5P0EVWE9T1WRQxc
LbhQzsM8xH0TI6qmeuWQpHAUam8q01lF7YKl4XKPIAiVxOVFPlgVpicC4RDINp1u2dIDKuRFR2O2
7dcC5Ka6pqZEOsYU1Eg5E8VTTX94xHvTCH8esCAHCs9Pf0C2lnVeNFySwxefDNhR75qMYe9dZkAO
rmMrS3bhZWrOBpuRrOvHJ6niJjTaB30WmP9L6UV1xALGy7BzqjpikA4JBUhbSGRdR0OgWn7p0jbt
QluWC9SPFzhB7XJLaCe/Gw+WyrZGanGj+nqIw9raSKEgkQRRiYDpMds+y5TSoy7UI9+LLKFx5xIv
b/Glwuz/gB8WAU/dqVfV/Y05RDG3zE8E62zIcNhzcEmFzYIEtHtSOt42J5/pvJk9ByZtarS7bMM4
ITQUN64OYTLik62F6Og6077KloCMXeVw4KxAKJyF5axzvflFTHCOMJDIL9i85qe2awGmJ7JonoFb
aDRBOnnALEBYmqMdDJmb6CUMQ1gLtQCZb6bCdd/m1jyvPWDyaZCSHrdID5xY4cA9ZecKJs4PzhOH
dlNY7aGtGzEN0Vyg6Cfq36FgjYM9KSf++hNv/6NTvNSqxwMeZYUN02QQEwG+nAEYkpLXJQvgTaOD
KU3U2Q33Dn0CfMWE+LNViwGQDmaVDn1zUCR/0UysOJrv1iZo0PrZkViS8Lp9cHBLFr69snJFk4Ru
4GeEA15Q0uDLU9U1RlzC6BUMqVa7qIHz+g0Y8hNyEI9gPEIFdSZ2h+R+pIaK0whVl75RWjXg5h65
y8jqYu3hxj7SvhQJ2G3IJkEh3M4+jHJjbFN1zH321aAdjlkJC8Hv63FXVgAo7rk+IHk0qvsTNnFv
YNjNfoWCHFpWP2aX5TuJxwTxnlJpIgys88ZVtLFJ/Mal4FGvz9AXzEcTzq0dGoVEInVZ18QRrTye
TaSH3qBq7xuH4yo04PUcbSB8kXJj3+rdoMkHOh/Q68pEoSxF/q0/+u5LJdjsU5ZFh9BIn0iGGShB
olG+bc7ymDsXown8RINaDBDqOSqbb6ArUt6jOpylPkTJhCrcuRteY2MA5Q0tZn5TIKu67KOzb1GG
NmFoPVKuL+2BE2Y6gvvd9d8HAjHVU7vOcwG7GxJeb149lQknuG0ow11Ymcjfrd5PlPoeUUyyVRhS
9FpczlLuft/iLIH9/92TsYncZeQ6pO5troCA5ZvGQw+NVaYa47GSpET4QPPUB+Qyir6UrDN18/br
I+39nzwEUvONAxz5WrX0uH2KdxVtH8FlN7xkPRuqJ1QmUYHj1BtqYBkzHZ82PHYMFme7qRzaTd/h
NsvYeneYt/4DrxodmRUVe0NSM5CNfwrUMdZXSvJI8iRhuUC5QBmgG9Y0vquOpGFoF5IPgiTvJKj+
D3MCN6ulN7Y2O6gXdOZ/dqpOjCKYMJjOgt+oY8CAsBAtXbW4Gw+FPGBXdPakULx7ROFLl1AinJcl
yTrYo2UPRjKa9zjJk7NRJiTg1WzfpFcAsEp8oZLxlLXWOfKRF9YM4V+SmpM3dj7q8GVLymzkRfLl
tlaRP5aGbdS9UPBtdMQw/cnJfIfnS6aU5YAmp7KjssGHV2XdSyt0kxyOCbYC77egRDXUlDkbwcLP
NLLpw7zvUEPcyF09FEABo9/Tu2eaXLq2Ax0T54vfjtgdmDwZga1NUO+ZcsICCQwizylaVdltA+B+
dkS2fizXo+rW+vOFjJFQa8UfwSM8HMcQBWIZMmp8zLBsS3UCY8+vEoOVWwqnWLTQsNpnLLyMHF8Z
7hYJHGD/wUT9jQsLuHKT9ZFQjkoeVNPElUfgu/qtRaUYcPwUMiayj5ZzvMc3Ey6q/oIEDHCI56fX
h7F8u/qyLQ/wzU8qYlYC9Avk/VcoBJHfRL+VLnZfB2Zqrw/ywb/GWmyXOzoAiFLa694AssAxrDJK
WdM2ODr5XeWG0VuowLJk6VGSg6Cx+BMfO9gtn5DXSf4VhlFnHz3W6+9WHnIOK595or+kvAQ22UNf
srknZZf+yb5Fplzy/f2dI40pZmltNBr9395POP4kOAhPva51xYRN1xP7Cvrms69SDglkxeGUqKpd
pDqUS6euyIe/t0D238iEO8zLzXkZSrly5uVNfw4OyKmv+FoH/mMink5+zoX4r+ix2+WOdSHUBJkA
0O0q3d9ojLfZIa8z5OOtLxrtPqjsNO0YiNGqexXjhA0BvYg1Dukir5riDM6kV8EjAe9hpFwnZK0P
itX3job7Jn2eeTlhT/Cxc3tSX44nd8dhOuhTcWHtIx3/0I1GLtsTk0nqgctkFnIRGgbAeeUL5G71
osT2rX/T/rC0sv23DE6PWx53nEko97XQAgXbxIFpTzdHILsXu4ja2Pw+5SkcmtDx837EhdPLRpTt
7wNAPF4W4tbLhEVNH6hpgUWSqkvRkUgjsNrqlyCgni4Mv2Vd4pubrMpoHmes9o5e1+YpMgOu3ClN
EttTz2nPB5NpUMf8GGTpX3M/1nOSkyTSt7klBl6zkrXjP7gd/Bwd2p5IPF043/mIjmgZOltL7o7V
EzgLvR0IOxkMm6wHbLlys7M3+KdKBRilHV11QSAq7qYVPEAWU/DCyPN/Cr6eT/JQMbGxMNx0DoML
jjrq+9c/X9anppU4/8yNu+rOfIoutNvY3Hbx8THYqEN8viDiRaRkf6L07wtgK9XZlHlW0yXTKOII
FTvjL2vKdQ3t8C/Qy4o4ZT0XKehgt4pxLZdYLz4Hav3lpSKLUR03y9jEyWI5QJKvoDomlhlEMYt7
xp2qQCBSvVFYmBgbYOSv/hNFBiYpUl+ZU6FXhN6N5tW1SsiA3kOkl5KmhCoA/ZjMceuLbJqlnszt
Or+aJyJcvNKD1jbHSnS067dBxlnGVZfZb12+qcFxxt7pkM3jceQTd8O7p2q+xTsm7P7QVYevTpnT
l1D/j1Ktv8xd1ogcdQtWlRo9I3smvB15OhNyAmsVyiDzQWZUl46tG0pnlz3T27L7MZmnOUWf8V2f
+y734JAK//WYXC+Bk5RvDTOzd6regEbOw0zEO0MVmfyARc7OJVt3v2sop+v7c7RHegmsP398qv8t
vqJNH+4JNr0PiYaupTlEqgXfMM81mutAYgssXrx+1ozcNYzenVxqjxIupWPeZUVzwErnV0WgsmjP
0icY8OQ6KrSPvVSOytDljwDvbCL/81g/kNFqYnH3+x7PGveJ4nbe7dcXvVOu8jXciOd7UjObUY6N
92GeLbjkZm+MKGdkBCaOT4C0C7keXSzUzQyZ2fy2Xk1nyUAacbnBrwy2McmHj4bfcyajG6H151U5
nt13morAC6uiSPKW3KRT/o1+fQOxkPATHqvDRCLjVEWa5PCRLNvinZMXY/Z/9y324U/0Q9v63Bw0
HO+3EIGS813iiVw+vI+bhzdVq8VRyjX2gm6rWPSQACD++ApPkjwArFo4/3UMq0olz+cW0YoSEOHC
L9eh9KrC1QO91+eB3qQ+Ub+d496Vzv9iEVMPfme+dPSlXmY40M0PTA5BoDOnsBsxctFScOB41Gk9
iap+yLV59LyjDEv6EUiDWqvoHqp/DTQZkCyQMpGQxm4QrppKzSRIGRrsSCTZ4Yw82m+jJPIZDtpQ
YIMAdg9K1cmKWiVIjhLcXCGjl0ucQOCRiiBAHDiZiQq31RZUP7+vyuCA1SLje5ZCrvISouq8wEIc
PjlmhsRI6oHXQSc5HG8ydYfxZrmZpIYkMkIsSX5CQHHwEdbT/l5UpiMZNwTfS4ZqiG8vVOh2U/Py
2O8iTbZED6HXqiUwts0T+ufWdy8voZr6pw7sfKT/0dbKVQ0BbISPbC4VweslAheiexuFn1At6pbU
o1K4R9H2o+0/UmatR6SLtVypinfX0hoZK2nn0Frae62obIPZqJgYmtr5PrULBKpClhzf9SOxrnsI
c3/A+LoDs73a9NjfoplxRHxVpyHCfTFOe3GS+Q36RrWY4zznQRZgZyvYmJeKpC5icW1oW6GBg9Kc
j/1B0nxA6Rso5zsuFME4uhJRZfL2WeJx/sF6yXzcNY8wzbCnyXUWr1cIU6iUFuSGRBNwuXUzH3YW
ZDUoYGc1aQfVhcy3A5+y5xE3Sa5KwKyIK3wt+DRLx7FOlJBuoatFCRUrBXEcd2f9TzacqgU6qBPB
giCVp3cHfFTOkAQOTdbgBxl+KTKjkQyC6mbxk2kyh3PvlNps6kOfsfEWvwwYUT6v1gftUgtzkfyW
5Si9aGzlAt4AS2m5c0rVsYi7w7kbwgWXnTpv8hB86lsY+9DKk204AeLfTKwOzLVi4tlMxPqPknVE
9RvD84TScBMrdEq6BzB25cbtWy+5IZ4bjYl8riKgxOzpuzrNuJ4GcQ21s0p4N7T4JD1DiUkna+vf
TPxo4XH5MGbtR3R1+PJmbU1f5AoQsKz9Rm4QCt8OLQo8rqN1N7kcPWhK16OjcA+sRNhZoQ3M86Kd
ZDUlUdYMIE3U3lzNxjLlRKllJ67qaO3BIlWMtWtOLidWqj6ZN4m8HwI8dj8GjimP3yXRIRGn3RrW
0ANh1oThsYNG9VjqM3QUnuF+0Dr7WBfX352v39AWaTqyglTWnQWqEaSXClbEWLKtbylpt/qg9SI+
NztM1cH7V9qUeK6yD9t1qBBNbl6PyQkX4tmFMIjBGe37JOYOaL0O4pcF+PRnMuuCPJUweJDO8TX7
Vypf7xx0LorXtfxVc1oTKNZg3uD2NuiZacC4Tq5hjjT+md2W9CRcdaVS/1umHHLPpf2aojApJPhB
tr4E9NIiI4QZxYVz/4YlArNABiU/d36H95sUPkTCx3j20oUukVSy/ZFOg7I2V9Ye615clll8uB17
UOsqaHwbpn74vdpa9X2W5d0cbATx0MyrEE6QSOlasxR5V4+7mkiyu4lgJ1Rhv9cx+MdinbEMnZ7N
Nu9yBzwdOYt5MlUY/878tJq3BdyTYsnYDnnvIo9jvnZXAUEVvqbUaXHQFUJhOh0zYwx/U/EIVS1K
sXNfEF/p9RRUFkPGyvPdej4lxz9EwR2QpQ1sBrPqljTijOZrUGZLxyar42qbW0lm46GspL9U3uTI
LWNdoKxFOdALQndGFmf7RpznkGAhJ3xbp7+EV70naswi/6DeRC9g6QsSqGhLfB1RW7L3jK+jEW83
a3B/WNdmZyYIE9A1TFIY3AHZScDBKwzXvrrQPsKOQrLgtKxVJ7iggO57v9nYtVVFSW/FB3DBd9h9
WtT3KHa3Qdsm3IS3p0OYnenh8AdYL514R5XAu3ct8+IbO8AzHcLTjC2cGOiNI2+0PrPeaTNZZDsk
SW6nKEaOGCxYa0gcSF4D8ejSOaTJvGuwirAnoJYJWONjMXjg0zjmKd9YkQW2ka9EGWUDezCVsXGc
jQn1dGUA7O68RY73iPBFhDC52MQvYhNnY0k74R5EMxAkvSIhoE9K9uEAwm4diObSMOjccuSz63Cq
fsODRALkw2wz7WcrtGQQzyDnMbx0cHF3IQpCdBarV8aIsFqyHXNNSENyEV5FBITe9ZxzmTxJm+48
NyiB2D2NIKA6Z2ySBwjNx0qSVwukR5Gua791WN0F1nWFWbzxrxHNX29j2hVgKQgsnTmTd0ss1rM4
V6Ov0zg4ijsVEo0AefoUzWfCFyNpdngs1FYMr40Gwdk33cDkjb8pdMSmYGtv5k1W/t0WjdLnv+1U
fGtTRzPW/+w4/CGnvxRa6ZOVh3h5TMHGyZX8gdxQMwX/+WptNSSQFpxUNMkA2JFttXvjutAubXoP
uZSM4Ojt1H8DM8gtOjPu6sJJ3d7PClg3DLU5ocDdJfNPoJM7/lL6LRf1R861Y3gk91dlG9+5M6o7
/+rnAyH9IbOMi7nuMfTGkf2CAWgOpBMTpF2tlgQJJzf5815e+Hsvm7mIt96Hs0Cwhym1K9W+QcW8
JPT7z+ho5M7k2oZYb/h2PO16cx0wtbS64GLFW6QWp2+gT84075flb3VcIbgvjCldJVdiFCBX7D7I
xNui3Bfv9CzP6vfvLfsCFRSOBgX85jFSOR9q0C37LSeUezrTh9JUgZME076TFJvCoD9/bXObObyi
NWD+b//0cBUIMndDl+ylCe9qtOCWbAZm9efhkeMNChL68zCY+MNcbedaTBuozM+JunJ0+Hsc+NNs
NSIIDyatjeGOVbOFi0wiWlMY2Rj/V2PVifl+8GDrW8KSUV3chctTIhrUkND39PpMGRrinfr+11+Q
cMLuIz7NCzMxz/BxgDVmjp/87f0iITnjDZ27sEjwuy882Y7hJH79qaDrQereXMtvRTuL5veGwpwj
ITjrumZizzv/tqQoa2k1Hd46XN9lr/N++SSddlEEjX9IBCK5nwiSmzavI8LXsSTJVow7M5Qwp90I
DCMnQNgjX/5Rh7KlP6olvVoCoiwxNpJUE6FS/xkhHsNBXTExhTnaLYDcou8fV/gDVxhQPNgZTk5B
s8Neyr2P5JchSp/7q8xA060YPXKX345mj2FelvdBrrqIA1PQ8NwFzkcof8MY0Q0AxO8rdlKlwBIH
TBSqYFC2G3ZJ01Ng3msSTOCo1dfvPph6dNaaa3rB5dszxHRJk21YpfO0GjPCkxUN0ArXdacfv2qR
eEEcD782bFpZDFrch5W1snyPNUXomrebrYBHV0+oYlx5y1R38u0oicTXNUEW4ciZTY+RKe3B+0Yl
suSriZXGjrStbT1QKz42cjhbS3FH9YzhsGvY8QcfVvzkVTreeBFIaoHquZ6sL4HOhGsEyqW/gg5H
GXczi2lpjhR+H5R0zssb3Yen9C42BWGBNcVsh5pMrk5nVhhbVstgvL2fL77Ky4mJkn4SBAkM8nAs
RSCQ6NmeVxJgxu7qL/vhPqUP65XYqI7KcmdYrsOK35JPREHWpU1RIKwtwcdhxtiiA7XagMaeFTzD
MS5V0zMtLwQsT/LIkrcylmo03m7JzhzZyR1OxBm+ipdOigIQpZ9rXPMzmqRzmefImZSokZ1SBev3
b5HQ4ESd13NZx+7s/Ko/KKq2eEIILaBhFdVlbsEpqgDojBkYavey6nrovNdzAN1R6h/7YJ0RnAY4
e54eqwQSr4LhvfqWwXDV+XCLoh49wYUniOVQy+qnFscrm/vM8kO/fdGjRkvRJqnL3bN1UxmmW6Zt
t3wMHUj2VWPUxpjXCguVA/wcanQkXc9psbiVQOtLRhyjTYS3Lo1eugdyIOpbxTXWy/5OXGhMAKRd
PI1BMuRZ3DS+J7NNE2LKF4bfh5V1/LapJkuxSov/g0lWA5gWXA21/PgOPJoaKHGra02Iu9GlzuxS
bNiGFWkEf7ApLdCy3kqwIMFNxJVLy4JpUQcztt9akntsCvd3gP6M6vG6MupiEM1n8pYGua2AATSo
1q++KvKNRKL9YyZeDNLVaJlrv3t4PlwbmEFdBdEncB7F8cXhZ5POQlp8d5IR6d0a5MKXdYeWafh6
SQFJvey9z4C53pf18lPCagdlQwxvETwEZ1bxUHliF/3hpkHjMWCNEjJzZa6w0fnoc1eMKrY8lVQs
9N9DEJHYabi6ET/YVN/TTGIStwVcVpW+lkpcanbouH0BDieXREEpj1Kl1ubyrCcwZsGmusjBiw1A
7l0jBeXIoOi24smQipWGzOn0GezSTgi+nYjMVCYpVbYNn6A5PSo6QzrDJMyMkG32l9AnGKIcQzNU
ON7Wi049wqZtCdJsbW4D9wrlISf5nMgY3VKNldi06IgUmM5dvjnSwnQIPps3fj1lrFM0ryvY3Cmz
1HwUpl/JJl9IBfnRDF9M0bFbNeFr4nuUeywF+OlXHHMuXSaHKx4IQFDIINRBFy2IbZ+Y/GvUXizJ
TFCZ/wl+KKWVD2y5Y2vE48Im0re/xtuIK4gh0x4IY+DRlaWQSEpFYBWm1YHjS8czD3thQ29TM+/c
SVAD01DZjDqpT6hue4xNU0Y8FpbVIoo2U0fXo6Tb6fXOuYjVfTWNkO0mi6nJQO6w8D5XGDgYfBj+
wXBQmNGtcSoRvuulzNAOmUKnltM1x3FmnpCFs9H1DW/0NGmXbokZNflzKcuSy9ES8hUp6dGTFXNw
F9inf9n/4xHclnp6m5TqomX4I1vEsFyhWoVvCJOPoy0XYrCZeSnbJVhoYGC466eEQaPi1zT/C9rR
E3PvdDYlM4M/ypxFeVThdjra3ypBylaoiqIET5S5mwE+bJMNd9eawZ3Kc9iF6R/sV9NlCH+vumlO
hDou76KIe1WIGsHf+qnQ+lcmW1IDqI2PufimiREVMpqSK31YEPV66YEHbxfN4NJid6D9wmxYVN9J
xe7kMwa49yjhOJcizjXw8uPOrCEnvY0rgalq04SUE4qp5ksGM6GE8nOVsi4QurN6U48kS//VUkEU
BbgB2r04Zi+McTs48JoNNLr8YDYem0HTd/yDO/EfulvNPR+SpR8iIOA175rnuSOj9A/KwdFhEfv4
BQhPhKGXEnp0jHJqG86Jc0DxVLf6oCxSYNQDwVsgXw3X4J5RJLPM8YNK2Pi4LQhRwDnwFa9Ek4+/
d0LEWzBbj2lDuNeqXbKosduUMvfkjbdOfQMymV3YdeIMU4LXGQ7j57YW1665ZlF6nydWrVQk8C4+
leuguR1uxXpvKVeCtMpID64Rc4QTh+oDYl5BKW90m2dPPnv+jdI8sqe5M1+cyPt6mx3L4Z83giJZ
13Y4qiKsg6kJHasx/h8MtidazOF8OP8M0fwH/wIQehzaB4TyZj/MJVHllklhaFM4Se3htD34R9X5
aLte/+YN+XgoJtJRu6wr41k679a/AZysACc7u4fRLuAysZ4U7cLDUC1l0At3rrIuggf4rXU61Ica
s9N39Aw4e1Vlws4yXXNORKDkIdcqapLniEDVdJMIvVmsUD6f60CbpkyQo221cx1RedQ7noUVXfGt
/TSzW4/fRGeUcBel7weGsUQvNUwikOTymunb3Bja8BIz1x1IdDooeoCcbszGonf7u32PRxYHIASt
6Xmowr0eXN4VrAlYi84GAuK3gpWAIGChHZEw/v9Q0WNurEY8HX8SBjo25s+RkbhtHrGsu99tNuK3
7lP8i3Mn4EzcaVuUh+Xi7CK8P9QwP6cVax5TdJyesFV8xkE+f7F76SDr5ghYgkpD1sNH7CVrJJ2f
/ndR86btkClXvCp8ovscSImv7xewrUutXkL2FXt6l+MMojlgKwDBHqJqNYGPzLfvo7gnCR7HhLmT
bbok5H2TW9kiNM9mQAVCjQAyXfQegE4FfR790ebTLys6OFHRlTTNN5AlqC0lB83jZ1B//5zXPl3O
ofscz3o/KoUXSJM/yVt3IpCF7nYt+TxLLqklsQ8u+QCXK4/FHg7ZyGa551Yfj9FJzmrI/gHYbGIZ
+7P+k3dTRzizKimiUK6ZtSuBdBHEPVDVKhlw8z9ADWC9095c028G4FtDvBbRGe5ii8kxQ5HT/hi7
jI7NE8rscVFSfbOsGsBOeCSGBHeklaN9O9QEMcmJdN8aA+mXWMPOnSNFj4wSUF0tR7BIaLDNbltp
8GXAP2azLxQVOwPu1wkOe1APFJCarclSUFm8nBY4TrFQRWwUXMt0GSVqJcE4f3H4Ib583IOF8WCj
5UIM4fu9Xxv1mfqCi5scwWqaTnOZqR2lMVOa6YLsR+vYXUMrT0Amwv7IkW/TzS/f+/sEjAKxvzV2
PNfpF7GUCoBdkd7DsVohkJnR8aDCNYoGLnzEc5PFybwkCJGpYznMoyAEsni44egWbsvwLE0PGyTd
qahlahqR0IMmJdTvHuuwF+Q0aXur2mMq8HjxsCCc9Dk4ayaWolWPoU7u3Z+z87m0hyeoKwMZP/LI
RZafSJsz2C9NG/x5UVQFgpNwtcrRqf9r+omFN5kr/JPSHlJwVZoGqKeiPFmziRcgwMP3MVtJjkC+
4GxzVIxsDKrkpte5KKvsBif9/aCCK7yV58RUGIggJvdTAHwIgDDXCUlnkT4/E0yaQsJ2G6f3O4Bj
s93PKUf030YsaH+4SBLs6JltmCHcioAobmyKMr5mZRn62qfV99Ec0Yex/JY5tKeyhhhlXDrBWMTo
nO/9BCH2Hx702KT5E0FNobVsRWO67OjlbQCH+ViDhaAqJwGnveNGAhi7dw9aW33luNJdMktFLP+D
9nTpi90Q+DSo16STEPCjJrzoyb3CJK5VE5O9kDWOtHiWnpbT41vutUwh+DbFzE+/8ga7PQ3liWy/
ROtsDKW7vO/StxSTzh4JtaBbb5PHjdvwWaLHVnm/2Fz1o7bNRE3uIHeOanjAxdSfhDmSTfnzZrCu
L5yT1Rj+7fByMD+PNsP5jXxprbx/F/U43WwFIFnQ3La+DcRT/JCi41P0KW/wjnRaIQ7wHmJ6CMrN
q4QbX83fEXnuFeMupo+yHTJVL0AI8VtMUA/Binr2XghCQ/haB3jcjYpt83CFX1l1X/nilWTzcagu
VOfTP6d3p6LJxOTM5gcyQGSaj7DNVG0R8qVC1WbWgywugPxpO6uugOlMNjSmOFDE9mlfQwICkWbt
stozjwsvWeLnxoINHBvrQT8/4MhbxPumYVbi7ozTYkmH+rBcecKclVxnguX07xh4PY3B4SyrTtoI
mwafoREQJZsvxSf0ebclenrTID9UIp2Ej+s4j4wySks8grdqaWVjFtipH3i2HUUXJRAUtz3Mk7zt
osbW3YViMhx3TVAzTVk0qAcuOB9CzRfwPQWP0g4KJwAaskH7hwgyada8sW8YfZIuOtKfbHgUYtn+
2hQkYlGirPdxR3VOHsH+FyZ2PNssf5nwOftpgZ1qiuQU9G4TNSj0qusWiBHOfPEPgrQcBYrVsfrK
XaGqSF3gYBAMvnd3KCq5+tVtKBFThc3VmhBuTEUJIXP41QbQ/k6HnxlTb9jR0nM/TulfJNkP+LzX
swQgu92CIGS5E3ixZRXfSxDSlQ7dI1TBCGFnu6nd1lRxiGFapRESdw8qpLZyiOw7ISXwWuXBEQ9o
e8SKXORk2Q6jHqFGmN7bstZ771Jha2nS46t80EdImD7YypAUZoQnGjQfR4ICVWbhhTw+HPCaY8br
YLyQvIk0KW7wg0OTSKwcJufin97A6ICxe2QIMrCUf/EvKeeV7z7ySWEX/FdhusbySQnfOACOjCFc
FBHZ+NkW8omkOeTx/t6ULxnAytXHbWhJJChz0I4XbzP+q5pNKVPdvV5MXJ/qlOosWKUeaZgr52Wv
p8fDuvFBXU++G9EFc5+NMeECPd30UJRLQRCQ2jmz3yBw3U4qDBvPtaeE0xExhAafGRGd+dykgtmi
BL0K96KG9ewroeVqMp0Jh0PVZ2jwBSkqWxMBPGjFocauh9DXM6v3goqrUICWtANMSbvV96jN17rt
Jrs3VwUcUT23bhUTLAhEOR0z3iziKHTgnkFk2y59+GGfad7ZBtparobYocDDz+AbgyI2kopCRDYa
cHNAqAGX6TWlUu3Oq/7UyLA6xWsNj6Ep+6xi7WvqyB5X6j9XBrT9zDumHaKNx9SMZekcmZdCmvkN
R5a7Q86dEuwpduf74TTHpbMvtVOHa27xqG0KxJGCktLBFf0C6xgHA3FIh6RK+sB6KnIkI969ybVu
BEGwXiCSiDVUTwWuTMIGrUDiecnutUjDYEibqS1ddd85nTRzZRpzgkWJbZk7zXtZ1pvWSjLqpZV6
vYQ1G8vkzdRd5arkVc/rHtxLjZr5X+Jy0P7Euqd18c1rDH1TTBUouedZdSku3foLXPmZPHYyXDa4
Lf4sfDIAOSYdS3BrBN+KlWVVrL6ur6RCo5NAvasjPUtVyLNGrS2nqGisQk7Qjw3atBFS6KrUbM3g
tpJ0CEo4bD/XFCD9S4+6wXCEEAiddnniqbNSgWivGEPBPPaONTJW7YwOLOUw/daL7uryIqVfKR9X
1qVUw/whtmHyTAA4qqwoGkOnljgtrs8ZF8UAFpvuR6AaGxqJHdR4iRBxRmPIEVCqIjtaZGsVd7xx
rQFcNwgx925wZls6ydkN9AlNZDaL2T01UZguoVt/Enz3Hlqe01q8+EJ43M+L4gHZpAs+hDW5MD3y
q2nZc6gIM3g12IGQgiZpnMZxs0aPaFrbfFdrPcMEBz8eeFgTwuu97KTN0tAEfRJYqFw1KFS3p9tO
jZae9OHXIgJtJ1ixsC/Q3RHOdAIebc2spNn65GpY4d0xrUeMEtDSmAS49kZiIpry5b9hRw4Rv25m
VNLzUO29LwWC0mrcmOndeYLFNlxQjdiT7mD8X/XbDQuS5HrIKNtmr1o36uc9j9eSC54dMvmwekWD
NjjKZ4y1jvybidsmAhLthlOfAYkxs8a5pUP11yE3DPsoDS/+Pc2aIHiaBO4FACkVC20tWTeah5PK
OobQrFfrrgNdApwNG4YEE8L88W1RxmDE+j2x/RtoSr9QbXgCcu1zSPyBSbx65eMRmpluGL9VBvh0
+eE81RfvFWT+cBOygW5bJPGJd2MfPxu7gvawR+shyv47ey7NvSG5uGI1DU4u26/n9QsWefLHbrxN
BtOxDhTh8l/VFO8tncc/519OJZZP0s86BJOoZACHddT19GIxXB4zjS1TI6A+gUHXob+UiVEQqUvW
zltpbmuP7ViUl7HGxyADRsdcWk8uoCHRNc81DCaYf5IOjRnh7CcHgqgeoMKeY2UniKUOUz2g4+ks
rEaHLCiuPvR2jlbkDuGFKYT0OpeuguXzLe3t15PgFH8IresDi5GgkZezRnqeMnfjTlrAyFwY3Kf7
UKmndz0+uDiZthemN9bVGjYoctgmoimymO1ZKJejXUoLNZkzdjZ5cdkXSCru9HS/AElOOUS1hKb2
Bh7+Ci0Q9ZuSlwVzB2loo5s8aDfdgYKjtrJHaP2K+0s98S5ftXgUqet/0rKaGYc0AGjDubSDSVvp
oxWQLReasuX9asvHOuuHPnkC4FkcEr4+gXHiraLDtIziq0ktQIwS5s46uYikCkYs1BvRnzOf+OrC
ViYQVDW7GebhnxeU0pbVBcdXqBVQ2eTkgo79rK/WeGL43Mkvpd1Xu2maviYE+i+ycGSbEiHH3URL
NmW/piZGSFRzVNkeY4JVqnuxsE49I7QUL08r3VSjQwoSB4rdE6wjtJpkGl8sUK9B+9nWdnu9KPCz
9LcMGMORTJE/kZPMgIRzSMg/vcO2WHt8x3CdtAkYx0m7N5AXPaw5cVHTMWTUq9SZulQ9gvD0480L
xtM0FdCk2DkMiedbdXs8BoWIS9DaWIITratzIpdI3zYRsScVgs+qyeVRXE6tyYArXsvbdLAmbDXu
wEI0RDQYKVVwYdpFMmoB//ECRyp32rVF25egV+EpRCE1s8leUE5FFLTId32H8eGUNs0cCpj9hHuc
Ae11BB64uu2ol+FHaW/I3GG2elDLG5JkQvCMeoq3obDbWLrCZQqfo93b+i1IaQp4Tosv6yq6ttmW
BGuByl+b9X1FZjoCFJC737arHdqF8OxyccfoostrhxiPAhKb1K7PU7rqpdQjeQk1G126D73AgHk9
VMJmL155Jcp2dFTxQIAcuIq8Pcpa3hVTxL1EgGCvSIZWCoLs4/Wb+YFUejrDNaCq7xf/doQz0AcS
iobh055quQkxx1rLc+b8uPKLzcmo5Nlayug57XlcXeSBOxJDefFTR1I51ptb/IPkPeoiT2+mva1r
I7rih5odyYqr27Ci337sMT7Bs+lN5vDfEA+Nd37Y1fLxc5TwREwc5NrtiVII8H6wHlwlzT6uiscE
70WA+zUrg3fUFp/L060iTp/igDact0JhjhbD5m8QJXzz/rBi6ahtSqI+Ipid45Pd4+AY4e/73iXw
jIs873rgCqeR9ju0WeI8yvNe9KQInhLykGHPvZ37MZC+zhUlqo1YPW3ogTHwEHtjGRfikeXovS7b
GhUt4ZCKlwGbYVJHbCGfm+FnVMRnyenx2sFYyfeayl77VCw8uugWkt4xut8yBaD41wYlSKI9rCsA
pddVbYL70+r4D/lKv8OPaT05g2eWKZ2/1Xz7G5QSQS/kghRWBOHKZup+OjOTHpkRkpjzT4YB1QUV
kfqao9i4nrcmtdMkrT+qETKodRjlO4DMDuF72RicvUXQOBUGXIJ9Wk7XZFVV+4bO7QXoY5hOfFVq
BG08MLMxsjIm/ix6mMmmvkVq8ACc4rNdPkJHrTaHv00mYI2y/TQCGptlw9cUXlTU4SWt/5gHTLds
BwIo08kniFURixJ5PJ6nTHwy2s+jBBueX+NsQ9JM5eZNlClMaxegJcwK4D8PuARrUFsJxGU3uYik
/bdnMcdPVDY8iPls8kCI296nW9tOWub8JncVI/pMOnLUE+h3V15k6eZ0x9sQrnT1F4/AbkXYXcGZ
UnJLhTKCq3ZBtxKyO0bCc3xowsRUXzLZ6mT6RHwtj9ReEo2v+eo78w/lY7GUY2rxAMyh+4PsKDxW
iS9tyl9kAvpCeJXPzOYxKBbB4F4aqj0+C0kGh9CLKkEO90eg0fOIcWrRouZEItlmKIXExru1OW+F
ckhZXyTcqsM4Qq2RupkbreME1gdJCrJj2hc/JcuFU0LLQMNkF/bM1TEEVniv2mcmXYBjaRkjt83B
60urgXjiumwc9/rd8oXrVunQT5LLH56ptKEWeN9oDhtVh6lL90GxUThpkRLqWXIEhBovArwfn3lh
iF04VlpHgnqK4B+88vLOJRKzxE3vnLMNIh5YRmDZiQUCbZdT7ZfpkS9u1x/iKITBOop2fuOLYL4P
7ezrXhJGV2QIFnTf7TvkRKydvfKaP/dWA3ycb/UQNaQuJA/rQebrEsbqBNsAnCoHbmN41CPpSlQY
kMDDhpP8RBXyHaqjFSBzraboqSG2ymm3sstiUcElOUfwElgzmSriMdZ3Qd9g52TwPGwIgwNekGR3
zXPAMvYHRaHIZxAQAbDNuMGsa9JPYyOwzrjIcUsduULv43bCmd8+758KsTjKym3joRYayDU/hqMh
kUQCfrwdkyPMgLoI7I1HCs9DKhERybdkVMBC6794LtQ68CH8IJUz6NxMNodPcSbDzzvjrNpJDYrt
Yb4W+FN+femh/38WpQqcyTLsgDVEdaz/KKVrPDn3JkMg9kYftLyP44spjyKVY9/lWS9KqI9z15J4
HG62xyUxt5hZb7nZop9q4unThfEZQ372qQ3EVhTiYiVmuWPHUjkiV5vK9wiUDlh3VD728hkq9CnQ
iUl6zCFFv3cXrgU84NzjrybtP1/CEXWJ8i2BAOAza7bLFfjNd+oFC+a3FG6gllDJPHSD04Kbrax3
6BtvJf7cbln826f0B6gn3J3wMjsmX4hNXTeQKQ9xkQL2zbixsSJ4LypcalFpTCFMR59VyTw7EYFS
jsdLYnik/93W97oWRT7nzJ/2sH4rWnJhWKXoAb3jMnisbd/Gqb2xY8ThFvchZE8zngELllcjdVm/
CB54RjeASNa9jBQw/XpmAm1706Zl8Y+q45Oqmw0oxMR7+vrRg+IkAeWAA7SpIvd7vMRjQsYs2ATL
Iaunxp6KC8g2V6d76mPYPdSGttWhk9HhG0L1wb9+VbX/Iv4tObSv0xQ6ATKkVgWFThlQ8+xS6AqE
xRkmOaOguU9x7irTXD6AismDDjzKSDEavzglO+Nwu8xf5ZgCqz8JyE/dyoZxlc3LWH/8xlBjtd5t
kEGFXpZDwA6iuqlSp3n/Ctvm1a3selzJILEZj0JatDb7N6wAyoaAoqdSseRBfm+1tlTVtWydnk/q
tW5dYvpBYqnaoNOP36MfCmajmqVp/tuIFrCuydl+nzBw/IRAT3BIdt3iYGSSAnkzw4MviYPjAIqj
i1s1G2C9HT1WqQXAhUkIIWDyqjobE66uvXqIsN5JQmxVcMQzmoAkvHOPpACUdsWSjeyOpk834l8E
6kah0Csqddr3w9gc9cP8H02FusJ8uF26vMpzXokdjdCPN6DLxNG5wptI+3aFWh6t7fut+ct90HHT
IcYoH65kP2MBFUWsRh+5DqjoB7v7teX5w7ME2WRu0ZVqPYjDo5xcCeB+R92Xb821ayQWIeWRcE5s
xIilIMC6gtOxi3HA7S55V9+P2e3cskoyij1ngiAmBPxEr/pfxGsH6aztQGERKABxoq6zjhow9xhr
YygunVkFIyxS1hVRsI8eqo1CfLojZY+Dfxr6SzZKAtT/iimhsFVhQ3RrwIRcXMQ/4osUUEXNbSHY
Dg1WRzZrnx5GodJAclHNl9iKarRlEd8FxLdXJI149vVHpzKfu+n5oacvwTAJshLC0PXyavlyN90o
HwiYLomHA7GTP6WjoGnEUj3TzettL8u6U8trGhcpSAdQIRtvNSGwHbuIeBpiuNxxyMt+BmLk4fnu
ukMwbX7WwjZiSPTpIZp2J7hNYZTxwU3Ze5DU0PjZ5N+HHItsQYmC5bL9M+8oHVEo4D9CigkbaqAU
3fCm6IMKDy/+M12luR8rs5XxelWiKYKPfvTapARKuwwfktu+fxsqRlJ3/5jbXYHRfFs339Oo2HdX
6+Jgqo3mMz5y2b8RM9kkpmxbTsM3Fg27cllvBO05jFDJ42VrEBAN35SqVCqGDjLgw84Jt3vYXkzb
MKs7clk3BKS9TRLaNVBh56H/Xt5m0Z2BWz7gOru1v3lIUAZmEWSDF4J/r3wRUD6inHSchBFnOjRQ
oFQYfSyWYp0Opz7RpsKp/hOCGXkRRO8bgoyAHdXuSPZv6p5UmB18bGGp82OicVxnUF0SqRTc4TUG
7VKBfD2OhpFN7QYOY5oYgMHHMb4AQkxoLiTQdSvKf/P++NsjOHxW2ZLRfUb4ZyAMWQirn/yb53UP
rlH/M6RwftBWTESX+UNdpxt7DugzGhxcKzqUueqBB02wTUbGKhOEbZhT1ZRCnPnsmP7ikHCF3QQ9
3XfHYBJRMxwe3NuI11xXJWrPEv5Za6c5aVFGms7Wp9Ic1oy0BR5ZJi63a/BQbYKrCBNqTZNMygOt
6rtYSSJhPw+DW94V7dv2GyMHNsSQBay19wtorxTLMSYxi8Z0bzwXGf3tmd21AvrzEvX0omcVrg89
qVlqyRGOytUtJNXFryQZWPOvuUNjtNIz7k7VkqGHFKkE8YBEdJrhm6r5aqyh3z5jEAcrvhTR2AHl
7NWaMhCmfz3j9Ft731D/T+a+3WTYqytmliXjrM9spKnMZCW3a2bzI20+xqpojEfTr0ZGRVap7+MQ
PXBNnLT9JV2lr/1xbXg4/z2GihZzIdlqq4AdfwL1JivRloaP/x7969hBGf43dVbYGbPeqDYMcBDh
eb+eq7xbmT5OKxlLR/CSgSZJbmcB6pS9njD1F/Ck1aIQgQ94tY8nxkB3rB6bc1p5IH2OTlrvG2O9
KRaGU2TzIyp+ba1QpUjSSic5N+MzrPPaW/YEQqFPvsFFfYxG5+mhfwCCnlOKXRoopwJxeecN0ci/
1T2AF1iUWymKa8yI55zH4qH3yUjOxJPXeLu713UpjJtZBSCQ9Zw8T25sl3Gc+VVF/5UdgZeFBKfU
aP/mvQvVdit8VAXHKpAcImfHyQukVJ41xqt8BQAN4pFfqt9ymyzaR1FiwhqY/agHPquDKwcjVHUm
dE+NnbswQzv6bXPykNIOwAraSuAepqFM9A8CxC+AAmONlnz6buCJ5ouvq5nCJaea0pxgSw6lKW0I
4ekiO4G7neNc62Pcw4eAYzoEkRSPkSWxRsMb3UOIXAqk7c1EeqoGOjRAV4JzrmWJn/UFDM9E2m+S
4GGUKmxlsIwJ3to7j4dRuuTekZ4ne4PnNZ7lI77bCvIoNgs46y8q5Lc5TZKb8YPPc88J2K1hlJQu
vIJEcfNq067SSzdjhsSn/tZDlLmCuvhpWBxhrKhzdEQd/lomgbY7ip7pEFm3mYkLvhaR7WjdWHag
PeHN44CG1pAkrhblpvSgBCsAXWCBbXUmu/dUQGZTd4Ws21R/KpWWPl+iPr0ECZfY3c2Gg5zYS4Qw
YLn+giGahqBsnW+lACYiB6eVRekRLjIVn+kRdS4nhxnX5cCi0q1eJowGLmtXQbNiPPrD3MKRYwXd
g1Kbq7e2LzyTAbCLNB64STFDn8Owtcj3e+hoQaveQJ2momIUEeKn1oiQl5OLhr4tgNOryZFXu/6I
4tFIGZs+HYJG51HufyOfG8KtdvZG6gucj5hybdhxDnloQ+jOS7q1ZuxA/LfPfXPyXfwUgpP0bMak
uyLy0tP0KSo8LvnPL+AkQMmwrT31j2NUO+aS/ZFWcqGSQ4wPc2kI8stGToGLj6h7mJRPlLCUUsie
ZLidxWvtVBHUOHPHKPtLcMLL/HfBub/0BZdPISEfkk3ESMjIqOjAncAGX5r7WlEVoSByZ3sxn0+6
bjwFu7tM89EhqGTQmgZabUaXxV+U7nce+/f07K7hJQIaguESK7VYO+1R0oMtcAFibzd11K/0Wn9J
TWLG7PVlBhtnXwJsy3cpiBgCk2Dn95UKTa+0n22t0kzWNhR5sSEHuSv0SIcEmQqhkZwoc1K56NlU
nkzp9mlZuLcGLAAYBhCsMTBlBOheA/BUqsP7p+sR5l7Bn3PWfUNqFLTgHqhYhuyP59Z3E/MC54EV
dhf5GgI2pmXQ2LwPgVT0ROoyFKICWA4x68kSs8f7bbYQ/LdRU2MQOGaQYxYIJCRt3tP4jrkOupsR
f+7PDes0I0Clr4N6sRSLIhdGWTGS5/8+W/oYEcL+ue+Wuev3CVMYVEvNnIZVSXALV7K+kn2ixiFi
plrzoVmGp2yEfxNF7WtaSTx8mqqq/3MDBY8ywMP/MVrc/CDIM4PR1TZvI53xmaaLWMbqJdEoMrMF
if1aNnjO0KuzSBUbNe9gTjJmFUJn21dYPHpF6Tu+61Da2jPhc7/8U3/75IdWbZJ6VUa1D5y1Q+To
KLH77uqt8HK98UCc7QNUr7znf+KVfjlUoFGsX4L3rKuv3aXsWf+Qi6zJ/T07nA1/hPpMoG8hkSy/
FTEsGNKGTj5dRyRMFdCRoI8NtC9zdLt06iQM4WMLK19ZMc+1c3VHJn5sV0/GAdnVqhdr9jR20gtB
4HwjVh0fssHuIbuQ0xV5RgmZMfw9SBOQ613TMwoEgr74o+P0Kps6xQdpvby+jV+RI9lQ1AZytzcu
9OxB2zU1wg1VHF19GOJR/QmfJPWSdGDx10nTORjKnVM4eXvLCHYMMsjGYFZSC21Vk6LbWnMwaOGC
TY6vimF0AaL5v3HfWhMyB0aNXvZWyYdObp8W2WiFLgOq1MXhz3GheBiFuKuZgmEZK7eHG+CMGvtv
s+T0epL0grRnUvQ9LqRMVe8zImQ9ZL6UibTTVBjoVk+EsSxGGEerExFG0SP1T7YFMAuuxOK+nSzm
03rklH43MR46wHpjzDsp+q3DAZWmGgSVCt+2p2Azpv/O8EVBO1U+UOe98WVuazgC4jyBIyMlIQSh
7ItQnt30brwQ/umKxXvTa4XPpykkM5YMfi03ebYgZfVSDvBso4V/cWFnClrMw3G/35irhZF2K72S
3KKOMTy8MFn7uXDEaGQ1d1vZTyciCILVp06yJS3c792Y3NFw/OdxzzQLsJNTUBFtPW8hso1HmiVz
8UnKUZpSEIl/6Yr9npW8Q6MN2ZA3PkjLz3YhtpCVCTAOKK9IlD3r6SUU07YJ0TsMxFsJ9qw0WsuV
2qRUVDJAEe1xBypb+eylTxPByghtbkXYEXssMBUPVNDLV305kgsi29+wdiNj96m7b+1Fu1z4v++K
07m9t6m0sLEgv1Q/LiufdR2nFmFdRPytOuQZLY4+0L3tKVcP0cmSnQebzbenHPHxVgryZ63vl7nH
zqc8M8zQl1f9Q1JlPwR2CHCXMz5JLNoT4oVPbZ1e9JH/otCApr5fqN0vmIFM9gNndpOsHqtvH6Tb
sI0lV6Y/xRUuC0QvFAAgh3QbYhKGfkbsBHZLLJgbpA8YKmi+cPeeBIXt4IUzcg3DnAZ2u6rLVaL/
p/1smrv4uKyTYzjqwgfj4zm1Qlqrpmdlp/31pUiyAu9mbn0x28xZSznFJNqG6USmpd5CFSEs2u00
0siZQLI/WBrfV/FROZE73JD5R+7suYSKuNC0NN9dNHmjYxy/GnaJK/NmsxQA6ThD/ofRSNrSntrk
LM+DOTZ4wScGpbygR+r2ai9DuNqVSNaggomMHV682PxiDTUFDd5aj5J1tRvYU/g7AeA0oIgRdneq
v5CkEj4OFB4SKd003IcdEn4QKUikBYd2Zucn5SfI/ggaeW/aT8elOvSh/HqM9XZoamohcEn8Jz6S
Ih8EDFnB9pWqxhzjEKTVPdCUSPP60duhbKDR5VlAbTAfao0Cm/iL+KwwaIWdywsT83l1M8S3ZRVw
B2GsxkLRPBNYXuis8BGrx1r1vhExGDBE6s0PuPIgtAipajYYx0yfPqPSZvdoIF9/6KKES3gZMK5n
PrYBUKqdxslAsmvlAb1wyyy2t7tz3h0wuIaFBu36wQxmE/3hq6embks/+CRkjo27EuvhugnYQBuY
y3loZGX8pPib4LRP9v0cirwjSSLA5cLDYBCENwbR0Sg+qBL2fpWLogymx1piCzRvPltunFH+eP7H
af8kvHRdDVn42Tta+0iIPV4vslC00fEfZg/BpnJmRT/ooqGhSBeo0N88cT7b/AQS/umeMvtp9rF9
YqEmXZTsP/1NHi5vemmA9le4jYcDH/zxdKD2bNA9NCoZnLhvk4K8eShN/phFuBSJ6s2XIo8KiwOh
ySlj1f6UmEnNdZd16dd4W7H7KagIz5f4TGEMNJPyvkapyiDmE52wynCHrlnY4jSs7ZYekGfYN8nO
KWt2nPqrFd/r2Q/3gH7E4fwkrkcpu3bT75U6lCxOM16ldrRes4LQMn03goItjOMHz0NNzfsbqFYA
8J5AFSyjrmrg75IMQX5EO2SwwH+fBunRZ+A6GP4wfmsIjRKG2CwRvJ6wmHDJm9Rm6jgcGeyN3+Ht
S9x2znAcCR21CJbv/U09G9QIVTo/iJzKZdzD5umn5Ev3vHaNjgr7BYZ+A+eFyThPnbwOfwcfi+8E
WYxnVYReNzqGnzUFQXqulCoQPAhC4OQqeLDsj8lBXGD70fzlnrGoOC3Ve+hbZam40tzRASlLqdyX
VSCse7tTtomHLgaTRDlAUrdLf1fbxdPvT08U+ScdNr2rAb/xi29Rnq6w3ANFZeQfMWr43GIDX9FF
AFLjJmhDJ3rwlrPH1C2l6awsKW+g0w2eMDiO5hLF7EIu7u/vFjTgreB1VHU5wjho1Xb//JGEENVA
En1eZs+xyzuDUIxNOy1GbPqThlSUq96QfB0IFuyb/E4tG4xphlkzEgtGhRXU2vOseBiAFjdJxpib
tO5x2PjGW8E8EnSaPTT6/OJkezLI6cSqdCqimzz2TiVp8ty2LP1iPEB8ks5nw8EyTQR84Cle2luX
DjThDvSRWanQGh4IdCZmi3H5op8l1p7h1ekiomxoXqq57ejphX6F+wNnMcfO68gKF/PRmlwlSTbp
IYTVimYCKhL0STmVxLUAndZ37E0E29UmG2NTV5if4f/VoITRQqd61IChmwW+onxKLDEg8bdU1ydi
gO0Ef2x1oDcVRILVsrUfdjTHu0hEWszw89c3KNJXQgfMXPEK1LpkBwlMCDJKbDRfD+aMFjK8ArXZ
8kdsKSMu4Iy8XMeJyRGyp7qWySqNDUQtfFFRSjs5vSgtZJVqOyw/RNli4B5eZXq1dVPOL9i4e1ez
djMs26jCakjih0OE9IFfUq5iAbEo+PjTN7bfj3y8aTJ//1a9J9P6bcGf3EbXzLIJ+oogUMJUgIP4
/NlG9d1rqcYI5ZHfP5+76N65Cvz3g01iVcMORFFIfwvrsZwB1848Dp/NrCk2NuUIht2KaJbTlMXc
i9vFXHI3/WObbJ90c2knPIqo/IptHxtev6+5Ci90J5yfIm9jsygL5JUtRIumUhMP5pEnTA8zYggR
d4fGnlKLkzMKJmVHPo6XGot81I7MyDarKMQLjI4OIFe10rX+EX4Qm++j+nqB3PWabOlCCtG7KmLH
qp7oq9JxBpNQdxilJw4zZYCe0HjWS1RMu92lN7mePcKD/oR7owEHvSP4iM7cFTlgGfX1OB94FJ7g
Jah3I7itN8pNjpWykcID8qcbesUq5+PJAz6orgYD49hddgxNABDzX+r2kZWbnDNjO7NTZS7etABM
Mw5faYzUEfzWOAq/YdLkTRnXW0KChJIyk61Tjr806JIINkramgtHsYYn3NXIVWjOIWEqlGtgeOdq
Ip6U45gTUHWh/BY4qOPpjlWN8nKHrl3G7c0ayWtM7RTafIxqEkvke8reRJTM24U/PHZDCd7h+BrB
V1Y2syCv6Eat6AIQkgDZo1tKNXZV1wm64wv3w8wbHqevcuUV9HquloncQKrHPPFnQnls5eAyAOM/
BA2TyIrofXe9G91IyJblgySKQhUU9yJJVSLUxssP0wpk5klSZSi9+HM6a72uloBgDS8H90bE4Xzq
8UBz5w3QjuwRM88dm02sXrbQybjlkctA44pUnIzqL/r22o/bEOUiPa1fw3zlnToZee68K5ce9BQf
0PHUWNLT1G3z9HxegtSIjrDwYhN2DkdjHynztRaSWOHdVAvDdmhHhbp7T5xMpF6hf8pHUoswP5HD
opyMnwpTbIbQMmis6AHrIPHxsY2Adfwm2ejNr5MzxyrYpeYPEAE4kNFlvEHrINjcgYaltKc44Exu
WKzjceLw/tX31MAr9sd7avHPIwQzdGlW4TAYXzGA5YOYtYSyfSs+GrH6Wia2fcq7UGxurSVi0Zye
ZBBm9cQE3tI2IFlSxXT3V7VFiQy89irmgWlA4uBIVkbTRdB+65X6U4k0zbbp8ElePzIp4qRdcBAY
/sW56jxDuEFKl/wByzIhluwhxDJEytjig93+sBdvwi6+q+AklekXSHBidX2D9iioXLKyLRGxWFM/
puhbJ0ut7HLPAiz0fQMnTSbTrJ+BEfp2clG4aCV4tBAvj2h37qNMLx9wgnjqjIfvbCP8YSLV/VwO
xGRCWyiS3YAxxPli/VyD1DDiUWGOhR2Nheh5akOKjRsWXH5emlXogzVVv8WHmdeg+gJA62L5Dz0+
UXNvE2TQPgo5lpJQhHvKqVVz8mj5mf/6FxzjpQEPv137/ujGx6fw5xDyOmZZBjEWwYzeQDCr8eLv
DFPCp3cYoUBrn+UAEYxD8wQQrdT7bNe4uEzS8GS4puCO+8JEWC26j6pxUHpV3WCLLjXfXHSiLY7G
WulctuvEzn5fYFf1T5cUskBD4fV1Vgx0Fl9eNi1Pm3KSyvcvx6xWcV2Uvzyc8bexxu9jObzOEBPD
46jOxpRVqopaVINvl30g9Mn93MSNGHvo3aZasaPWHh3HSnL5Omt8DFz5ERXjrO0Sx9C2T+5BArBJ
LFEhG07UUI7MCbDntSVGr0Okqel1aPYb6OWpnFoMiYqxDb1bTjjpgZ1k4iN4n+GWELnLDjLqoyi9
uPpc7AosqAo79dLWVV0aasyFWzdJHJGRa2s6+shaprpwKnBOJ2sIAnmJO/vA8zIbjLSH/iM14e/4
fLmZRe5bVIoa8jIlkPP43X0+i7eZuVAFyrflMw5Bx7J4wrwV9qbAN8Ydz1U+JME4ZWirRLDkdV4F
UlfRRqLRvb/5/CgC0zLbu25dDJ4lJqZPDhvTo8+gy9UvZx1H+pZkrqEiFc0/wSfkHYeYM4UEmNrw
psD93Ia2LWNuwYFRYjY0zMPBM+V5VCXrAgvuwaDCqmVMUjnJ9LV8BqxssxIH0mdct4reXG1VY821
FJZjbu35DRM4DL4+sCzz1v/yaKBByyyYZch3YJjpIJAQmmxPsQkfjSU8x4w7mRAggMKPVpy2UTQ5
/3SyCpwp19RA0EikO2jNLEXAscjjoouLosjMA4H2lB8Q3K028c+70fTm71cQFVk/Ye4Et8Lc3x9S
tW1xTuq45GLgEfcgkkoU6Ht++kp7S3o7r1cxWNm5ZXZpU4KvX1iUxTg8Xf/AspDh4rOR6Vzv5kEL
otphMeOLA7qAVtK4lesXGc2RbHaaEta/7ToIpghnFmWL3b2tDpqkTCeRB9EHtkJYR9HUFN2XH0R4
LgROXDQoVY0UtuOvnnbGjai+2LpMnoa2h/semU696kWNusMlGf82or0ZNuNnLm2l/98Iaf4hFsyo
qUxvOdNI+szRWtPvxbUiGtu0CUS8or99nSRpTAnZQ0j+nHS35hHlLRuqmgespdW2Fgt1ElVtsCZ8
Y9Ss8pb3SACj4QQkqiLxZL3nS5KvkBGvU6B625O8kdKABCJOfbHkNURaNvaWBTz6UVdxK78/cSqR
tiWAMD8yCh5CcpRbdtWbh0YRuoL7vM4M7aQdqooo69ZFLqpaE3o9ouSvmX8VYka+1FdyRP15vRTN
Qf+GcEHUNY8Q0rMF0b4YzlWJ0zuXMzULV2njd64v3AFnvMZwID/6+7sfK46gsQ9Ou2XpLyYYj0ac
7R8uGu9Z4RDGrdo2wwXDctFWj+oJSVyaaUxOFKPnoKfDP2DVLLKQJLTJq+BFA11wuwanXwpHYUzb
yYZ5fMct7zimqHzniMSiQU/qzWKzLeF0XPAOWtKUVgHCROTddypLYvK/xHXvewWZBepgBBQbMu2Q
WEIip0YFBDWKRKJqFO6aUWhNdmbWwNMP09ZwpooJo8MUp4eqOncOvcE4ebi6UfXK7Gg0k6qINsXd
PFYWhyh0oQ7UMAMtKRp5N2T6YpqeUhAf8WpxLQVqFK9LmwjX+c5eDf+xT7cyPTP1tOh9uqkNTTbF
8OZaJa+Wa35bo5zrTVzEeGeWkz+kenEdJkr8Pa4QJCYkE/0v7KNfERVLK15Ic9CcbFc2JSu92735
54o045orpDqKS6GfbAPqmw6+dum1hFZqtTfg7oG1Lms6tYmMXgqqFMH58OVVvz/krL2REK8q2M5n
pu+OiFBHHSghnFvYXPPM2wzKsziMgzE7GKO06cuuaemcwRfFydJYCYELkC62mbXGSzxw8Cih0K1u
uOcJxdGU7rQAwpGrIHe/ZyKwSD2QV1TGgWN0GULKBzL0xqKYbAdPM+83/RepwQ4TiuGZIdFrzxxM
XReJrssP/31NZMVgemUnz5hCWCJAVoKi3QCe91Rjj3MV8C9FjmCCSvozS7JLbO2s4OSd+1EOI4NT
qsYfNAdYEOOMQ9IdkTAb0Gi1e8saiX5fApwU+My8Fbe/al/LBEFdv8oMKm+++ntIIe4pZ4fBup3v
Kc29U+507BmwmasxdxiyVYxeJcWQjfRsovV4V3NiSMi9WJHcpf2X+cewMIviODuDzuPKKFQe7WNG
7rnbHK7D3P79ARxllvALEgxUatyLFZrp2FJsP7fdyqqWRwkj7sn1HCclbTsIWAdhzg5dTuzDxcsL
JVDITR7UGrArB7w1to7xMUTSaWvYUIRMZkFD3x6LOqR320S1+H9LVAeQrELZi3TYbpKIv3mZUcM8
5o83/6GsFzM3KQZnjJFIA0uDgTf5qeEzm9ySi/r3xXQv5hvYzXLTXEMOBJWNqrzaHTCHgEe/CY5E
KQ662mKFEFFSe647g09HDwHZoZ7wDPc4/MPkKP0AO+NDhgE4ZnuNl5AC+m3NpyykwAJiIcsxn8aN
H0aw8n+BTzuNQPZ3ZQPBvkuDAskMJt4jVUGrC8rvhAeG6Hb2+pxmwm4pGyqusPr6BPdFhmC2g09J
DiLt6FPhtVz3KatIfqTFjcVI2b3/bXx+ehBp3ZK0moHwtCDACeovX7XSQS3sNq3lXnvfuIBEAPCa
ONgSU3+bwwAqMCll1FG8YSXPoUVtZswwmZVYuBDeHscLn8NtQvTp59nnOGNvjDdZz33dxzc49/a0
nkpSUXBDDZ+r22zTckSWkmuiAHYNIUcsir+2LQN9YFKg8o5dMfKmtEGKyPCZfhaleKpAo1kZPdfS
KMuR8yG8b9XBe9VOz/OQUoi76JPBSl7Oxq5KLCKf93YR1RZRPZjwX1R2GSKR5Odkr30Nk3d/FqaI
4JTxbJtUssLgIfdLNQ6mUOtG/b4BVOED9108gH+vIf5kzyB2DqW+JGN25kb+b1fAJlzCzNh6+Gp0
ISPmFZ3JV3jbEAWdYUhnxuze1ahWb2/6+ZL7abZhInIv9ushZpmMl8DffJLu7CJ34Dn2UZP/m2SJ
BNANCqQRVVwUD1i5IDbOr1PFKrnRpXbyqmJdRNdVsdra7YxP2AolQ/H92zSuxj+RmimGjmMzrZGW
broWQw79+9wlVYnuIg0waU3ZtXACX9oa9nBWeoB/v+l7MCAJe3VDxnwDA7pesrVj9uBzurjAbF2/
a7qGDp+izj7V/MxxQ2VZiPvgJuEXZZhU1AqS7jxiNtjuCY2cNIdZXgKqwPN9rFhZ7gJ8WCgYR3Ex
qnmmOvSBNBNXqF1pB6BtMfDhrZ7zmoVsNGsEjIO6qmGlgCBlOj6nY8YNpwJPskoX/P2LWie22qEE
KQUa99QO6oLF4q/prIDmqVkvIUOE/6dmhl1tOp7oqEBgz4cxB2HxnqS+UC2LuuEs37+rrIOJeoM/
65Ejtc+heF3WxETwgmb38cXxt7m9P25M/+UTaZZjRaq2i6NtNab78Yz9MxbA2XBJQfiD7fVsjoXc
BUPGI3XCakfb4l531VNIV3QuU4AOlBjMubv4vLMQcO3FeqBNpIBbuDn8jh1t9//xb1Q3cR6dUKsi
f1bjU6WsTiBkxjSL+eQddrjRcY5zFvVUII/TC3yOCL4BnI6smEbCFwbmx50ZgJRquExY/YkpV07S
xEYk8O6t2bngoFVE7+vd2juuZogTzWTI0+tuD2adz9hZsLHEDTdrU9IdDMQa6si/OBJDfUTeBcrk
oo0v2Y9CIleF50/M4uTEo6478g+J4GDN3EpaxeeDbwy/nX0ZZADgW0jq3hA8avNbUEATFv5E2lj4
Y0Mhi2/PyDXu7martteD22XOujorYwQ3JRA1T4sxPx5lbU0bvfq1oxi+BWBnpx8HCS/v7omY3xdc
nUYU2rfxbYUrd/6gTuOO0GT0mDcEC++7otv7kHW6/MZbltZrvU8DlcUXiUbh+DvsirtNT8LWs9CX
H8WgQtvOJrMm4g8c0/V0a5fUG08Gu8zHNMe5uSiFGbdIi/Q4HI7KREtVCgdV94KXyvbLr1sB4u8h
32xHgz5U3jJC06mH4rbW0Hof7ugZ/b3A+xGeQ/fg+evCS8AYFwhyzFz3NFeu/3MhlSpe3WxN7lrz
JQvhTrb9JJNlhBLhd5EAr6E8XMWb+/Z8Q00bORV5HgCXH0OCY3NCltlfOsnP+NGvUw4zbXivHeoW
3aaFYffis4ajMgCA4MZnMdzcoXmURhqIu7cGNMNpmFYNqcd0SHVIqe6lHq/ktRqYweZpZpCOIKx1
owcMTyir5c1B2+0dnH7TOhg3ZQmEx/sZhYCR3Z0jOd7D3KmDgTEhEZ7G6SpMFpRbxo7vYGVLjLLG
NKQRAGCvAbe/I2KF/2SjSYbSUZ8ukWSSJm/qeKBa8bR8Udf2exB2E5w2YzyeK08713XWUeWA/SaZ
5vZETeO/HpimTSyf+LKNOkk9xQG/dkcP0oQJNGsYRRzZag+U+BoxbjRJF/rAn/cfCsNG3WPrAQsQ
RqAhRDNRMPE8K9ef4mNrZqqT1aGXA8Vvkv015BZE4ydV5mF+uj7gRWfIJvBIoWWfXh0epxSUlDXc
3a+Tmun1BHxeL4ZiRcmzwjUgS9yLAZj4wvfxvZ5RZA+W1Vg/mPQSKgYR5UctWCvfdWJO9m7cF7md
pvY16IRTdhelF3NPHyzZKlB2g33nw562OGLqgsPCsuDEG+wsxMAnOw8eDFterQLdz8ax0iIa/0uo
NvVF5toTOb90PaU4XJBw0C+e5yFW7HhzBIdaz9PXvUKyXyMJxFM17v03U/IiRmaVqK+IniQp4oxU
atXrXJJmSTvSdZ6M9evrK/rew66ChPmZxk/dMjUPKuafDAZ7/GR03dt+phRqh9UtR2NkhOdsRxnC
EyN8rHLadtMVrMVRWR3iODI/94wVY6a4YQXwYvq00EhCJScRERiHzU3VydLwDHQmJlelqRe+UJ/s
ywohLxEEnhpZDxj7fK1UifIARWdYnRjnj1D9wKbD6km0+uHbt8g7oHc2oM/JcpNke2ag9DzFIAV+
dswJaAgV7bwg0uYDXw4AevW0qzqGSdH2mBuxrWkJUMdlOnOrCS26Xg2m1QQ9jmxd3PRHobBQecU2
efrN+HPAwcY3tcs3zlt2EpKdh1dNvt+Tkso9rem1ELRA6yWIXwhxXSqvUpdoO9G0jV+je5+xiKcK
dIvvic0O+IY8GUW4KoBI+Y20mRdmwwW6DLnJNpq00t3nb0lKOBUL4IWWZkXv75TfvxbZqIAmtt7/
ke8h37cgIfr852dzA0+NMpAcBwJ8nMY+jFQkVg0ktfa/UHeE1QCDkXazcThTrjCaSfMhlCrYdRDW
0on5j9qQ4u6lDJWdhu+mMifmTQwUZBLecCRe5GKWCjYwPf8hqgv5dcDI4LVScCZkvrGs9e4jdpHx
at9SteGLy57ZmgZkJ07n6CZHhfnze+SP05vk4U0/bB3GnJiLvbtNuZmiLVrx7onossL/u1+W119C
NgtLk7Zi2UDk0DYVvS1F+r+hyphVAA0gUfotdp2fsYNhZfWzbGsEElsECuE94IXrqk4uHeYNXBNA
A8xgf/RxNK2N8CQiSrbjKji3DZi3j5Ic4hwAT0moQiCy7u+XYMd34GyVw5x/cHv+TUqxpXIjMOuk
WH+b6geuimXzWXksCtJxV6f3jWrOOXrkM2HRHo4aCmEQSAGvWvTTrb1ap00QZvvFsKeczAo8wCg2
GdeP6gD6fBVZ1D63DkhVuCcmgVxifJKlPAq3sGl7ngzXIJS/d8ymxJAasiPRa2Oi/DOR+LptOKx/
2TmvumCKFNVFW0uFc4EvjwC04nFvywmA+dxVxtyZQRb9HOPri5a+Ly6J18+uI4pRLPqbOfIWhH5J
gIyxsbkziguYQE9REnPyUlsre/kAYYSUEx/iFP4wtCxKV2gxkwXyVd40tSWRgV3ibzfEsKZ6+a8v
iltXlrYqLRCDThbHM7CKrZzIesRN/4g0VWP98/KBWCe/REwcFZR5gx7+hHW+QdYzE5wLQuHX96og
DZK3U4kfgxr964lSYqJIK2IAhnZa8r1DcyW0rfoZ5hmJNK0eKJy2f6waIW5gUoREazKDlm14jL7Z
jhQ5W9m3z1XTs3i559Pwc2tIBRhegtyfHeTPk6/ZiMRT+EBJAMsvPIZu6kbzZq2VO4+Q3vY8gChr
8n2f2djLz88VvpskPFc59dTia4wE5QJMzuse6U/FnAlPQqLZ8Bqi2Is5fBkiRWPwkqztrdBTVeYb
FJ3isRTJD4dcUKfGlT/LLnJkTmX/zdB9gnwSC/TbizGeVuL6wzti+/7n0C8vqW4e1HRkfwgMSpVp
gQJao2jogI7rDnEQdQchIT+1NT8IhV5P0m+vCmmxjtxnuph8zH455priFHwOy0SjZGiEmEDtWM1x
XAj/vEZf2231xwUUVwRi/YC6C6rNHVJlHjG6oGcvZXCSgvLxMOVz/cVuIEN+iCKYz+aPN2HX2Fql
EV3Jm8asew+AxdTdlFYTwRALLtHzPz/3cu5SEx5C+7mr8vJEOKsOLrz9y3NDpnY6qbWNFoti2Bxz
G+WOZsK5onJWt1JV0uRnA+y75LOHhSYc1g/gilR64WiQ52a9wHHn14JFqOZurZTOp9WKHhw/D8nA
VF9yApzvGhkGBDluaLLul7PY9/NSMpyTnaAowJAfG8zXXZgvvZM+r4hRNUjcweOci3CJXH+rtjdY
YYWZTkA4lWuqFcmiqWBv9fPwJH9+d39eoL2QZY7HQthGseGO/58tdiQmm0xurXE0Mkt9cQ0XWg1/
LwJe77L57SFCwMpkKOCRk7XLzG3+LmUHQXgqq09kG2UM7jKS6rMWpXxr3AH0wOOwjVhKScIalwcX
WFgcqgmEz7XE1P7jotyX3Ur80XxtUUmPVi+z6gsHDg+zdik4KQJyPOTPym51qroM/3WDbbR2ZBig
8gn2rSPA7FnOCWoqoGXDGmWRyByhWSja1TFyyyJ/6ujsM3u0F/X5oz+4uxi5/s8qGHdbxzkb5wgc
dtbZvs6bIQjvTxipMKC32EVRZARd5QA9MgBzGfPN/gXviTampsSr6+P6IERxrDu91mfeHsZK/Ea9
LXdG2hjT8na3glY9fpQFqeeS+owZpczATyBGXLqgy1CWt1MIbbsjsHmmfXg3sctlIukKpKxZZyhI
uxcs+7+l7+CoI4Z7k5hSucGMOaQoDXHSGwdzhaikfzKqNXDpbG24ZeDM5R9n34vos2JwtPK4Z2HL
Y4y0TUzXjuxFPhy7u5YC9JinINxtLEUuJpeJhnmtS8pojdWHeeCcCBFTjhk1jxpvTawx+QWiQYMC
RP6eX8iooQT4zgIIsw0TqvRavB1zArGlKmoTeg8Yp2krHWor0qKVW9BWRtPKkv+aY0X0pU7OVWa3
9B73kLrn3glcmxonnI4qQOKWW5azl8/9UHYBPaF27nO61Y7g5VPkpWgaaAOamzO1SaS7Hft4/AnR
5pTmaQhxWUhfQA89B4CNe364RbMzqufQhE8ZHPM8MpK7pwytPteJCtdja4KV+0UQxd/darOdhKDs
c18H15qoW5ESCXEiYlnyxgh1tAS5wyTD1FCNYpftALfoC3GobVblkhpj9H6n4Z7A33GMSwLzcgvp
s19YnoLCnM3wqm4Ju5QJwBl2edsQpplkxrdHeHDemWZ6pQ/VWCPjbmZO1gwcOJYn8BVoUKf6yQDV
kZ0cYth1kXfzxtkBV5b5KzZ8tYSiCrkFfJJYrLUJKAlxIiewqRU0XLs/+u5dv51maCT42SfM40lT
+q1epAk6ub/nnrwe9pMK1d1qQomgBKiQJ58PnY1Trpfd6fQ6XlGRPKMWyWeKlV5FPln55kIpHGQK
sVS3fnENpq/ecqOXRWqStaJ4FkPYEUiLdhbTVI2+usIgDGQesgkctl7F8JnMrG4SViiU1q0fQ2zr
8gB0RNSY6ufqqDgeljAy+gmTq8WAsE12+BM9l99PF38ZwXR6S9+NRPXO6RN4eWmyIPLzUl38nKhQ
yTI6HAAJ+uegAJSaFp2qgAHvIKDe/jmSnjrRA4t6j+WWnO3q83kc36aawFGxXxwEqWshOZOQNri7
cjfU4mv3YZemYXw12WbxL4MFxb7j0L9doLSwPD2kt9KnyAHXGHIUvNjuLnrfNGBDM2K7ZEBT9q48
wH0IHpLv8jiXuJql9YIGdE+590Su2pcx6vvi+yRmfcyNfYbuun09TncD0lUngEywLTax+cdZuZ/o
3Ah78H8AqlfEpJw18pXnsxOVN/8rE5bhDyGFkNzqfgnUCxU38j/vrSZHZfMGCjEm2bcjhRqE5Cuv
0UTqHE0mPwCUz0ciQmRBr/jZ5dkGfQadia4o1OemW6NI/11mqgNpmNLBa4hWhTi7p/yurg11jONC
/k7mtsM4760S/eJMAld3Ko0bVnAb60aDz6itVCL4iGpVCNPQ61mIM7kQhjPyWBhATmA+getXfF7/
/iEm2t4l2mkphtmbryKI3qMFf+psB+5oLZK5YPR6rt9Dsgiw8kzB9mmgfED5c2LqBTGcZYAL5I/y
XTn8uX+7TdyP+MroVejkYQrAptof0Ooi07W9ME2qyVEMi9udDhMvsutsG7/QmwGHIvCN+pIDQdRP
8dHqv1C17eEIh++NVtAOajdtx1cUJWBEaiMXxaQq445I2aEcr2jb2u2KC3a5lLhPWelNCqGxOPA5
dJ0OsSV+Oo2S0rh7Tp40asHYZ9mL1pVRNhj2TqCoqoP2g3/A9uuBpRMp9jwKWZkYU7EJJ7EIOMK0
CDMUOwRvUZJ0Zrzmx6ByN416eVOdPNbeApZkdtQc2Px/tiLQ+KOPYaBww/BKhvRJWjdW3VhAnG6r
4/jzZ0ZaphCxMreNraI0VTOM+Nq/RySkbL3H7XfaCDVUniVYni0MwQ9GL15iZXTG1yv3LYBG82U3
/t6kXxXboWPbEr2MfXAoNkVxrC0IM6WH92fWaESCHjkApm1ywluDbqscm7SBZdtIXm+CniocKoRR
YUHwin39SRlKNsWXHTF5oYYSOgukIh/mMkbeYcVXmZHFaslpgzeIKj4SrSYzNotQXlOT9hyycOnx
gZPzFn8UJxNlIHKW/SksAV8O7i4TKfXPuuNRYmySh8d1onj2bwemdipT8VkAfqwnNERftn4wP8Hn
iexAGDqFzUEsMWzUQsihKlWNAJ9FlA/9TJxrDqyt/Ahhg60WWu2uwk1O8wfuSshnv2J2pnQUSige
j1zXyrXgEUbdLDN1VS67m7eq98e+mPKH3bm2ZhLa56//3EsRAUtCWkTAtnlOGJHm7CxSC05ES3iC
1n9YE1C7EP9WgEpj7karxZCAXL4BGTnoeZDf7oZIe5v8cSNdzP7Vbeh519Mjs1lAtkjNecczT4ta
cNKRCHqDOzBVqof7G1s7DDY5ojUkBMYOBwZ6P9o2SjSFzcDxrGFJEogHdPAcZUKocHJEPqW5ntdh
wrAOZYSDfDEzxAVK3k14RDEkBKPW/Yk6xwV028t7XnF12xJgzaB1r6/mxFBat7zJeNlMG2SPzOUM
yLoIKNCU4E9vapl6mGGpBB8bRGAc7QJxQUIpGbRjpQk45A4uv7pCvq0SgRiKIb3x7VEOUs8RE6mM
9bOLfHUEm8KDYeSnPSZ6E+SWWr6tgB1UwZYmbNmpjTUI4XvrxCj29t6Y+SmJvBxbmr2QIh06n1gD
4VBEdGBgomlaMznotwPGltJ2Kpoj9VcRq7i3uZedRSWBncQslFjzPUlr0YfwgJaVeyx8UBk/E/4f
veV4TWLpzqjuc9iNBO43Ymk890NFeFakpKGBqlhLscZ9q7mPWZAzRp9AWKyCnYy5ed8mnrUyIKS8
EOSOWIGoZV3JOMrzn6VL/3X26vHzGgRyi4vkg2/0Vnr0VYx/XdatDoAyk2eY6rxehfhL/tVzFeSX
8zMVE0ji+V0hffkRMz9MpJeRln3/3ygT9RSKjLyOxr4SM0lmzg9cA9zF/gir0mLHDDOc7kQ+W7MV
3iRGTi7TaPcCcCoKBBao1VBocpwbl2ZUWTaE9vM/AhbbZZOhHDe9BSXcFP5Yam/tm2RANMPNkOoE
QLtjjqwICDJCXGRSqW46KQBOYdTK77KFIR2yk3AcI7Sx3T2DwcMmZeBg5y9p/iO4llCS3GAmj+SZ
k/YDEhelFxi14kKu72vkpcWNvtDd69zPmso6a2lkhyOsNvFasMUs6mn2adLLaOHCp2UFeu243PR4
e12M9gccEN+Dpgp2rTKQ/ipgBQoliAxHeAuwUKYbiNjHMWvLW8dQUTUm1RspjI6nEBJ5FbMaC6VC
OoDg5sWOI4noTMVVsBv1I3GRTJHHMuH1zKqWvmiABzBhMgWRNymg0Rz4FCgMJ9Ysqa077F4sHfRE
XKbzSdDqCbZC8JPLXVx7C8asQiMP+InjO0SWbY2A+nVY5Sacvnv1T+rLRW7ROVAlcLAWx4JVmYVP
2OygZzYAC8GW/2ROcphd0raLBFpqPkjmX88wgD2LEWAfmuG6OU/D9QXY8+CLjX5OmAVI3jWr9Gza
nEn+i3lqW322L39whVFACx8/bVlsUozT/6BiVbpzCrfCqmYWr2TFfU1uuSVw8T0xkT1eBGp3H0Gd
9VDi+eztKuGfMi6NBpawuu5pVSWQChD09CWTR/rOQrw9YwoyabcPa2NwyOkeDi1DjCZ8xgrfZAy8
efFLA57WznJdgTOf0Jv775ovVxs/p3m7w0VRxx2bW40LeATVg7Kdp/kAv/S6UAD5dOre76eSgFTX
xDbXW65a7JR8B6mDZTk0m5OEA/v2gwSw9la7qU2qcqYhpgFuCqkGpG57E9iyJL6doN9jLXIomNFc
IF6Nj8578QTgzQN7qpJb5VJzmgN03jo1b0SD3HK+6xn6GPLKYcBj/GDDYstWPjrBlCOepq+F5+I+
kd7I2orITC10h7q1MoRrarkoKxGbIdYLzjp4OZF4dOHBUqmHvoBIvdyt+Jw8iGVWBe2RNo2uMCkC
YtBGUtg2RgIV2eEItk4JyrhkdcKlUJ4iEpckBzF+CmLkWhW66ynnB7fLBJrTUS8MnKui/Jdb0sNB
5DKklLtIGX/eK0I8jqI7JSQjjEX5cLNw/iICLfAG+82nR8J+AyTvkJqn3PIsM6Ff2cS3o7RO10p+
6Ey91wzVJ97KxkUHJCn2vBOR7HhV60FZq4TZ8zJ3sgTqD//IQw4C/zRRdDxRhJnDqA5dOQM1ubeT
o085EJvRd1dyU4VfbyjCWL/s3BtJ5D3t8LCGPnFauQuoM50zQPr9IPtpckHFnMIsdCSWQwr/xutO
K7lyi3b/35ipqCyX6DvJILH+Cdo/iTqD+dsh3RKoeId5ipTgCSg5y5ZWUnsDtuUO+4gMhwLi4Lb1
9vPBXwbg6J8Y8Ty3PBLlEwK/Xuzw6jOxq+H4+8GifQ6itOXrpdxx390ByAYdVu/U2PKZGMN35feb
FKYzt2kOUU/1j4cBjZJcHWkPBi8IUbp5AtyIaJepEnl+/w0vsD4ZNCIa6l1+gfGCH0GFvyLo5YTh
W0ZDIYHiziEDbWuGXESBZnEsv1tQ7QLwrCSVS5bQk5LvEw//5e2mDOC9bc+O5wHApTtJP0uCNBBT
xcgh3I3z8p5dTf9ct9uQ88x9rgQfc26Dao/RyRjRonPLoF7Prs+onJJnumlArZoFcESKKVXtPAwM
vgKy4VPqWiK9c/anARiD461ht5IHoeSMu3jMQpzZ2C7umeQTNwcFmUh68/d5GOvmRR7liPKSoUza
pKfiK7CSpCCa99xCf9fvIg/EAS25Zheiu5b34r0ThssHoQyRZRng+04MkRy9w43R8ylqIQ3BEqMr
8NB4t8ewbdDKKLjF9FYMI5UUDvbKLu7q82JHjHL5rW9ljoU0RenyUFymU0H/wgHV2w41aGyOk3i6
Qdim9JBsydXyseIpkJMxjNdor8HmM9sYvjpaEmb6NqInoS92p4s+dfmSygX2Giok4YLRTnrUWPQj
0eIcwCMC8DkDZeYPfw1Gflf9cN0NuxG0wqq0MVVJmYOAQRp8wIdJ7LFDy560/46P6FeHGGIe4HLp
GdmsORGrhlJk9mLWUqgjagtSbnjIx1SxPPrQYi8C8FDOb2BcY8MEv71CVNv6BMZ6/KXk51jYNY1d
KgAaqYugDpq2I7QuTikNm6FVckU/aBd9ct8lIqYVKFnFQaFlbVSJLOqfb+CzCAzK17wy88ckzwXl
yEHPrKx5DuH5JVUOG+kMAGdf78v85TPzegVzUoHBKDWAXdAEnx3YGfgvnws0lY8FToiVi80C9Z3t
SP2rAgE+0PbRNXw4tZHpFlLettQSQeOZJNotjQNgly//aXLoYGwpaHwCdAYNGss08J5LixIgvrra
xmGo7oGg9OCtWdHzzF56NfKHLmrcpXL+IgzXcjBR+M64z8cnvr0izF2wG62c+MhydB8VHQu0gzGk
7quuQj+/HESVY+joQxDkfprCpwc6zt3zTtlNZeIUEFIaEoOQGHyWobfcTwVxtzD0kNLoOuoIrTyH
AWjJsEJ74J11L8O8UnZZ9xWeAo8CPq46FrSqRNVR6V/Zsldhl7FMF4lUORvmzqN5Csfca99kNe0J
Y8/1v/ssC3sqBejryVB0HJCdgNpraVCnWXZOZlXyaFSwx6q5acBLCG2pXqFZuCtQ+YNYY+wG87+Q
IcC607CMG6AnSBa++FK0H1dKLnLQoL7LU1EM5TY85w2jfK3Y4LCAEXSHkEbAIZNBCyt2y/SF7frI
vCfqBQTT/LZTx/VyQVrskrB7DyE7/lW17aXQD9U6xFKgfmRPe+7ew0SiiKBB3NflQfC+vLuw/ig8
A20Ppa+hsFTefDc5yQ+GxO4AAmA1W9cCn0/pSEFulaDNDZszPhqNK5OzLodmjMg271zL5434gUrZ
WIJR0f7dpJZtf8AJdMIjxg+0/MiuSJBStUnWD0XZ7kTFmjCmON3W92s+5uhBGmqlJ8vcLf5JyRvt
2lf68tHUjGdJRLzu5vmdPTVxp7LxWY1al7/8F9i9uX2FOTvc99wzzzHpctS44+hWeIA++Y+lYmaX
HUXQZvy8FBQbNGufwWpsYfgBdP8C0iqj/x7ElKqvyBVWETKEgk6xHffn5FE2v2/203ui9MOZfr1U
BaZYar+Rx94IPuO6znRe1e64tFt1JgXovwvIEIMwAFdMVVXq6/CtNYIaaRvTTq6c/CssW859bUdF
xpD6Mc/GEucLT/Mr6VOnW1ah76td7ct5nDUfI/4OJtoEfujLWN4UUQrtcOCk7hRMI2YzEN6Lfsdz
RPcUWzjeCVH1hx1fA4iP3iQCLsi3QqQD0HuVikT9pwgPF9Ft2i5F9vnfVxAmgs1Od5EsOB7p1l1V
DXBE4lIKwXiCXoXHuws/E6RIJZ72KWgBxkGqugBpvqjscJto2JoZG9kirbUrGzaVwog2CsE3S7RX
db+otJG99wSNmJhO0JAY6pdhr1VWo3SxctSo5YRhLZYI+OqVrgv5Pg9hUXz+PhivXeLGERnqCk0d
v+s6tqj8OQdjDFnBZdV0AgzXWAp/qQgXNbbmN85HbPUwRIilqw00F7jYIOFVN9oRsEk2W95ts8i+
eN6rhf/35M+dU80i3DvLsVXiovYjj2IBxjD0aG8bHpNJt/JkasO2oUYac7krrPfW7h7uc1gOQJWr
HIAR6ErubcnTV7IFV2GJDpP9akPdcAJS3HQBVhu6KJv6RqpQLGCkRzq5R5ol7qs7vR067Vnx03Cz
XAaw7g18mgYZMzm5V6OcHQffGQ66Yh+x+mWqSJK1FBDgUuzJNWwwolPeKuoZWb1mRyJlBIQgOiup
0IaA0SiiDylmHDjdrLn2DhGv2wi3ypv6eEhBz+Isa+rElSGBZ956enqDqPlPR+vF06+X63g+jRtN
N7UuPyMdgkibFyv5GDnUk6WT7269s8IBPjSAD/oNiMEj7/0wrpPLaQhV3xpVi/n20mwiVVJtTvMy
fDZR9LpiC3JSUKHrjrg54N+KYGYV6z0L/7R2Pe63og9g0ZHVr+TxxJcQ5oFSz3GIQr5V5ddzKbBp
xBtgaQJ2GurVFP22x0EwLJ0+rKfcEzhXuDzPBNtFmULAclNfhFv+X0rMzpE+cuBFJvwljwYXje9B
9DnPnfOFTYdGSIgCFpE/VNruqvof4HtvlZEZKrG6i5WZtJ68JPQvG9TaDdYkpnRydpJ69CY9iSbk
9NeF+tyYF6PHK3R+/jGVzQrVGHB7TiyMVeoRI4BxNOz9N00ztVR43yDNBmL3mFW0V52GVY9GNK/H
wKhJrO0YlVTvdiIJ5ffcLMqQmInDM23zB7pncH17n3wOZj2F7vxTeY34TkpsmiFdKPhmGPtzA6rj
u3c7tX24SKtbz7HX2ReheYTiucnOw8ElSiZ5FD6fMIFSlVJHxH6Sso52wNrQW5K2+GPoz73N+urv
xKRVjfV4rngpevaac2z4byXgAIcCadlYksp/nxDo66jcj4mi8CkgoTnlh+aWCAK5YbfAMyQmrgs0
VC/yhMUYOt0DxnUMPPHI7UlOyCQNKWkOqnfNQDx7teXzaNFzxLRdCZzJn7ozIvbcQkH+feM5JgCI
JK253tPPfJcZHENZUfqnTcC8g/JjttlA2RWcXDH8xZAzfCAWs3o8JiYjmOj6rZkMC1/Ner4QiTny
uNj9QnTK/b/jbAqRPXAupQnf6wW1kL5Z5kw1HGl3hmEKX1ez2uB0x9bcpG/ii2nti/Eom5CBqkZW
4o/v0v7LbV4lTWeBwVSDJxOx/ZDCoysqWZaJYNLoEZuHb2iQzDASLRNKJQbNqy4+oSXYE6FYJwws
qLtqCeE1rumXaIrzgnjROoIrT7jlNAUXR4re+OFmmzM06tA7yE8Ip6A6zpXzzk0RwvXOf4W53sN0
9q+H0+2lPl47QrXzHfg9d0uC6GyvhouepiNsL2lCS+zLeMfXw9zjAhUDERvJC4mWLAr1NCBmvGi/
P/fDOzyg/yXLRAYJJAZIO++0wHriZJY86qcfP6jW+Hc1a1Lg1uRd+nUWys9ME72wDGBq0gzL4rbx
EbydXamY6DR1QuBGuiTQHPfwjVGb/tHQzSpOxPdmnx7BTTExshUchzyFdNcuIqkEUyAM0yJEpaJl
6lIKBb8aIDxU8Es/LpDFP/fsRicSsNM3zAE5FEvFZ0e70T8mlopJRRSsk/9jTsk8C+HQ42HxLFhe
uYlfrHTUtjfYOsx3YXEuyZ202voD+mMVOBNgDMlANy0DSJ9tkff21Qn/LoM2jaqGhq0LmjnpOhHx
4ZIgoWtxgyHmzqJ/3WQ8PeeI267hp2DPCMrUJRfG3x11Ote29ghP92s7e2rqmvVcWwC8oNNu71A3
+HDGCX0m7aslAVgZDJaSXu++K9OMBs6ZH0KhCqX5XayQiZEselgNZDXnouYk6upQvJ6oh16HTSyt
mCSPER7F22PfUrKhNm3AbkcSJfRNi85dTknQIxSy0syY7XWh/t2OKH5I8ZRmXnX/MXA8G9RxHmbL
D8ynU5JP9VSxJiRe1JYPx/HCSR3zxBea/BfKq9b72+a91KvxhjCugm/+ytGW2JipOnBSYl4tccwE
XvtQC2btlXxeg81gMjF74TdsNifYTl3u+FrSLLKzXCPC5UOLPjuv1WCUpDcOxC3oQ/0YYUXNYFLM
K4jzIcfjdrf52R3Zq7LsJGKReyAc/w19/OW5qFcttjXrBUwmKxF3vs+6VuivVQPJR6p7CsC+WcYe
R5viu/dfzFXGutn6cm1faTkAMXEBWk26sN3PXNLbr9fnJngLJrR2rbg1FPedftmsFMJknIEf1ORd
TmE6zyTDRMs8onCzdXnVJRVQn5uSR/WToK/raJXUe6J7xQsqZ8Z6mm3wxTUiIyw+Hg+oO0KCukqS
3p4KFwhKB1tQ3+Yp2UuluxcS+0HQ4Uf6JSrNEXnnadkoqTAYOfJWkI4D2k0DbU6DaHWCo9+rHs8R
sm84S15W+OlfpZ3PguF1zB1Sdpc4BXb5GvrHoddsGEmxp9CSnmz3FqEPIRpreLIm9Qga7gGy3p/a
Vh+umxEj22ao7HTh6EdqJ1qhenHPuJpKpASOIPnJ7+5apgWLJWQfIFO9tQeB0Ptf/xystaTw+XXO
NKzhOScCaTQ1tU/LgIa3tVOlEFj9uwbFZl36/itBR5hQ+2PXCXlNfQZC+ti30ShdMGu9t0iozN3r
pcgzmrcct+I94JJj/4/hnB25ZygBb6Mlz2HKg6aQrrTrPdW2751bO9OF+0qKWim0EVpPQz+oZrQb
jaG2NdzlsqH27kI2LBaOZbtoWBZ75UhtyBs23pOYDOZ7kiLcd2ZQF3Z+yCTMYd5+HY1Qq4I2Kb+Q
284x7NauFhkdsYnFd5/TBE6AVXae2qZW9kwi3w3RW+xv+Jx0/TzSKEqPsfvKxAHwlf9vbSYdVld3
MNbP77EoVbNstExmBmRa02KbQcu53YFz/OAcWkWX9GgPsoDYKb9Ml7HuG4W2zN1KMiD3xbgwwKtx
VbRy5O7V+Nv9XTleqOvzuNoIvINu+K/3RTdh8a+qAzPbgD0EjiBKjTUmVqsKAFW+UO2s/G/pYrKf
3mq7+3u3T5rwzvKY1WI5nZGiy0oCAm35euigu5ZJHvmenH13cD/Kp948ndyrt9Mgo1Tg/0jSt3Zb
NWNaNPle5ElnZTUh/WtF7MSmpjdtLykEkqoimlz0pn5vm4Zm1WXx/crew0pgn3puAvFkYM5ijhO1
bh4w1InHtu+zmTvIFh608IHeiY/G7xs1EDwwpxoOMA1eBvZRv83DqcRqBF//nIlVWXGoUF+aLFgg
NfhBHdDxssM8JFNYE3eqMMXMz6hBzUQTV874TB8LiF3hO2xxq1MfVcCAjWHn5BBhBpYFJ3SKx/rS
Xq3M06h8enWSZzVv9Tf5KBux66HjTXATaSvij31FBeHlz0brMOLSvn0/DnBDo5K4wRey7KNxedqD
6VDBbWbAZmZMKHkUEDCafShS8v6VnC2t9FRpuIKMf6x/iUCw5ae37vKFlUo9+qrQ/kLwTmqRBFIa
nBkcVHPWTU4P8HfQBvgJ83GulrTI5JMaEIBeRuRAzF54qOmiuePaCymPwxvCys+xIDHpWfr0pv6t
ZoCz/mL/p4zswFcJ/xOmKBLBSewnmVChTU4qVwMfooCpHTVDyvM22hF2xtaQMdCeH2JObnjxCo/l
ukQRwzbp/duXyQt350Bc5ujcA6UPjWMdxTXaXUpQeZFyuXmiAqAu5alz4QCp0AdCbnq8il7G8OPp
SgNbgv8fMLhq1USFM2KRQupAvqh+L4XMHDHrdRgCm6KvEQlcton+BzEN6s808srzwVxHDJi4nELC
ZCK6NtVDT1zJpV5NV9yuEDpIleE4VPXc+GqBnxrzJ+YPUOUsP//mVa5qOo+xFXShJBTAJWswXFFc
xbqaYjrzGoNIy/k+IRomywSA6eng4kCzEMItBr/ZPwWu1jLr/mY7Eoxobm8fW9X9t5QQGlJZrgi8
PaS5ySLZMTdGhEQbGFsF+ogMyDBfWfzhf1x7nwUSslvKVrfR6EOr4bh1o6ybn8h9bhZ184Qox5cx
DaR8yvEqUZmkoCRD6ka3Wfv+y2Icy3llcfZYViS66RwqlCRjzLRY2IQ9JlHKr5TWhtzs04OUzd6p
4bbN5bTd6/5arogdNORPXauE5jNm0ACsOw/KVFdrZCdpx+ur/K1iIyGA3Eo/F1qVcvyN7dX+IiC9
PkTcOPFel4NT6/lwdnd5Jd/BymYxKjI110Ttb4y9QODgekXZI5RVu2pLvVkCQ4271tjyE7Okmz/k
Z1MqvYnOqyrH3kUDaXeBf3G40X/20TWA6NJbLLR/VXmrdhcA+zb4iJDNdSVt+1ywyU4+de0S6oPa
LTfSWWJydUnT5ESHFaQNknB4L5odqNtJE6AeM+sDMFgm95/xJKjrilUX2W49y+j9nNIjOj0cInxP
uGvCAPoEZCqVbM6/lSSTiwmbdMTYRwwW7uai2C3oJZpRSO8RGYE7aIMLjL6/Po3vFFRhl3O9QT3h
cHW4A+Bx0EJSdHxZf7JBgCNWOfuzwqK7ICK1KXPG2jDEgD2Xh5OfHhklTvCG2RBbwNhVlKI048hr
aqUtwyNkKMDHOhCOZ9e6i8AoCrnpvHT7PljlK56h1hXy3s4UaAZzq7b815psX2lcgc05TDRK+Yyq
st5+Bd5JJLhfrsheeU9q+TLuf7Rzbs3OARCGAn+8GH0PGuo62McoygvosetGUAif4LvTm8yaBLRF
laaC6D3RfUkH1ilMO2kywLUmorSqDEBwtHkBHSjCFK88NiNfdCUtN2mHGyE8SbFI0Yuk2y/POxwu
xn3kM4Xky8I3ahIAIo0SQl/bVyfGGrevPb52xlQF8CehNJKM9s7ODvmajv1COaUpkr4pz/LXQv8o
MkEWSf3hny1EyJhTc6O3JdwI3ftK6D8pLRSI2oUYQ/wRNoh/XJlhXMiZvKVBnlvLat3L7tbXpRSk
1owp2ewzcMEgk5XQpMCWO+CyevEqEEQ6Of5/xTG7EtUnPAqm3ewt8JGlte0JpLKmTRr9FH32bqSp
oItg06IGkENRmvTwtt5um6YcC/VcU4VuycT+ge3MMzoXOkdqmxGw558aurL/56ROWkJJbmRxx35o
ItxDQQmTnnsH8hUGV5jP4TDAlMzoTh7bX2a0KKn+gTKWY8t3gQ2xnCLkZuMsmGKvCdjfaK+3j+M6
b+fv34JYzzWgFGG3dG+7l3ZDo3QZ3HFq01P6oARNbzpX5CXNt7eImixx1FFvIU20n6y48h1bw+Xl
DkQJubsWEzl3ntP8XO8BsPofwrn8thMDHG5Huqg4nR4mcRib1CV6y8F3iyHjt3+7lxV60SgUMy/d
FHwIiXev/tyKrd3iPKWGWp0Pfp9avd94Pm5a8+2MYMAY5NAZHlELyYpwk1ulwvbMjOzQABuceY20
YXTSPkL4rP+Z3flyfpcIZ+EjqVog5hGTC6Se0ionvSFGqjm+MrXOFFgTM5D7iEk2sRpP9WmEozKJ
tHCfnpp3qPVsv9fyu+oMq20dXw9XP4lO2w33NYoFWFNnXBGaErp5aLdwlFf5+bQPQHlvwC0YPX0Q
SsxCt+O05H3H6OsxgjW75Ny11JOw0vEmBp5uaXdOZ4j3aE/XZCVVslW7HO8TfNN7Auj1vuI7AX+y
ONCM8ACAINYAgP8cINkg4iNrey9Uk9K/QP00I+qxz0NVebgbDC6eD7Pc5Z6xCM4jPQR8Udp1U6WX
1cS1YlbACMyAulBRqVh/lSIP3+3daRlJw5rfMVOkF8785Lq0+1S4jdUNsgfsc7i+GISNj0UgfCnn
PNqg9vudtmlUN6baz0ITwxXNMx0ILxTV5E97kA301JW/AKkUALqUQLfKomjY7dt1InwVP3Qr3Wfy
GJrUu6DYQJQyV8JrBfdoPiLHKij1BA0iGUqF11W3Y0/nb4AKHGv365rb4oU2utXHSZ/eevs87/jm
BzCu9EkWYsi8RBDoB1egmtQZ6uouGTqiIcvCKl4bLeeuR8qQGrVkI8YRvqBhqgc/PtMzQRXj3w3J
918CDFOHi3z0nG2VaZ42YxXLHAadTfYILtWwOnIi8gQGUT9qCQ3AfDW1qLcKSzlL+ghe82Gwd5WY
/D1UE1cBkPgdS1+j26Tpm1txB4XwLfdswWXVsY3AQEMnyfDsh4cjAzGRW+LDCYVSFFcZVsTV9Byu
pwHB7TOWDsms/SEX4vriOGUq7uUXw8x+0C0QsYTBN/otF+eqCKNeaH1XMBmtBzm/xY/lB8MvQZwS
J2vtE3GQmyDY+bKctj/ac2te+w0pXA18jwLzqULVD22FR2LTYzfEqLnF49d8XeiiJB/UqbS8uOAp
RDh0ywLk2MBa9/gJRlpCg8BAHx2XwmxCDNjIwE4kpO1P+zF/x4U/3khSvzIG4K8aUdQwkpHlkE/j
2qnZd09JXpJECB2PFluipK98TJMiai0p3mVhwfm5Xlm8p9cC0uCjvbmk54WpkwQ5qsRziIyMTiGG
OnK0FuJy+xb+esyrzM9pP+vyz1H+ILAYn2kIxGM3c45LoOmLqxjGhNhDiImT/VqOTQahFCcPfTsY
ZuqEd/1ckLJal+t+o17rSchl+Q3V3dK+CDJZ6dAw3sVMmiL0QVuj+Cf0oOu/tTK5d19Rqp3+SD9I
xUodVIay22s1Wc6geRD+qqWOxI5uB/sey2SbuptYSp4mugwDGwIaqaMuh0gdpbxrHpPbPcExChka
NwuK+m7ZuzVIw1USy0S5kaavGFrdcj0kb+BvpNmu+8058SybL7lqGzM3zbzJIO1wAudJBSeHB5Iv
DRaKz5Hv4pmqBRS/9pCycFpwEHQrQzy0WQKtcTGSj6WYb9ZP2wZqFsp64W2jv/aOJ4j+SMW0tWfZ
NK5SD33xjxPzT91G/yIIJol7NL1IddVBm5V2F1mcwadeFN9vovZzVOuUl/jzit/Zu2fvK6yKigLL
bsBZB7uvjlc+b+ZSq+e46RWjxrC2Bvr5c1CUfEb4X01TVQdSV44cvhAPsgWfQ9nVq3ILJOQodrqv
1FrybUfuYVl7XWwDceUelfsqNcTC/sIoYWD3aLkoZmkXmGdzP4LtoOknstKOmqBm2i6Mw10ep2+/
OvdxA0nHZhaalCBHj9kSNDGzVXoGQO+98DXlq5u4cpWvJ3mzycHEeO1C4wD31q4NIn6H4rhwcc5x
0Dmdm4os/vdUYnj9Jjo+9YI6sqsBPFpCYEy3vaUuf4B92Z685vLAJDM2GubPZcIyMaf8iatjGg/I
UDSwg3eYKMYuxEge3mdqJf+VMhU6kdgkH0AU+v8/3ClfBs9QCky6ruhSny7YmDF7E1zeaz4DRQs4
HPgvNECq4X4yjN7VEPV/H2V4sNPLWEWXzjkuthr7KQ2t/ymDBmuzb2FYJ0QFw8auJQufm1O7+Tdu
D2rDJh9i3ROezTsJUEOhtAM0dbQqSB+nMS07SVDLwubGr0MMkxYssiAhSpSoDk4M0rF6Qc4ZpCdu
CuxenVwvkIBaK+7pjDc+k17z1okzU3EXdLVJUVy0OtSJTNolClnYIvffpf8XlP1qqc98xoj4T1Vr
SpGtfa+w5STBV5EARK2cpqJpdYlkDm66Pmxh5WLrnTFsJWM8hNQVKBPft/SL2KWryd8w2nqyUo7N
Zw3goAyaBDbVe2UDoItnB/lHNSlGQD4s6W8YmygyIxDDrwVgBNUr+B3C7lRGqXkiE34quhcwbkWK
MHdMmMc0aZ23eFQLvmYL4Md4EeaPZkmpoqRoRCq7Kb5mGnNV5EySz8wzhoIsibtAzDLqMa6pWjMi
/zqs0lG7YPC/6pvqD1DRAzUj9Ao8owQ8a1kQaW9HwYd+CtZLJnBM7ZhzZEBqN1tJyv3Mf4PesaOY
/yryGj8uJi8hMmHMZ+ylhRxXTC84yQnvuVnzNjEP3MAbjHsH5nS0lvO8gCZoIpfSaORI3am4MzVX
HlfqsaFsg5mEGUErD5fTdFlECpq0t1zFhvvtB77G8o6p8cg6N0ko8RvooVfeut844itBFoHKrheB
wCC025jyJdrMtq2m1B57n27F/LGa8K9NX89ZFnkF7f5YeFJbXuPeoUUQ7CXfrz/FuWmsdYhMcYk3
Oja5bDKJIb4DauSojovWtKNXPeLgSnUkb9PxZK1ZRnF1keKM6uCKmQuAah2lo0dQMYKtOv4HK7mx
pN495EkFd0lXPiJBadFbq+2qljs1hn2fbl9XZ965L1PeZauVb2mYv0GyCGKJo0Y6O4zcs1DHclA9
uhjT5jOY6VHH7QoKIe2NFCnxDi6DTM+8MOBsqQKJkuEeIj8haH8x7pqQNl7An7LGyQHPtOnuiJ8G
A9bpS3w+qnLYDvUhgGpfscLAWSm576PRIVoi2QxXYBbYt6RrqRekBy0DJcrorKRPB4x2LU1p1k03
B221PF8zldyUz48eBmh1maCznrqa2F0EZNtQfh7nRxxVeDNDHhc+dZwv7MzyaqonN0p7opOwcvIa
PdGRGCNaq4DEQgySCBdsECABJk4uMhPU+r/VDdNSQBoP4iSSEPjaD17DulcH6x2dXn0XUH/O7ajK
OWEWJ+a9CUXMhNTbPEAYbEcEFJU8DAimi5VnsRoSX7wuLBpvijjzMYoE5Akn/lfH+Lq/jIGlNUZQ
8U4WyI8tzUvDR0O7jiOAwOltXIyd9g/NCxYp7UUDnBdbsgNAggPvzqgHJ/mHjIkwO8WFyEEO5tPD
yBDOft/IucVm3VAZDgculrJ73ZLkcAaIN7mF6KrDhHpq7YplJAcy8zzcyZzOJEBUqDMIcV2L5JKJ
nLiCJUcDFJ8WudigVHdRuIdI35Dl74mYGerWJnrqnX04WSwuo82y1rWaMwQSF3/fw2OXgi6MpIaM
vGQxlmsgvNTvgMnMMMwFw8Kn2QKTAWEbLoi5Xtb+fS1f35cJMvs+0jkOo9S2OP63CX0LcpC8idaX
MVTPc5uhe2xySWp5YeRQOMag1wQipr7Y+y5rVByYHhr8Taf0C4M4k701/nSg/vcPWQfsHPxtcium
tEWBx1HZofJfQ9cwo6+SxbU6RS1uXiG+P19sbeMzLYKAVibSlgYWR6Qo7bXPOnsJkwmBsNt9VueM
Jxbt5Vdp8dIzrCZmy6M6AZ9EGFCs7uwJ3K9cZzDGCWd2TA3ZDYu2ZSrlj9UlgslJNgOe2znXdKNo
N9e5mvuCei7tLaOYnS+b4jX8ufrdI8N4JKUixNf1em+1aBtWW2mbNjKX5FgX8JjBS1bjw4z6rsPZ
kVcO0ZwfGOnF7SHqXFwpuUcFNGZADlurP9i5clt9IJPpG+C0Y5i5cBavlcby8osVLVOyP56qWcLz
Pv2ci26SRfNCM77vD/fq/zpooYFDf2HucWJYHh3wbPC3CczRFU4dMsLTDEKnNjd4iDQES0QCbYur
LzIraJTFtzgjMYQEc+KH47456lE/U1PpzDPa7cu1g7w8VWYSM5HC9s+BWPtoFy9dU0+Z1sPlEVNR
WTeBte+scFYEIxfKShhODrg1c+D1Y3QxpZYYe9GbZrk9cmgvf4HZTr+0BFpx2edHans9c3X3TSel
nOIcalUY/owjL9z92JZS8oKcjLf7xDvzq4OgpYj7aadfmHIWdQwPPGr5wSsPpNYwzzJQSNethrN9
RFu0rXrb9sH+YiFVrcXPRGeEhkAgUwUqww8x6nqyz8L44lM5U7yagkIt8OvWvEdHJpUpzKlFzLvA
Itpgk4FEtI8UobmXm867vIUG4ehprQMwl70l7adejxhwOv/NPy/ExMNUigP+OobILlZN8j2nNJnB
fGHk8fWYfYyfzJXqIAWbmMKXVB/jRfNRBytHRztD+HvEoBU/1P+oC65cr2ek1+aSMOEHgsBlHBQG
+ohVjTZFl/sp8kQCR6oSKQMUudn9lGIkUc5Cz61YNZ+IJW7/Wm0RT3h97epD0Y3vAExxI+2B7AGD
31HBHLEzigRFgw3P28OmdSTJvKgQh27XkI8llJ5GG3VN4Pj7sdzMsMsvM3Il97J2dKtud8VjpVTq
9r2kWcfewNdCC/hGkfvQ2O+XjPIBAXnDocqD94qhsRB+apxQSt8HdFN0XyFviv11YIuv0d+0Ch9p
SJYGSvvpqow9wmAKAB/DY9qIDwIMYR1ynmCGSD95XhP0KPQ1kdq+ie0J/6o9Io/PJTJHT9n8FiBk
edMRxgMFxNZHmLTOo5rikkam7mCHLEwEDY9zdyBa1XA4ZIfTZLnNuROGAbNFb7AKDu+pdaGHV5CG
bw6U/0kykMH/4S8S1dG4bWF5agn0ClesSbn8q0C5gmG+RBNqC7haMLOH3Yq5oIOA7dEeEwwZfgdW
8LpmEZ6m3fY3a4EDSW7u1eKuP9tc4UN7VtF0TmSOJ1Fu5Ejfhin7f9f8vp7Wo58rfMFbPOS45gVV
QWmwsc5w7Q4DdN63zEa6HyhMO5dwmkIBAxT89u6ZvccZCi/XbilHwNU42AewJz1obMnxHV3D1e4i
zkAnE3Uw89HiPsLH9itwwpLcX1eHGYp9HqCTHN3aLAhrb+4oIZLRsSl6lqYUCS2TWN+iZ00ZO186
cWgIxibYp4V2E4RFfnqoeGPu//7mqmCV7ZGfF5E2qxUnUZ8Hmy3hEyoRPNbiY0CK9+bE3VJqLp/s
vols47RY/P7Hpz3Ne9XChTKlkpkDpQ1QGdORJFIO0uZjd9q4kjkbY4cC/oe7hecQqKEjKy1kLnSR
QHYwScn7Borr1b4tp+KCqI+v6ahRbsIytRpM+3+xZp85nYLeR4uxRCy423l08hbPD4seHhffel02
HYyyqG0mpGNeZRFvs5WpWQGsqPQCATDPvDsrjjHMeuWD5gTRoJGRPm275LDSR4qQU0M0PVXurAe1
QNbkR1xX+4qW0Asst/ZmrYcWZ6hdPvTc3tclUvSiClQXFooBR8aDFmgwzxUBR8T0yH+MrBfa9i3m
hu8Odox/WumNkPVwEsIdD5Ytlf1Gw8qr7pul+RTGM3geJnIsPPWYjytLEFCcF38rDtISwfE7Dv7C
cr4Vgw41uKG0x78A9QHjUGBOc1SGQxZ/jfYkZNrbxQ/7ezPo2c4EHcahvpIMH/A5jYHU6Roo+MjU
jzU4p7ypcSNwJwVnplGpzQNMVsW8IKGgOTNxcnPGoAria7v/ca/KSKdpmR+px5h3cYupkPh0HGX4
uBfrg55f88I70doxiVgX6fqU27uwjdEuiWczf3D0Coxllk+ggoQolXACx8PUc1g+dETpls3yKGEZ
lemx4GmrJ+IFDO99j4A2dLhFXWGysr17tdlwlaaN1s2anprDEgLNKCkQwHv8oBviW08aGiruz+Jn
s4fsh/QqOTydOqANUWMX2V18eGI6V12EMnjUdqXNhvBcj4ARKhbyiP+IPNcOkm9QByApMhCNprOd
QcTMUMr43TaRPcjZDAHd9qALapZjna2PcChdLIg/oWzwKk0BBSstTc0ZDK1yADghtACee3hk38XE
kxlbMu9twbKHMPTnNj/HB7S59pZBPTnhHlTLOEq/hkFVIEB8tGFmqMIOy0Ag3eAl/fKNn258ObKE
KKX7lqILFO+kPnmoy6e3zg9pfPLuIVDc+xmxDzZYfamRB3JbIIvJZFoXj/Gh/DsdSlC74LGKgTh9
HmFoFQQRkgL2pvRSw/1zC3OjA9QLBQ1PB/Tz3bV+C7u1KcdRQ1fp5ljFuXL318ELecPwZpD/xdGG
H66BQ7ILkHbMZP1t4o+9taJ4HBTfQeZzhRtfOIbypX2qh5J2mC/BuLKX4fBdJ2rR+qSfJYPmIwsL
jDG0prRBbJiKxjSpSaqEm9uRzXk3War5yYZpgsgxq/WUHwH16Wd3qkdTplc/pCz6sLFEqDuF6Mjp
qYH9GBX4dR4+kJ41k5pqg2ySkxHhJA/vvo/sfn8FMUOCtqi4M2SMtEl8VpgvLa5jaE54iIdVW+P6
LMjjC0S9KxEkGKCbdks0FJbFhiYjpVCKsVmjiYhOY+/fPPF/bcxsUYmD1ptbpvntVSCAF9XN6F0F
jZE4JGLfmsNS7Gd9zKHTrtzIoK/lguA1AuN+Yy1Krg3/5S+CA5bgoPvznC+7B4AzdK22ujPCj1AO
2VFThGN7h2A2bI3auCsP2jyRJUxYEJZmqLs6AJmqbAzwQvBX7O9cW4FF2flBOrtfimSCCRDN5Ae4
ZUgD4VjZJQH0YZQMDCFRJm0/E10r6olDKCoPFfOkBqASPzKQ2emFOgIPo5BAzXyMHX9sVwVYbFb3
ezSJOAzD1bMcZ9TAaHctr8Kz/2RpYt3623tvLJa2+UmCfQi1WCtH7IcJ055oKbsA5cq5QrM2KUsc
CFOywO/61FKl9kmLtXGr2YJdnMibTn6JExYcLK+PWgE+1ZwoIcKnafQu0C6BDtlDj5Q5mMSe5cJE
EFDDS5SlbJo/55KMWrfWBHuxgECIOvfzY56BN5hbOCFv1zxPqjtbWW87icCidFZ9ekqH6U9eVwmT
27DwBUXNccato/dBAVwkZB8fmY/gcG0uFE+qCYn1+LU9L8mSaFoQLu4VoTaiSJ+VJK8/mHLcFIUg
r3iYZvk7aW+bTx44DAWH/70mR+IcQ5sDEmS/mgWHMP8IJZc0pvXjQMVUVYsBXyML6Y1ctd0f7YeH
k21gkHFPRSPovy5J9uOTwa9TjCJWBZJTX1ooa2CwwckbYjF1YWMSz5ESoS9E2wKOxB9yCnp3ugc1
hNAPZ7vVFchwknZgH5IDnoIfNCnO7cdpVi/HLELzcfNkVLTh1z34WNG4vW5MdaHsfqoakfSLsHsa
lLLb+nJbSB1KkLW1DvnL9MIfWaoif4bxC52eWxOBlmvf6eHWhXtMVEycch8FgSPixKs/teYEsCZ1
Qpe9/Rut9ZMEcKv5+bs9cO42OhLyO07dnZ+MvFW3vV+9ct4b5oMbs5D0GHKD+0i1Iwg1JwW1YzVk
hDyP2sUS19QTlfq8LqFUz9WSw4ZNBf3TdmPsHjFZn4r0jgO8gVSF5CTlpHeVSisdh5zn0qjWJ8Hp
5D3SPGWHYpoMbp+xZAZIW+TXvAjBAxXi2JnZACplw3tLADTYo0q+jBFrudnhvOXBnZQjdFB+90p/
WTNJZmcgELRfgdIsqUrHcNNoPeon8TNnk+K+/suNsBBXhzWrY5JkmfLDIrGahHuNaek7Sh81Khg1
Q64Au4FStuLSoH4dMQAqNPOB+WCNegZDDy/Ssvgi2g16KrLB8p00ktChazb27tU1Dy2paMLMMKaa
5K4w31Cre/RigTl/bxbtJutQh1JStgoFNV/F4Fev7zTOwH/RgjfYubQM9E+tyyBWa7/jQXmPgzcg
vLy2djcKo0Yy6DtwiuMxkxL1IdYmb7cj09bQTvQpmbzxmyh4VheVL+wDPzh85Ib5atzeKEvRjMiQ
FhR80//jX5UeUMNOQIv+ZrM0/uobIa+6o7ZcKfvwobvxxaeumK+uDT16rnWf6cgUDIySKq3iUSAx
Piehr/TitxjaWKOM+icsdoWYYw7963kXxcBFIkJ9ZP+JWFLDPej+viLr8K0J8WqH9p7AY6JDPn5k
4TIOMa1qpr0ZZ942w3LLDEhmDVXKLa0YS52eu3FyMy5Lz8EmqQCT1vsDL+FZYlpNgVrQvCQ2kd4Z
Il9aB7AmFuRHVXLb4mKsfz5L+0rR5QA/yQKGIQU/A+Imj+xdXttxMIP3BmVRVDpV7mc+vAjl6aNQ
qr0D6/liTgyAC/gEKYINUOGC/oYpnN6Yjpwoo21Aqk389AQirNfcYd4Vy80EDvx904nZeq5rn8Oq
7R6gESV9rljJibNCOzsQ3kdokbQLvPQNMnjzLioccH8Y6rr3TqECOqBBCp5lPHTv+WMxi6K+60mV
nNfUEsC9XajxuEBACEEagRHDA067v83NhTCf/m4wIYiL7dFFfOGka3Z6JNXz+CdbNmKYK4S3/1Qx
FMNhUX2gdalrXdX1kOXzAPg5T+N0ObvFgqVjGs8t1zC6Qtzrkes8sKA8hg8JlBvvrbY82RB8AfCO
KQrkctW+1zPHi7ATU2UTgBUxJq09466PTj/atPdWwYsn11kgv7u9JAngA8FtXva6fBwgiGoJSPsJ
8dMOLqHFb969AKjXmJvHF6uiwLvgFkei4aqO5AF+9Gk6LgUwdfGj7Wx7TXaVpCEmBGhQYYJ8vsSM
5K3//FGGIFo6cRt56dOH+T5qPqHATICkBB39k1jUqHtxhCbnG9L5B4wszuimD29nhIO1MaBChPFE
+WWW0mEEmxGWJTb15S0dHi1O1vw91OJGeskFLz84qBjFIcyIiUkxUH86sRvbZIN7uesr9hp06665
DHaVN5iwjoqZDPhvd8fNtD04ryh3iGFruFuwb9d67KMgKjIKN1eK6GK0S/FdBhvUdbZ2pLldisyc
bDb+9WY3zqKjILE7NsBNUIvPplJrUoLGJ744Xfuy3K8pfIXbCSL+bySRjQKLbQ6QjBSMHL14lDTj
Ct74LqpjChJta9gnV7e4XNNy/zkF8LHMX/4rm8pukfr+tK+GHjfO2jaYV8NnFCJPA+Fnh5qzWT1P
r80l4OkY2eYJKP6YIENV7p4DgwBDMnkh8oTItFpB3zggNi5R/sQiIQj3IUsEXJxI5Q3mkle3pLLY
Yc7jYppgNDUjdOr/+/jwkJKi68bmoKLMTt8yVsC+WGiEhg2zYSmSiQDwtOUVSj9pwOljx8YsMGd4
s8bDwxj7SkPtnCjVpWfHDnsjhQ3W2HBVfPsRgg/qUFqERvh0PIx6jF7Mx8VdwxAV+BK1yqBU7+0O
dVkGRIbgUhkX9khe9NG8FhZYPYC0TY9mHtchibze18bZooQp/+62I4iwKWVm70ZC3hDACM6ocSlq
O2NqxxaU4Xb19Qjm/tFRRyi0CpSm7agAgokItf6Zci/UlRqkVlWuJvgbuNPBEGOt24FbTcGjIXvC
8a/m2NkH+P5ZzBEOtYU29L3RBfKUGdWOS9UROrNEdLQ8imBXcCzMvQP9PJ+zt/gZqLAjdIG95v7q
AZXI+IzfmLKB2bpYfWytGFmqblLTK1xr1nDlwsUNPBxg8NNEKGCU0H7W7Lcn9SzasHA7P9xrPVXS
INbAJGow5Dp/3lok2kz5u6WPULCPQvUD40zHPC9eqhmB+ky/PczlWQ1kP6n8PZVW4h0f4t+Kn0UQ
J475RC9D6BZv9AJGRpVXakE1/K9m0p0/rDCdyzbx/mvaBvCJtg9pYNiXf9COWq5YdC+nD9/HMOsE
u2uYp0jwR188XjAkeU0+cGMjQZwF/3tyeICfrdmkZXgLBSOwLd3ViGFD2YCNjIlHZFWbVhj4q/k/
isUyG3b3uMwTvaRL8Yu6+MPke5ce7JSBo8O5jfsKbBubsUJHnLL0lU7f4UQuxjgrSkU1swgsWdit
8o7Y9teKhB+jBnKZwPMVPQ8Vy+fP/2BFohVInLG3xDCnRd3Ax3+UVUtTZbFeOjc83xNIsxMB8Bxh
D+6lNuojss/7ZmwovyIkhTC2SVkOiWGZ7pNuDjFSWBKBskPdLFcHDOD14Z6QXRvtYEpxLiWh3+mK
3enkf2S7i0pwM6l4qbw15Lyv7e8e88rngBPEkQNu9lf/yWwUdcVXphV9dU6FeK/s1A6PH0VRypGe
dZzWho8nI7zpFZ7QDii0N9x/n+9TIvuL81EnIioITkTdQubqbcgVOI5QjiI7KKgyUFdDe+owQ326
sFNLKO2o/5Rfo8zxgi85Q329Zt3bztJHGuB9+DJ4GXXPLtjm3iJDPg4jGkKUT+06DyF7qt702W1x
k9O4r6cGFwsMAWRVnoAHyP6NXJOF1818VQ7vuEMC6E7dGrhwHiNkJ7f7oD80q6Z5hUL72a5VnVVc
ud/59H0v5O2O3k9Tyct95zQL9GlzZafqGRLtoflQoU/QOmCoZ2pPIWI+E+faJyqD9BDc6VBG5hzZ
b/VM++W4XoHLzNkH8v8/Pk/CtJwHHujYRmXboC9upyrM/eEaabypZOlUH2KdgFF0WS7LGbb+CHWe
7762PA9l9vB9IN6+rUZVWYf/AtuO2u2Wi8QPXyJYwkLOMGpeTLsKWB/VpZGkgus/qj4kcbAvBHdP
pNZjUyQK5iqCwNuECH8uTPE0lBRZy3npKJEHX37dJ8876PV6uosjo6N8vwXlwI7FPVKQtbfDB3ey
58EBEOge09IUVqdGTe3GSVUiw5qLJfUQoF8OjyWoMm++1BekeKad9o6+fWO4B6daEmW3rGohh+jy
bUjB+iKr4xTe0GCNL7NQV0MgJO+UoFvKiuSi7WU8jlNbSDc1X0aLt77qqBbwpro3K5w9sv1PhqGO
OP69p29P5eAVl09AbqAmYNabparNL03AJhp38VRC+9pYCAztE831oMYdx44wnKiNzt3VHdcq5Ism
Ca4UBLc8D1ktYcI7e7liDT3LeIUu6qKFp4Y3xseSEOjgMBevmkoZd46DZObiehqD7SEYUiF8DsCT
9xyggzR58ZTVwFV2y/8gtrO9daqESuO/NmnK6mWhKli3y8iKCttcFOZSYto30pEFBlfmY7kxnEfA
9lHuLEWjTEIgdluzaxcunohuBV41ACGap/SO2lsIZUPz93yEnCFEco8/z8R2OZLphUIquq/bUFP6
97itsYWLVF/QakiNWInA01er+ruHAWKN0SrhPWWzL1L4JYZS0PMXXSDXQnqWkgPmDHQXJWGivdDx
Si7W90+n87kuoHOTTc9eEuUPQbEFeEWUp+0Jy+Bzav5ijSS/29b9jWT/1bFYOsW0Rnux5w7vReGQ
hUgCAm6mQ7puBBtLcY8K1xuJEPw7Zr7Plze/T91E2rKCJ/gx1MpMsrjeuXuQ8ifE3vbjKwZSjq2q
VxSKAYcTL0crq07QYoTpGp5ZYh427WvIyBz9vZ2/Uvt8eaxZowesMGXUtE/5eCZR1NDm19P9Tkx2
JS68ZGdk6AnvZO1ms0CLtO2ZedoVFn35hdHSeXZ/n9/eYkshrP/wK2qYsB/V0ZDTCSZfuZliPqtS
Yg/wjJmp9zaSBBpsmDt7AunZHDTwiu5IJCAx6YAZlONAHt7A7hwNPV6td3PfsGn+cQs7ZiFT+7H6
NQZ9yvdnezjWtK5NCfJZ3ql62QRuKf8PJoQkHkxjbi5yJer0xDA8abuxZ1tDhxgbt61uWghBGhzw
vEKy1p7z1It5T4UkhrNSH3RqB+Vz0D8z1ur27hN0DWBLyKRMZkkIzGeuWtHSlCfE9yUhkONoYJMP
wcUWPPsPIojLVMyQh3mypBCWzHM0QoGS0N4Gnd0gyvGC6R+zHi68X6kPgQ3uc3T1MW0h6IC6AEWZ
W6R35TYdCg2tNP3zYRiAoSsgKiVdF3wDflvZMLq5xQGq7v1m3cdsCmZYCgjbuk6auWYvPXNPCWZY
Bczq2cTS+KXaECJehuogqwEZX29TDx54vv+8KyuJM0qpIDn9j9ViekkOXiv2xOzY2bzx3G7YguIy
lOvwUI0j3aFKrUtCW6I3ybBFMT1YNU9HBXeZs2OIFgXiDRNhum/DiJUJkQEfjwSkK+xuUxc2JWVu
TxixBlQwYgr+d9VVrqwBtop4JAyFtLi7y3YlhP7ivNdWdLxl4sGgxouE8g/3MjVc3RHhpdthhl+q
ByOMI8ZxCr0KJEtBl4Dtn4ZctO4FbSn927efUsofI7RK+Fw79KP3J9/EdyCw5zlV0ykT5mDBOorO
/uKsr0AyQoQ4V3jvqqxaKOuY1oPP0RxPqmQ/Drc5XX2e7ztIqZBFE7LcsRhFc8uDNdR0eNLoKsMd
CqFCgtEyO1RUkpnhXvc5htQ9l3Ml4uvjtxennyRivEQNppMqZSeqrOAhmQ2vZVp81h1XdnkW1Mct
wVkDzeVrDllN4EC7B7ig9YbN/62QK9dbWqcTdXG3HqLbpENE+/ZrQUoQx0AVETD5ah34AIXa2ctK
kszx+R7DC3i4YPOs2kcew2wj81eIaouhUKEyfkLx0V4jMEhRWfpT5ZRDM+Z3DFa7o6mTyq7z/liI
blcXwL8lTH40Msg3sL23wtc5oGsxI7lsJ8pskbtoGbdjoM2Mc6pLPohX5Js1+eezJUCbs56ocLj4
XIWNRjUWt2mUXjThGJzeWNDZvLNZpfX6JyFXCFixipmsdj3gvoNea8i5xgEw3CF5aghjqw29pCSg
96k6oWKpX+cLGrx0Zn0pzM/jsZE1eWAqBPrCZUsPSSsEe/p0zQoh7yJHCli502A3uEHS1PfC2OxU
+76r9+djGR5mj85dJ5ITFH/pk4uVvpekL7Iyy3UtlCD9lP42qfpdn/Eao7AhEKYU2RF1ugZEYojy
fb1YemSsfDV+aaY+crI/32liwnPlGKgoqAL03RDd3bM+X/DAMIph4z4tmNcoi0detKIP9zfvJlGu
qYeuZi8HHMn4i0HUsoybZcWGiTY7xNcb63y4p/RIVgYa/9LJV9hmE+nS+GkO/bXWfMZ+nTKsEiWw
iDRk6UZG713/z/1ijEjAQPvQTYUjWZxzwt1TbYcr+Kbwk1CQ50UA0xRsqhs4ZOKc7aAyO6DdBQFi
ZPy/fAYCmfAOAsE2YFBN4R85HXSE1x/rvcdCf6NZ02w/8Re50s9a0tSps3fvUcBO6ZK70Uom6sKJ
0hBAhi5WZe+XKzRIiuILHk9hmU7VobHldvP60O5THy3pxc90jI9WHeAhZO9AKr55sf6pjOzVDWX/
gwkzuSyJSrLJl3YrgTqw4JueW3Meo0IHc6sfhgVjYaWxN+XiPShleBSuFAWiOZYixx064zLlafB+
UUXgqp2wZggbP0SnMV9jWzZYM8WrYp6pc6OPzwWJLGjcZRCQJ2DRHGY0EzF9DprncGzBCSMmetMj
LMmgJe3LnC+KLfcfm0JYSxyYvG7HI4lg96vdV8mOeR8OER3SgnXrk1sM55JswpPmk0Pqxl1y47nW
poWUYRhUIe3Jg1VC+hEYMFeWAGDvTI2qFbh23qFOkkvVjEj6aGDuzgOst8wvjbV4QId1tDFE0EQ+
RF97rF6ew12NHkBdPqteqYa5NtZD8hRv07AsmQrPoPbv4t7VqppPtNolZF927yfMk+C7IQgFzmRs
OeDmiGvLXbCbedsGK69WWf5SWsVSadTHOm1ToPfD/uXNR6GIqPDZt5bnJYlcGUWflrIRSqsRuYzW
1tunR4t1LqDjHbgWVHlnHhfQyd6dt+X8BNC2kEQmP6788EQQ5Oq54I0S6RLCm3kmfMMwzNy/nOlr
vL7EGW4czTw5xWlMKpOD2xfbMV8oY87pNjqIak9WPD/ftopdb8aAtTbfU0vp4oRCe35JA450C3tj
J5pvA3ENjYBbML8vIeX8pqM5kXcTqnFpe2YqGpc1qDij83opnYIxuEbJc9UB2awnnoI4ouoVW8cG
00jYYn5El5SyQbow2wyjNgns3QmWA6JDgFq0bpZuJJnqbCvi+3CjgWpRbrN4eFu4Nxszy0CmsSIc
MRByqtl0BtfyJ2VVHLG0zgmxGU31h+3mlRXf7w8uEnkSHPV6lmQ+NQboe1IRspen3j+1zf4l0RW8
DjPhc+wgZut5y3NdFKVCuzHKjTxa8cHxFt5dM/t0eFAZJzTyHqDqwxEdtq6kCPUBE9zwvUl/S5GR
5ZLrwcNfAZWHnNrvnmyWjyehWLe+CtYA6wwbt/UKeQzOumJAagnq+YGZFoO68YMVAiSL2yXTN401
nG/IsKm9343NswMOyspdMZ9HkADNbOh6835aqJrfZATP0adxOkDfmolSxiWK5+LFxsrNRWEJM10A
9G/n/zw6S4hRQitTb1AAExYyj8F51/ogA//ICMbjvFWOMLB23vO4EC22HZ81c4hf4K8v1++YcAfa
eisCa6Gt/6u70VI9oB2h1TFmeAeKQW3+vXYDMNAjMphZ5pidA7Aq1skHN1sTDrfTLc0L4Y34ZDD/
Ryh9a7oaQnnRnZgBjTKFrY3J/QhCsWwXEWA6keIV6UGXdIYwlxdgI/7gKrJN132yts1VPkayWzSu
IVT8GFRW+4xTUwWEFpuezr0XXy43JQc6KVwjfzQQMExSCgkNxrrYULkBKTOUCddisaI/IGQCFZjd
RF+D10o95hHLWamjsZGSF9Cmu1yzY1r0nsfYYP/S5YgUkpEPwt0o5rJ4N/T6VwZo9pKG8Ir7yBb+
RXKbb7Jv/1XOXzQjg8BrlXZkSUcrMNsNLcnANpbfU2HNlQL0x4q6U+bOqfSu+75/uYKudrc2N4z7
UpcjWqL8jsJmMEmEvYECjbJCKA/zyC6HtiwxVdMemt5yUkWNWQ9OA2krrRkaH2fKC2sl/P/buuWj
HOizaCQzY7ViNF4rameOnC3kVWoqfSjwgOdNfgWwbsvG5M+Knw0uAaC7LChppiJcitdxjxg9fHOs
utOOas2ImjcDKTqfBczyb7mrkigjw7ZuRsG3KD3XD6kFE7Ak1a5CyzD/jVltVrLXpN6sH5hEwlGx
gOeLv/rmwzDMRGV+qKiqSG8Yy2OrncbUknOT1m5DK8IZKwdnnhFWPP88aNEvp+UMg/joaPxTyHG7
z78yKIruzOEfHx7Bo5ZmV9sUb7Q7X1vFiE38QhvHJe1POMdeVPoXViNjE+7GLUYbNxa3uOxvc1Wz
uISteR8yOyn8H1XdO+ZeYYvwvInXWER/h+VQ8XYEIn9IW85fyJTlOQHCp64T6sg6MaAHfT8HFFfr
1hFKTUbABoI2CEG6T0oV+gHcJglhAzfQUJzZHB8AOXONuTgcAJ0YjgkG/CgGGBw56ciCg2MEijeh
VFgvXtXd1PFeV3YG/j8o+tV/iB3/dVlYrwzcc1CNc9IBnVFyFC7eAafvWMe8+zPqoSvnHf5D15HT
X0pXYikB3mFRncKplZV2SfTiiLEDqfzGkGKnNnEaPZ+fkiA9HIrl4OqvollR4IM1P9tM14XJplCi
z3lRSD/3RJGUhl9NpW5iuRR21AY/5oTI80keWr1SpUE4AwHUUxsV+aR2Zd7fD9wYMX6uWUTuGzfb
dovwBNLBscRuzBh/fPoWR6GX/wDlfKBy+q0pulKwfJTj+HYbqweL3WvI8EoLijtpTJXVGjfZZ4X0
4kRoJt3zwgwmqH19DQdAFYHsMmw73ymDO/nkcNhR5a3YBrByrL6uH5ZEJQhL3EaTmg/rKWIfYOGq
CG8BZuumGGWJNk+zPSoyP+J4AMW2W0vZKSzs9SoKgHqSbWcp+f3FuIXdxzL+YrH/ASr/hXX4ihXk
V6aeDgD6iMIpBpZfTOnEV4F/JhiUjotDtkphbUmcB9e9UqKYWeC6P0babDCmctvlkB/Py2aqHpgT
Hb6Z6nl8UjSE0ZP9Dj1LKSJi2sAsm7jdAwIxMSgG+o88TLHrPg8MfWbhVNExmGShaC44EJlgW3NV
qH/SO2N8rCtRPH3LNFT2QahuU8hzFKYPkJkGX5jFeS4ED7/XMPv0CO8+8ujeYRrWy85oS4Ix2MPN
ouZgVrYW6AMiFfY8ZWqdg4CWdQznZl+4QSFnJMjb9TZOaDxavwXzS+IYgyMuQXxixIMHvkhnkjJd
VNgsjN0vlmdjDBcQCU+ItZbZ0TxhkyjiR1ELxakQRBJxb4jQEDb6ezGwGYPZyHC+jLHi0PlEj1sI
njRduVVr0VR0oivR5jVib6aloEtoZPsOrQCuLRHwawYBeuou1yimlA60IiqxMSkq7jCaSBdqcB0R
5Zvk2ojy4/rus9a12Eg+Wf3oWSKmZR00r/g2i5dWyBu9ETZJM61vbOqf1WuhX3TXg6/FPS1k8oaw
VbTWYpEwwqPUBVPCQ5uzjQ/VV+6fUFMKQnRVqND8FLa97RaAy+EpYNyuRfKc6IA1BJ0BmgN1dXsg
weisPGYL7v0BTv4x0fKUU1fZ8mdLMlU7YuwY1lEljY62tT1vsaBZNaHzXrcQbBd1WlRD+o9zuYN4
uCskZy8+kKREhbeqgX9UpEYb1HMXVPw0g2QW7KF7yB9iMaKt7wM3gJljXAOCnOpguSWlnU9NHC1s
WeAKAE11KYzjDom8ic/z9G5wau5YAPUeKKaoXyFbCgfEtN8l8kFy+HcNfGFxD+HoxFqGtVdDAH9J
WJvF/ZCPJtc9nUDBwxEXZvb4Nc069u0vUTjP/Ojum0EEBpRzCM/WF08nTintrkNPsIF3SEBiMVG+
eVCgF5j99Wo0YTnhj765L0OUoRFKROg0SdP6VcuA15rkCIBUayVutCF/sUXeOvgh4/52PsgbegDD
F6ytWgPUCVhnCxDAk++3SX9EeEjV9mKrcB9bR5HcfHuc995vlo17/zWygaTPw1JIvC6YfXe5jDLz
YAw7w81rfIS7woVaElX3BlSZahH3h2zUDoS/flVRdXsBvWv9gOaUakyTRtka2MdbBRpKtsXM0KVb
muMCqMlTEturu8SpDfovYCBDXhOLPAw7EHlVzJAmBMw7K+qeNIXO08sBSXb1E+P5icFhR04wl1Af
5C+g0teJmaVOTKD7a/fZb1a2ZtrRaQW5hUaL5EUH6325nHA3daU5LN++ueb3r0MY0cQbaCO54jzs
/iq+Ek3E2I3V5jo6wzaPBGKiF5wUXeefKMXq7DBojNbnZ/klWZZRuKBuhZrkJzOnib6/gBc/I+KS
2CJBsCgl2UQCTNbTPF0gvgkzBFqSu/xiioaSmIbtXiDwU0TcddIpIz0h+LXvSASwXgakhK9U99qI
sNV9dU1T+11lXCog1D+iJJpOOAIC4cJl6SPFEEDAmKdidXtiXhZF6LZNKkxrU9Ep/xjIW27D1qHC
xZMV2adtwKY+bhA5cfb1fCVsevVy4PMoNWYsKJNR4FCL5+Z5MXpi/gXEc2dYaVCYErMo0xTrgcts
qJzgehGZF9fK5mo39f3JPOV8P/hP9Tb4WMfIOih1y+0z8HwVRfqzTF7IfP237h8Mc5JuZy0IpVuV
oSI+ouhcyPKKQmB6X3RJsHlAupA5nT2G+aMnN3GMCp1Gl/Hkt6GX9xCj9Dn9gsH48MYyS3JRtRZD
30aiEgtS3UOg0ecU6b0iVvpexpdBUyfVus+0Hesal1dj47dYtu5x8FADKn+UC2Uo0AtaQadUqF3J
Gh3jRaQJSrkatE+q12w4p/3vtARbEVBDIoKQHA8YZ3Px7mT6p96Dp4euLlFho7cLBGW8VTpdoval
ihgetHQKlLlvhJ3vEoiMOB4NTqef+WaJYafDLH6VSmPHi726/Djk7E4Lm9XacYmq2JDDg7WQtbd+
EHlDdL+HGNFL1RLWNjDzGorzmjK2ACcDyINZD7U6UA54INFMfq2z+jIDpcP7wHld/qLnkXg8dc+N
b73VUq0bsn85OMUZU8une0pI9OiJ4EknYrePNA4qMRxQamM/R9KxNy7uZO9CI6Y9WUgtK2zIU7aH
4KJ4FBhaQKm/+h47sAL31mmST6Td2NKrsyqVxUoCgO6xmJa7G4MoLoHm1X2u7iDd2otUVtxxYjSE
OdvzbJfIVTpYLP2cQhflHUwcNA7fgHDszMqWoeTx+l49HeAQ4q6iRJakDezZtpPrvwrWdVO2JUQh
EBDDV5bP19yaMiOsxuDfFGWtLJBkcdgS9d/U8keHVhvPwLLlKwS5jk09l8G6sUK5r61f4+qG1+M7
/CxmIi+D8lSOWPktEVt4XHkLs90dHu7evFqWVB3kTyJ9DneO8aLB1BhytjggcxznaVvAaTr+Px08
wTb2hl6D0O5aj5uN4vy/Bb7YeHy1e9zv2tNpnlzaNRMfUtBTAhf5oV8uZsn22q0Q9bdhJ7WHQ7h9
cXzgCLKqq8A1Kw2vTe7m00VaQ+5fqfhi48toUSs7odJZm6o9Vyvbh4IgpImYK97FMW7HKVkRJ4Sa
jfBeARMWqlIWELGncAP37rIeMEa3JEZde0+jw0W8o1tnWMkGbnIeFLwHxBbByIFplHdJmVlhicK3
2bIHZnU4Cey7sxAv9oYggqkx0THOx0jspqjGkWXHMrXjQlKsnQZcWrRxykjXuv/oW0UguNaCPogy
J7AaQRw9eB709yfiRmBZwV6+VPGeFUxlvsFp4cVDRHeefHDx8BgjwtddjiJw6J3vptadDZzGDMVg
wV7LIujks8pQ3QRCKnxKq9Zw/bUDc9ozTy11DGk8HnSq5TVqg///IDWVpgLfRS0x6V21opJq0QuU
yz6mbRYdjCB7T21Tdy1R+IDEZVYvSW/avrDJtI3ByV9dlQSFxoVCz1P2fUS+4mVDWQfvVrgvgVp7
H3UeQoQlN6MeE0Yeo5yYrmpFDluBb6m7uGqJjXsq1XkZ6MuFsh0pFLeK8t3BMjRzM1xc5eAGakHH
NAvkWOlDGWxSXuEuD1yAewOPexoAJkWbzeITYFsq+yKoxzroTI5ynrz8n0BYrJMxUcRCSECbJ2dg
koyMUoujJFA/eg/ASvGxDnuDHjtsY8qaJFV4u8VNRJs0bTvF3R+Zu3WEfLThPOwPDzDKn4CbUe1/
jCKAwJEG+L4WdPcFlFxOiQR2S5w+181lbKvUsaft0ZLnxfhB7/T6LcPXnciZtfVCvKnv7gh5jdFy
s+TI0fBbqFeUfIIMEM5dvulPDt9Qz/2YvBuq7Qx43sNhJo3+01Y6q1q5streCjrWW7QL1dDog8d5
/BTvBbYIYxZ1XsNdDp9wcQ8u/yA0GhJ9vXgo08vMgwpqsCyuaANVClwpq4uwtoQryTjVkcF7C1as
OCEGFVN2jI0kOXNjtpIfolOzJEa+3YEX7YGVerFv1X+bbQq0ZTNM/StwjjwVufYjuI6FYLtQwwC5
xdL8xzGcSO9K7v3OEjeI+F+gIP/aX+cMndTUQZlzKT7F/OJ/JtMKgat4RrQsmtbevBDnWmmG+fVX
hPOrO2Rvapl3U0SSV29lphMuNo0hH+jozKIQ/Lvt29uwBUlwnNsJcwkRbeLug7xIHGujvvqMBD4K
waYXvv5u3eS9rKEnaGihZOL9jXx7NDSibx8Oj3iFE5dHy0r4cqpcC4DlZZT9ZI9/m+vyCXpN+kxx
RLg7ZzvraeRUcaawv3mGPg3jZbAYwgmJDJo4jbI7jEiqWxJcappIxLrBsP6QhwwotlLSaPbLIs9z
IQlX0zUH3JsHk7xGbjL+oOrvS+qNMXMcxphIXE49yHBfdMG6JNFbs5uSCwcZV+WzLQEGZ0POdmiM
+J7JStGEHyamoJFdwvrczFh4t+SCjqr5n9Lmg+6t9LV9D5PY+4Dd5wb7aJXl7sVBgXJbrEr1YVqK
E4cRG9B7QW81AKoPANzxvduy6yDqfQ3Ga4WdwFIiW9FnA9Z5gyF0lOPjuC1nN2ExrhlLELO2dtlE
eLJnowti/nxLIXiNL+KjoBMFuGVi9lJJsXYWxVpavbwy1pxzOHXgGf52F48+gUTF15fWnrXrurQD
kyLhlsK8J/d2HJsk73SmdMaE+n7mLalxPVqBA9o2VeJx2sfrBJ+N6HvV/7Sp6iezDvNsHA/Ce7kI
3M/OMlj/BKrVG8seVgYHq+HjF/GByFDWwzXTgF1RDHSrYF7uS/S6MiGOAmiIBrhbDIJioJ00B23N
4jk0Nvl28FGD1xcEOIGB/RdvcrVbRoaJBokc0cRBW1udKVocd4NL1NZ54FglRpbm2wqPh8N1B0Fz
CJTH+IyA7+KAMbwAj4CmUieckG/gGStEvuyyvUAL9lrKRqZ0shnWvEMuJso5CE3BkV++r669dHYs
1YVWDxv9RoTPeVIVv+FKB0fE6Z1zaU/1HEwJWWzN7rlG3YABrQCMo1E70b33LJYwPzH6NvQRuT3/
0dN20j+dak/0oDFZIh3OTvnA2+qy6zfpbJwSZw8GivOaQ0UCS34L+4BwLQuaeQAdyba/br4qipd7
YbBzQKicyDPGxt4BSyytihO0tTlxFGwHBcLpE4CWg9yQuzVI+rNz2wQm7GK8yqIKtrRCVDk9fly9
jyUQhEDIFBrFJAzvgZZmzKGGPM7jjbO8J3PWrh7EpP5r9hNqup6gY3std8ceMPhjIC1AAvJEJWRx
EX4wFckEUzupBKEYgJyRApqupMd0w3SeBxzrbD2y7/5IE+LJ2dwnjrSdMCDoCRi3E2JEIys9akXG
0aWrkN2dePYiPDn9xXRrF56s7VcAia9tqty5zTD8CGsFccqL9hUGM0IXjujg0g/6RKACm7pOI9/Y
zH1e9zkaVAQpBvJt/1OqYa6mNNLJsDEi6X4YUHRECfI0vGqwqJ+HL0IuzBtvENWd696bICMbLvYC
ZGJRUHm/tJgPROqawYIqExdcW43nb26/7YK/uwtlRTfVxDJ8M3YiN2wW0XDrXQHegsFOX1e1vFHy
TpHDIq7xtXIFC0hmMcWf3LAK47GD7nOn8QbZ2wCwO+lwVghI8q8Q962XkHJDn1uvb9dcL2thVAzM
wNxv1HKXYDIswCWVuSqA2l0R7H+9+pYkMHrpanJN7srMjeYG4lmRXkguwjKE49R6peoZCL4+nvG8
eWRQ8atHb7IWR+9JbT7GRgf0xhsXuetPHKfu0Pw0ZtYlCHo7EHOlQFRXIKqAPXhJNHYagFRYZ9a+
Upvbf4VET4M+UecBhCUS5WxPWvaaEskVsQ1x9VfGpP5sudk+PW7fgu+aVuLdBP2Gd1crXr6imMNY
bzB8qswQENnWgU5jc8TZCrPYUskZdR27TBDb63kCcwvI4wRgO0oVJc0uiDMCD7KSccLxZUGGOmw3
I3lRpj1vN2PWWpxYM7OXLZ6fN/NkPpMfwYrR4R5ayEyiIdRCOQdmmVlAcQBUwnzRTAktoXULidP4
nrTRRwcs3qavG+3wcnZtRp4EjOKCvBzbVPJ1dKYj7++dn3HbLLaaNAKacwEwx9WunZsJ88mwyv4H
c7AQd1CEZdD/832m4T3xcfDFhWnrG+V0G9PG0LiJiDnHjPG3XUKlIQnJl8FIJ09vTWZRlA/1hDis
luMYE49SebdZnAeQTeYLfvmuvIQuTdMOdVvy/VVy3rnLX8IdTx09i0LsDbuunPktTPDV9F+eZRjW
eduoblSTFMPadXydZQ2kDbXkzZfS2sex/b7GusQNWoC+GzAnN/dnnswxwgnrA8npldTTOmTZqMPV
od8i1dX840kM/Ymt7LzQf6eadGhSJ0ftGHkurIznBFCjUlToNFZRCNJeqlH3upkF7eFwS/mYUmo5
YO+52dBqNCUSTq4B/Nh0fXsF4W/yL7xHDAwAxXXKvHrv/KQWcWEuyJi+upnZmACXTxrXHavLhHZS
dY6X8KGQWYGTvod7Fq/9tliHiBeZmkNx+jxawXVqQdZ2sDydZcyA8luX8OjIKiEmKvO3Rw9QD1im
KZZ3idcKb97IcmF2F70bR2SkLzgl1WOBGcTXzSMJ6UHTlFmRuEBgFpQFqmsyezr9cNc7ykAKXt85
LrT1C4X6S6NjtTgZFkv5/M6oQdpuKk2iRm6XgbTG2f5uKRsYzBDUmr7TBHqzHBLGfNWNd57QQ4W/
PhXYW5bmi0XpUeS5q21vbe0XZKKVplCdRberU2gjoP3D7OknstMtUAiLXnt9i68G+Orqq8mfipID
O+zzE9FGn6X5wfa8K7BcoPLrLtERbR/73eGVuaYnE2ui/8nR15jbOF3FIi8g7htr/DHOoQOs9EXl
2JoTr0IYuVzdhpYpo+L66O6j/oNoSYbxKbwmaE8KLiQ4jYMnQK/bUQGW+R4N11rwZIV5E6CoVKqX
ADbLHXlmpcqoFPGACeW13UuKrIvshQVTkSqLQS1Ie6Q4Acks1o7+I3rQRQMWe86CjMw3pkGL8AEO
xSUfrf3hQrGYr5gZFfpUKy8VlQJK36kLHV0+rSIfhUV1GfH4kU8QeDLuqfJoL78/2rcVWK15Xn0+
f/1jehSWqxd04RZS0QFMsSjYd5Ju7LQGv3GSZDXdVkTXPbQVxL+Zw1W6kCkYXvf5Yuo1gqoVE4DK
oCGNaW4LLGtMgVlBm2hgl4C9lJmNava4BQmQGTDt4lDP6f9vOpTsNRHl0sU3cTO8wLG2+W0OWj/x
HSIn6ne6drRs8LfcnWWd+4HmE8qZKE0CWiL6ZWoZLwdm9fmBceLFIi9k0OzIOFxwvbnmtkmZjlQS
QSFqiGm0otKzabPaDFAcPlE0d1jDvOTs1VFOC8DWicu4DDuwXrxU1ZOjhgTq9gIP6/7xuraA/P7t
pXbNkWi1VU2DV7NMqYMqG8c1q2kznFe8GAVLTA34Ef3K8IweTcQC6Odzk0+biwfB/xm0b41GTOHw
cTSJk3ee6+iRoh5H/pKIEog+5WDbIHL/DPfCP31RFNIqHg27KSmRvyuTWw67F9Wht6gmV6dLmBMI
8g7/tDa75w3roYashmn0l5XqR/Y9abXoRqMv4CNFyvlYm0SRFt04xjyWt5XZ6p8Sa3nZuo49YJxQ
UqxcK4mEpf2Qt6shP5HaSrc3NXTaoYIwjw1vy1lrzUDpWvNgAI1zOpXFMPB+AFKp3KBtlTmWt9TB
W3pbcMp7x/XLlLQ5tXVMQeDn5NeYYgyYk6lUC4FOFeqc8CZ9CfYnr6IDFsVNy0aeYliP9hb1Xgb4
Y4THuzSRR5QLsSKz0VYokNaIM7FWRSWkWSWzAefxKkbSaSbEe3hLcvuQcNcQKZd9223qOtQLAWVh
CDQHEqBst2oOSJWVmeApzWZy9YgftRX5HalvnYmmBuxKIBt2q4WBhpYemthnQDAh515BpTm/Ons+
SMEuMaWW/yJj4yVCL/ufPHQM1eeIWNmq4PXtkZTK2lrwTx3g09ag5hLI1zUIMYq6LbeVgQn/sKoA
149H7f1FxE1uWDKMGApadVQckqQIRR0FCbYvwWrx44k+yVmCYnQo0ek76150AyFY3xFKfgh8Qb9+
3UBpg6nfn4EYjjHv6EVhKpMGb9UwvsEOjgmZTT93+SQY0eqVfc114pJDiDdFPvZi3oJBz3RaRpME
LP+up+YZ7I9nxKgyIT+bAU6rlYOsixuwO+5fjExO24ouqmKEypWirPLxA1/+ztOiimExABXWEJBd
el+SfTQs5ydX8b2pi6tgMjn64jtZ9AKue80kZm5gjcXqyciLj7L+n4uj8b6DONoqicYdWXm/ASgi
6XtrJM3/ULl9Y20y3KOOxhKwwtIvo+6WhNugi2sRSFQWjA/yuv/ISp1W53XaqxOXi/W0F1SIL7h1
xZJf2GMURe1UKyCuVNEFC5uccYMIUx0H+t0sC2F7JE9oDa80JFY51MyESUIQfgIm5rQBhaUEUuEQ
ruy6rtwi39SYIKPw5mNlnL+hMLPhisxMRqSGjCiYKTjE1pWxXuclb9GWXfIwG912/m07MQ3lk3hh
q79oWj57jBXipZ65jlvJeqc9FCa0J6Rw1g9G6BDB+QbHl2J4k+sAr1D0Lso74ZcAMrI4476DpAQv
jUlzCq4pgJrwAlZfP6bkd5BNVGPoPy3Oe3yWJYVdwixOvKrDfVthhZv1UCHGgiRHXjmcH/6I7ZD/
UVBuRzrCOMrsFSGz6IiTEhtc4qzbvF2fwpt8qpfgJYQyfzSx1VewpBycoOpgiftkxHOzt65e/Cvz
JPDlMLQ2HPYoFWShyqLPgaHnr63c1cyOUmwqG9gR0t4aPB/mD5KS+E/iSNDP+u2TvZzxd/NeIYEL
BwnRyW8pH60NjRAvv59d2t6l+VpfAhFOBRvyv3g2C85MnOkP4dYxaZjJ88btqUOwAnNV0PxYHUtd
BqYVCCATBcfqU2ROPsnnUtO0A5Juh9M295hyq1lCikV1o+5Eiaf4XEXikUKQZ26hvPWzs2gUd5OI
vDvjKogVSLUi/+gYi06dtNYzri/2nMHW2RXrnbK0Mj88VclpzrUx+RCMHYtj2l9si6ByoSDRP+Z0
Dqrypf7KCLOchqsbHJvUyoJSzFKklGdwX1adxOGS1CEqkOYiEUggKc2s0I6gDcO5iaI3wRHfne25
vjdqwJrTc1a4NWvzi/z7wdU+Fg06fhPNUUQ+pB6UyDrekCqeAKXt+im/VYgGh6FEidnDz3GXqu8N
edx/yNVT4TZVf65Qv0+xcmh0iE2vRkQYFwRiES2jIzI0mivW+zrD9DIHAfJD2unAC+wEsxTRRvBh
QG42Ci8lz4QR3RUlZ1WNwFMJwJe1jiBYPMg+y61crl0f/7T97kmJa0fomJz2OMvEy4Cb+oqfJHGC
vJ1h1foC/IAfA8ZUsmkWu5PqolqdYJa9DeewBsrKnB8Hc+4RDpmv7qLGg123qkI/zXYJFm3eBAVU
hljsl1kM0TjECONlG0AaZf8TWQjU5T6JHbKQWgZr2fu521pa6O5T+Y6OWcya98B27sZHGartGsAj
yOgYoIYcI/LnKJq8P2+8XAdtbuYEtGVwW/TQLEXvOpXkd2X1z8zIx4bnq5AOJu2BuA6zvcNx0MhV
/ArHyImIXWIQRWJ2LrcttjN+9pBMszFjue73T3BJzprKm/kVuugrEmLjRM5DIl5oRp9z2FGIY0/Z
L+mnGUNG9mX3AtYX0VRzcFIkriXFUgTTsEeu/a5hAM5F6/Oz832sThE+cEk9RiadgkQqe1Er3wK7
Ks3vDpblWLP4EmqUJQ3WSniSBJc1fVRpeo5IukbR/2fmu8TAlMRMq209hHsEbLOalHmwjkn535Q6
u7gXtOCvKWTk503upZ16gkHAZgC8ub1tOMiJJNldTvBWd5KGMH/ergaECLWn7HEdnZrdbm7Jmtrc
EOAs0IWFD/+LcoerBXRV4JaNqk4cjKc6Zv+UtxIB8kFqIiqs7VyOR8xvCbjWgvLw8HsE85GBB379
KqyCLgKRGHAXUyza24tC4CALKtVZWGGp4rjy/E31S5MZzOL/lsH/8+e5og1SsdLxLYx9kxwsXcBX
s4/7nQ4vMTeF7m994hQhvKZA8ohZDvQ8Ij89Eh9P4x80UEysSrJrsYS01kzUFal6HjN5ct/9ECpn
7AVZ6fngtjUqGv7eRzMnh/7ngiYbqQyAmuzGcIOHmuN7nTwN0djzeY0dq21BLlKeOuffCAL5iVtx
sQTeCRj/zurnpG5ItceFk/y8oqaYAFC2XmPZm2uI9SO2y5klegETU5nkjMSmfqTw0GZpotyqLvoP
hECyaVoPPXJbCs2IxB5AtK0vr0ttswq3fYaU7Pdus3HDzRGOFdQIZ3jxeyPKBbOaW9o9mckV9mP3
sU1i/8a/Rdny6zkF9qryTRp5uainT6VEp3WodHz4AL5ZB8OYPCZitWrzp9U9scEZNiyz3xe9z33S
viI1N+UeDJr3orDr6CeRCo/K+v6mUaePwupgtCUZNk5+jwxi1w2q6FJrl8pYQGLpceBiE8EM4Lxo
HcfH2/GJY0tQ/RC9qP8qFHriGG+iyEQ0oSfzvHdfnBJo8o1XvlXYbT02DniodSyaodMpo2OWZrdH
baXok16a92Ds3ktYFrW0ascLrFNL21X0CDtl9eOT+zyk6GK0O8bdcgp80BxzQE4PY1lUj/YgBc/E
y/pJW3pxS8n+RzU2ovx4EpRN2qMS5CBukMoJJTIdncxb4ZZ2MiKGr1ylo7bcv4AdP31TxGnOODc2
cbAZ8qj4w49XafziuVKVm2dx5c4lq48EsDdypb+DGRQfBoOHfOMdBgwK4SsI3ANwERQ44wfXdiJf
0S/FudTSRT2tFdjqpeY8uyOsRQvfaTZIN3pQOpOXk3iKym7qvcy/jFjlqR1DIB2SDqibFMkSwCso
716LYIR5Hjl09jwOVERea38rESfeRGHwKRl+KporLY68sMRTbm9wu+BTt0TJdc/I6FQkJVOPExzs
9el8rhOAkh/3qIv40pkairs5w2hg6oaH1HpPKMhGWvUy6mKr+ff4eOc36cngRPomVjoI3/Fgq31m
zpeiPTSemNemvops+r5b0lVjsbMkW2WAWenfR2Qq6okKPdIAnI9Vzhs1L2yjKqBdBmeejN1nQ5XC
L2wM930lpo4TzFMyD0z2QlMxNGyNeB5CWPO3oyczLg7Ftn0nQ1SlRqkELETUoGeC5pdyKXSGEMlL
AJjVsY7qqcbk6if6chnkDS8xNROxuy+r0gvg3sOFTEAY1AlutJv8ZN+VccLEvgVLD3s/Hq5Ti2hh
d8EKVE0YczgA9oaOW3gG4cZIgt57lnXULoQrSzRcS8UNgD23wa3LDM3Yd9JOrMVDBnvRW+wg8Y4b
uu4GnnTgGSk8SNTuj39unLb51q9KtKUOGFN7ACwXgH6nppHXHVft6l0RLE3RsTfgdgwlRm/0gYp4
NnE3KUDZBpFxxBr0sWgJuwbkrmZ+L9Q+u/qpj2nFToOk3I5B9T9/GZDa3/4R3rT8+y2fGY+6ztA7
/59tOQkZzthtXhHEhB6FJUA7cDYiiyrqMig31tbQms3rz6Z1tgpu80/bPxFYPkwDTRfcAv9VCUMY
aYnz92tePoAftL03iPOzOVBZFm8xWUu415kRTBRUygQv/3dHRbGnC7I4WtfYGCjIM5TMqi6jHmSe
ulTj+sbibd6s2PlICoUGdBREzfNFNPHSqFGVmTN9ppdfDOQyafog7hXyv+CtN0yrQp6I5dEIklHY
rbGGGe1plWQYdX/7DQ8J0Jmt1kTCF2mrewRWspbBnDInE0UUeALijik5dlReht28ongvgX7UpSeE
fWx0KH9ZWTRGfwudVHlgUeFGQweRK7/A6x0RH2j2RyBkcBsmjvie8kYfyYyLf7fmL0PTyacDWJuA
//k20BFHqtoc0QwXHV9NdqrfZaPSfmm+e6n7CV7IcLrvK8L7GkMQ3FpyalW7IkUSxR6DrfQaw79A
Tk5ymVBldcUq4b95bvbg5oJ8z3MzSusWXeoPYnGrSaVlP7GR8radIwRNp//vDrMKSBQn9B53y57N
3qqguxKEX5RPeh9g3SwcaZfs9ibZHNLiS/lCwvysdLuxsGPnrJDAOCtE8+U3d8dHV+eybFxNilBV
KWPXjV1iKCLLIFwAcvvFZ3V73uLKz2uuUHIO8LQjRor3OzBUNc9rzOjmLeLh4MK2r3Rqv3rmHWLy
bLWbrJA/At+CyLTvrzepdlKXMPgZKpgLTocf0UElnokOhVG1EkKWcAq3ltFxNtxouDjda3Hc6wYT
5wTpI2qbCG1qk8Zl/hyU70GpQB+9D5r6OfX4hJczYoe75ZJChi9x60vbY3z+4qMCJOGZjWf9QcGU
3Q0ZYDt9ZxjoXhmNfitm6nE091gE2C0NAKze8sgpickzaPSxPt/Le1bsM0RqBV96nOJ6gfFmmfCn
6qpeagRbrrELhUp3k2ps3YPW7UVjA0/GHrJOBfsetYc3Q5Y/vUKfLIw7bR6cA8ziGQ+KvNtUrmAR
lZ5YdVS//6AHnDTZ+enp0g3DhirIE0ue+jIaNnIRv/we7Dybi76G9lrpbDMP6SllrQxYUrWpJ1PF
F1Gp9SI5HR7L3qQ9jP64UhCx4ah/P6Nc6pXvmCxpthifWGjoqo9mULrkmDjgVfCm1EYGP3I5r96y
PZYDEyq6vCmzWGDUU3C7VkoFq+If43POxMnoQzuT7dqyz5MlTMcbFCtGM7Zn4Rh9bICuajvhtTj9
WBF8+XbeJT15uWUK0LX5HZTFrGK2nqJi47yNwy29dSP5ApeLE5uJlP+HjQ0ytGlk43OoKLk+H8MA
VmYjM8jAk5wukLEMJ8Ed+z8oz9x7mEgSZlRnRHeZoHr2FM9v3UhcE8JIxX0hDL5U9GkB2Vg38sbC
SbaYlpgHXUS23L22J3kVWfkWsqyXReEj/6CSuNKSIdrYh7niLP7USjHts1wKeIS9DrkNMdBmSTJM
b0cJkUbx40U7EFHvVQIaZ8qq1IN13++iEW5doYu9jqc0nl9C/y87TV62CKFsOVuDOqBYhN5/G4jq
NkIt7EDGOWEEiRB64yIs4jMEmZ46XpX2WtXHB0ul/q1s1qoYH7o+3biCw/c0Y18YJPuC5JfsfSPH
H/0yuyGFMWLP15/HJ6sqcC7SO6vRHRzb7sreVWBSoteefYpT9/mMkupAizzLmM+20eQ7PGYwjxkP
mSxeFKcg3uGM12h3NIEvvxmnlRJYEwpoLe93IViPQ3QHM4kjaxFMx3LM51l+3KEEQDsjSYWqOBil
kMp4s8QCB8sjuGIAiXBFWC8pMmcfB/hW5oErMNLtlScFzIStHOMlhafzGtQ/0JAZ4WqAChry1wco
dJmf8rPYEg5z+K/BJKSK0lv7vGd1Z8eGS7k8NIm4obLDLLpeoiKQ/Dhcx+VgG1NRSnnvELLCvX+S
yrrPfuljLKWWr7Uetj4bVksy3YDgPMQtYLqkZVyBQ0sKQaM0sraAbfgXEnLZvULiYdTOHTz4dNrq
ChFdthZS6XRmYnMKkjOZRbKjcl4Eowh2/6QwevDl4qPDNgLbk97nCx/HnOdoaVUVSdJk3nPJ/p2I
abkguHAbd1mAMiuyJSoUJZWwpbkbuKpP2fqqGPHfE4alpj+OFBpMDQzQ0Qe4wgATd9hzscmCnBEk
Kj8USl5S+vbh6qw3PVyKOg37Rnfcg+Hw3WnRtYVJEmxxOKUGOTpLZDfSFHFZMtLkARDRF5caLyG4
vSpasDiSuiAw1PERGcah86tZxTyUD8TkTtbRMv0zfJ0DgR0KmMS2/lCLMttLtT+utXDVnhUHji4J
qCvGDiRKzCYooPMY7DqVsa+SqrInV6euKnj1JzQ+AL8fhBhq7oe2JaZ1wdZ2pZMEbKelfj9aAvPK
/WWtoryq1psay5Iz5KbdXqCtTPKNuG/g+X2GPNVSTJrJ8PfeAmSR/fei761ZGrorAOXdsbJYDD+F
bI4CV1asF3WobNzIKP+ZKt7dmA71K6XVe2vqS5RU6WMmFc0ONoP5elFVz2kZH3wsfQkJvDu+bSCo
CtwtWgJJVc/XXGTAw42VzCWw0U4J69SaqGJEtYI9DWO0H0KrAp+xqmGC+wqH5xFpUacv8f46cnZJ
cQb06Fljb7wr88t8UrTdfnDW4+bmQjlzl57YKI8rsxru0Bx43BAmqxphCO7If7tOz3a3a0PGu6hp
gQxl/SuTqCAdekGos3AaFjgcx9U1iSmTqtPqfDYutMRpnRaz/KmruLCg4Fla7lpc7fDro6gwBW4n
HffH4JrnNfheA3RgphG/wRRnAJaY19DzNd9lL1dptRH4Lo53sxrP1vT9I9dr6AJL3Wq/p/ry2maH
y9CWSk1rKT5Q3JG0zdyiiVE/Pp7kNkTQ8a2SLWFl0N/Nqq6NDrdoh4qAmkH+mNUN6V386NiMH0PC
2Rm5oqMyerKQHyd2W23I2zIfjL78iQTtzdnEpnLQLsbCqlGPz2R1FoDu89PT9g5gAnJ/miwRrmHr
JipkzG+Qz8dgi+GQdrbUu8rl7iZtGIFk7udossLSA14/dk2vn26/ixB/6ZYw92eQHqSPr1C5oFku
k4KGFibwpaweagVxZ+Eeseo281RbSQM1WV4JufNDTHf1kfBk+6HyCC6+IErClPGrWjrO+4xfftyg
giqlrtFKkUxuJ1Zs491Xi6BncblmQBpe0I7Pj4BrrRgQgoYAv/5Yfw8A5N4m7ApL8o1IImioCFiP
Ff56AcCiQnOTSGXlrJkBnTAMbPQ628DQta9msTF0e5NW4ROuyerJ+VbBYM9XeqtFIeuPAlNg8qA/
ptN6b29ttWUMRborbwx6VhRz/wpzGBVzBXluD9IclSmXEawRkJeoF5rAT+2upMAPlMCNQEfPG+c5
gUTRzTELW1D/3yY9KTuA0MJ9ox1eC2xbdiz3Iz7vTmOlt5grKZwNLRJmmCy2dmJ4Drh7Uf7Iz7OF
0i4TXNLOsbt2au+5NwrCN3y2oWKqkQzL7E9Ubh2nWLI1o4rS6nZWDE5PKehZcUNX4NvlZqs6YaGl
/DPvyLlQPsZ3EiWhJuamIPCkQ+DM3qTQXcWJTVtcmE8rKBJ401OSEr0TW7YfbGjFha1HYZujLsAf
6tRR1UlWRV6ThrCq+kiEwTBVhhHmGX7W3gIvrvx6G+dH5v5PJK9funcnwL7GHBmKC8m0BZtzcTay
dax/jT87RtYG6dBkGaqLi3/tkYNP8xzKkq83okTTl5xuP5XblJCosBlDi2SorUQkrHny2Lx2c66H
IbSsnN7mM4WDwwgqfsTvTcmXAq/HYZ1vBfssTnf72rhyAEEwS5Qph/yJhcujNjZj5N2hBKighIw+
7Eq/mYDV2DNjDBwD/Z2ta+cLSIHlb9hiYG2NTIH76KJDKcaUmtFXm00V2fvkbhTBipvgYFI+Y/Cs
crhTpGce+BDTuTaHlMosE1NJ2Ojxvvo+yz2uuSbfq89/A2/A2QDoWbChDurgpUwG4Sr+nvY0oiMb
l5JLdHSDFAY+Inl+E1pK99fmqNHF6dJGQWRSE9TtP38Tvf2uwN7GnrST562mMPs3VqXgjv4yMa0Y
g/RNNlpNIugs8LXvDKAOwwpjy6rLvBFkp3aLdmWsV9EZeYpUEijfY20rngqxLYDTGp0iKwu7tp0G
Miec+bw+iQQu6Oy4uy7s0+1eqgIIztKFiOBM2tTnKm3TSywWxfMIN4xI1+UvtiSHTqxfChZpA9co
b58FpjyI1DhSrQJcpWKtIYsKccrla3FdOZ9ZwqE6718HqtdWRYVyoW9TPeuV39VySvU+lkut/qar
51A94nF9OW/HlITMwOaj4qDoOP2/MFHspvQH9tuia0DIAZsl5kuCqyESA3Y/kxMc0piowSffySdx
kx1s0mPZDKq+OGLT1Fg+evQht6jHCF9wmucjuG46GlR/UiE1IhwewMn30Y6HCY5zhLPno5BtEsxE
pAPP3I0nzApsFuU73Edvr5+Y80+CT11OkSSMtHBsLnbcA2sk/cEkJ40aRR4IlcRhFr2uV/5hs+ZZ
ibXLuxE6MXqAg099eM1YG2stLdz+B5QnJiZCMq1zAOa1gXTSRwUhiO6PMhit76+e/xPujJLjnvql
+vSRjWe/QuA/KQZoJaeuseNjeoMXv6TyHiuMnlodhrV+fq1vDWJJN+YDP8hQZ5QW+3yqkim/y0b/
dnNklety2NRPqa5inX4YFHNisAUXfnHyl1gB+WP+uKZAoEdPSHFwyEGja08ZRKR4MVXjKicunaUh
rCCgvSji3NOEWvX+bCfWE3Io0kW7WKWJ8jJBWnS8YZrMQu8toecMrrNJMgKCyKMZG3DRnuwo96vS
ZPK6RUSfjvwsMb7CqCeJT8DeketpU5tZy60c0rNq3wL36V6V1R+2edT4TeUODypnpniAooFEdLRv
rbxzyLXBr+imsLYv14s2+y5F2dufdpICKFiUyUdVi9hVu/iUPAE6QpD1KfUBZ++e7FrLMdAkCNN5
jFZyGjVH6QdinXj5lrghrfH4Ksj2VIV6flV74+uiLM2AxaQ9CVhLLEvWSmHIAij6k2CYBgMHGChY
5QEYqfsv87F/70c3KLV3wY/kbyeUiFIOvAi4g1W1n2boS3YXymPLsRpNo4vM1udR+Hk9SGiQRhyH
aboF6dgu+6p/Hc+kLjLJznIJ+KerE6DFQpyoma4tJODWx0twwTcVp9kzSJQYQxcFbtik/NWk4K0o
rCc1TVUH56v7TpmH22Bu0fPRS3LySwFiC/R2wsIkGa8CxbA8BjWycC3EdVepUyQhGC6UvCc1s5Vs
qKHvuxRhiFI1LcgNzj7McaTF4JOQUD7vtvD39zq2Fkdsq36sQzOswzSc5xiWcsFhVEeOtiAsSNsC
0Nkcsnan+5QwC1HtjItuGRkMWmtDeXgT5k9NIHC2Rx6zfrVVa3erD2+1KHuDupPEPq8VyOtQAIk/
4yqhIw0KNKan39nyoDlnxSvdug/dyCDBFNpWkBRdLqm6ErX7PveTbUaT7mlrpJUkopKNSKvoXDUA
oYdqo3qxNAUwLw4dNEVnbRyKGTtDT+pGwHzZkzhduvBqfALYwgyRD6WYhb9AmTlY8COS+XmQCei8
fPWJLWeY0cSAp+x5hAyvZTcSzwKZP1Qu0OSV6Pfokf58rh3J108x1IuDqKw0nsx71JMZkTPVkaL1
G9Wx1Am7lYx2+BZhJwzoekeui+Taw6jnbnDWCmDuqNDcsl+M0x+YXk6P+P8uRiIA7Qa5JS7oXA07
AXzeRgJbfw2DorDDcY5fHfnifInkwLn8YKCWOoCYaKMCc+nbQSQAjJ1apmuBhE9MkLnU32I/FOxL
SxhQfMSSU+cZLbo5Jp+0Ead2GeCIHIRADtFlNmCViqiDUWSaKuhK6r/hVC8EoUgls9wf56DsXU5I
K/suOLhr2Zn70NVGW0VAdq57oU5UBsSA4zoIVjMgYNGRFtR/yMtP0Eo/66Oa527/P6qUVj+yT5IE
i9vOkH5vifg94VcAW7JN8Vfmsym8e6/e1JYUJUP271PovKnzmxhqbOMN4a37gpak5aG/fDwl5L5a
jNeM9K1DuhnSNEee2viBqyetQwJ+9fg3vpDh+bixpPQgKpOiUGUKCGcDbKxWDtEKiuCFpPQv5pRb
mr1xCPaXzrmou4WnvjkrvH/EaJJPIfN71Rmz/TeYQhr75n/JZW99fnIQu3ebfS3YR9hg+Thht4nG
oA94YHRnVM6wrXgBZqi1dfIlKZ8cupSvgxP2A1BBSepiFnsJpdxvJI3vo9Rp3BoX/OmHQbXw4wnw
pi+RcDiW9+eS1GHHoT9ukJ/UkjmyoZhEE/rmIzu37bSkvm6ADCPE+3IQNjZWeQN4OllKVP2UDxFt
8VmmSIvY6QO+cQFusABmL89IR0YmZjGfYEeMCknZf7HCUDohtlxU9UVN014JaaqQHxsx81wBRN/K
f6YXLZrxRq0APX7moi7i7nbQiBR4QQgDSWY5DW1WZNz1t5miTY52KOeAf84iV+NRsSO1LWI61/md
WfWGKmufA0uPzSW4XieWKI6OyKOq/W1Lib1ErLXEwsme73HbimpK6tfpiLZNcTYgHlCJoFEjn07T
FPArMudzdttfoZXoo3/mMtDbMbRXNapBlPS7ezJ5mJh8Bwt/HuovjZRUlw5HnuljtygGTPTSbnN1
t/O06qmhyhoCi7KCFIE10VmYsgctSp5Wb0RLxCedGvNwqIZ5zpgvS5YPQLFlpuDDHzNNgubNuiF1
mQz6+Ouo0A89hQnbYCowHnTGOIzJB8efGc1L8Rm8yD+ndNHWhMcs1aq1FG/KFPbIt2w6+fM6trQx
nzNAS8wR02HbV5DGKUntsFLhHoEVB51rgDO0BPi+LPCqyN65Ttj8TI8gh3m4JlnQOoiBzJZIoitM
ylsl2ITq5CiJJak9kUft892cEEW/I+PTWoom86o0FTLpgRzj/DD7xweSSr1dhB4SjWv0Pi4tGbq9
cgFLQ9Bohx/dQcvD78mzGLJXE/Uq9xL6eqWK639Nt6fQT1x/eMlLtZ3WJhrcvvjyfWhz6f4n4uc/
x0/PfPLHnEIJKw/piXv7cyv/MiVsUq9RhVCYEOBDoLxuR650x8ndxxejCUdbqvCs7n+NzYeE043D
zV5RwW7+qA8LQQgBkflxFs7orMUbDsgbhzvlq6stfhcrrbOKvpnJn5df2TNKxDBqP82ciKnoo6yw
0GWC6X70/AyXW+NlAYQiDeZFqYVwleJhOAdLH93C2xdkdgFEFfUffQ3uQzG0ooLGZjAK9UHj9rOM
QxFS8rp7lthWVOCyFE7wkfU2nafY1pCuTZq3Ssx47KngHt0uUsMPplxDdZfEWWks05e0AjI40X83
GQxIrWSiW1bGzBYv7NZ7LJBSS+ftp68cp93/x2NUasFVChaZtH7NKeG+/dOc7KKRMC32TQevv3vJ
sTpEmo0Pb3B4wHvDkh+YHxe8N4MKngsFYzr82K4ZWvqBpDT1Z8f38viNcZwxl6Od0bnAAUdAMErF
OIu/TdOctyN1Ah0OEg4VxsmIi06nBLU3C/53K8le3nevk5RkgVKAK65cxk9C5SWFs+Y90xddoEnb
D8bEHieRTQ7rkTWQMmib4ShTgMrFL6v/fDtAHAyjxKC+i8OmxmisgYBVGQmxD2AKqJMhOClLYA6W
LUgrqO3+f4Nfin934jQe/Ei1JcCmQ8/tB1sA1jZFbJY/wHh7YT3AuxWBbqZoEoJHrG5nZjpms0Jt
Gbalj5UyJ5UrnsrjCgL//z6xxmYhmzDbr6PuhoJgWVzUu0xvXfjYb7NoKqfDXBFBM3MSw5TlwRJy
VZuwV2wAH486/NwMmrDMGX7V0xa1WNYG41Zy+Oq4K4M40srJQMcgYbvbIKehL11fOPVlir79Xo1m
kW9xCc2xs+y01y5Odw/kmCSdEYB/7Zt4cMj9URysFTBk4Fg8b0wbuvJhKkeOgED7Tiop4zrlxFty
FkRpUXw6bq4RkfADkYS4Z8WGOjrLpgLcle4a9PsyqUpTjNq5zQ+s3PH/qm8qPm6W/f695gNkXBJp
JqLHQfdnKVoBe5a2kbcFPOKsHy6lcgvMRLjsT9TDZFlrfUQMGh3FDsiqMXfu211kgtcTva+ttAu6
Fa/SnMN1QWB/vC4BQgTw6vX/tjwaVmmH6VpKI+kiiW1fuOcn9HOhNu7rjkE1Xi2rI5Fd8v/l6nN/
0/D2wGd0z8yb1AUDB4CL/e2BxUBTVAmhoO1K44vckiTUmRNI9RRDQ12FRg+DdhgV9GtiD5f2MA9K
siFGKqY7iw87wktsRuVaFN88h/Uau6ZuOzp6rUxqyXPeadtDYH1ShXGjcGjmcNs9ZAqzuFsMtKiq
hPEto2WHxR0DhzR0LBWR7pmeNoCpRQkGJKhHhR8E1Hyw6OzQXGVpLKJX3n9gxuTyld61w3Rp2x2u
lCsj4vwfYfsTNiJTw/MiO+zG2PR2LH+cobbAaTLKe0b/Nf16cq9SdevxhlGkZqsx3+HzqQdjaDYY
y0Wt+dUSGLXmQSdyKi1DCsD9ePG6r0i+Av28JodBZoU7NKBJ3E2SSvLLPBdnNsusoMMsq9SwSsVU
RRd5SiWEZrFd4+GUTb8hldojUbwkvLzYagxlgVhHBsJMSVKmLBmUM6adS63P+l17nziiaiiHLUt9
zdTgQkE/s5/BY0kohD82dWoateJjlAAT0krTsVpITf4ehTHdSMvvA7F+kDJ/rFf/ZWGBzabepT3q
kX9vgx22Atl9Hzt665MTNHAOEB6bpTdmyBlXg0VB2yyLBxY4+8YNnyCYZijKrTasgTL3th6emBlH
rsnOfGtEjaL/UPvyPQXSM2M510gEfLArl96VCGRpse9L0fPLjxx5hQnuJZLlLuE9+dZhG0lcKNaT
ru8P5RllpCoQX8VB70ZKXJoQXEAmqpCMVSQZN3hpjuUQAGMd/ArqT+gzedm4Ob7b700CWFeUDBhD
g/pIy4PlnMEpQoYXZsyCJ5WC0yomD9NxYPuHsDhTJ2+sfTOUYWMiYkh4DWiJL8VhVvuaisVVDkEn
oA5D69rBFMd3gUQwUvmaSbImK8s+204VEc2QR3TmJaeV7R4iycvsH2SuccBR38DP3UdFdSd41UHE
k8tXgMpL4EUy+epeFGGVOPvd66vkT65OUXjZKE6qmxMi1miIVRKMTKTpmN4VKo1zejyzW0ZUbMfB
RJNCyZpoAfm4YF+Us/t04ZRDv0fT5dijCe+SGl/uXck0MvKFwOyWu+45xbv0f6XKpywsw0J3OLqP
MrZ8FwRjye0PBRMy8yWXfSDPcfAlluBT4qnnhS2ryZ3/HYm63nzSaLIfR3Tlh2RgKKDPbUNnQaZQ
CgOVcSYDrIeHQEJCqybjm0LRgz1cNjGU9WTl+M+Lz2mEoMwCjNXiDTbE32HbYiElp0I+z931Pf4b
eVYWXhCsNYGo9/M2EBqVpqrIbQL2XvvsKACSq94k//9Hs33zkPJMH6jNuy7tonaYg6ZtkEktXe74
49NCoL1JdGF4rVo1hQBY7rp+6cqEJ6F38caEdHqFv3RP/W4umhnQ9wnpHj97QOW1NeS1BWdN3HWK
QubCcJlI0TCguSTplM9SjeG0NhUSvr3kS/MnhMgl+P2lOuxNyfbp2oVFfBMfFictb3vLzL2ovOHe
l6nY5cEJWVf02zOxetfpTt94zc/nM8pVWA0ydEzobPEnyaydO1ZPKpeoo50eUCAbyIauRlW1cvxw
hdJ3IbF+i01IS6Kk2PdPYAGSAgDdlprmVSN52YQ28uTFvR3CUtrvShnQj5NTO2LTadVAhXFfudm1
QS28jhbi78ByQ1FfomRwP++doUCADQRhDdLjvXd+mcNXG1H5xlZstg55vDyAIQxDvdxqXWDWgNdn
jmJtvvPRUkpKaVbccGRsGAnRAxnzXubGkpCSLk4Z+GkyOeaj4iMHBMrBLkfugPsQ4I5kLAyv7eAD
EPeyEBMlJ7Ff+J7L07p77Ag8dZEUsKm6uiptXOXAKlzUuGsmDtWnUE0wO1Yr7pFDPVhFOqAdr5dl
STBWUuej3aOvElubthbEeBFnHCMBIFFINkc18H4quqJyUegHQ0Dc5my5w+010G4/AUbrd87fyMNj
Ov7LY7oT1kn+LP7J41HtbqMWnh8V2w/4p6lkiMnDfjBxcGqHnlXHyV1bFTV1pvvKijHxRnssbHC5
ptwBE47nk1f3wcMTC5hmT/CzDuu6A09viuElzZL1TkVt/Em4y/+K+DeFa5C0/1PJupzak0/ZpdCB
9pRkFOJV5sJkLoK5mJFd0E1cG3IGL4TBjxQIFAjupVQzSS9PMMHfcrtE5jdYPCOLrrw74O+UEGz3
BJ5nCiqTej2t357CZu9r+VqGXQJeyyRDfHXksZvyJ85klk0eTE4x1uLD4D0kmoyVbn/wrXzUX0OW
z2tAtvh5hoamBSPDd059Wa+LK434hgVnGyfIzSaSXN4DZG4iBvt61rkBoLzeoYGhPh8nFt+oTbvp
U5TzqA4nKTO0vI36ODzFpnZEKr0Eia1DUMCM329+V/KDG8HihTjFOFoWJpy2/FWPCKZNs8rTzlby
Y59ZZRHux1E2ZsVcBxz8nKnQ5bhB2lWntNUKM7ZuSVEHuQdA54uJOu3wSThgNHGEemh1IAE9pV/k
oWv0TuBT8jdB68l5V047k9LzEcc2hy55EB2pVFsgqEYA5r26kT3YFHbvOynd7XF3hC/xbpWRPvze
6airhYnxZcHZwkA4TOsM3L+c0O5GdWaHxlgByewmZxluaL0wTcFja2lpUO5SjkyoQwTRxiCHrWf4
7d7o70mh+HYVknGZVLqomTXFIDSkBn39Pv1tqpjcDYXSkk84kjQVfhgY5c0Fu8OnfqEAXUI6Cggy
oHCaqe1ZpbuqgH3r9SJWKQPeF3O3wh2DLWNNlcihiUnQaSguv+Ya/l9QEIs1CngVdd8lIl1yejtv
nGqCFaHpgR2BKT8suYW9ABO6vQvE/XClWFyzRXWyg5xCJzTnl/8+jaajhMfqV81AJqp9J2ZlZJnm
ELiYn91uAXX2ZKFJEN7MmZD+d8ij0g9+Bn/7X30IfBrC5YdflWMybWSh0E+2CD0VkDsU307vRXEF
ha4gurNaowawRSadUjLxM4Y910H8iS8QK3PSjN7rcimcQH7Y7MgbLokqxY8oULfmlHAgActdeRIR
EtLrwqyKUd+MbDH3PoGKlFzRPlFVAXoE924Nj2sNmgIEQX7aNQH8ifizr9ehzbOpIujtZ/9JFJk7
kMUUQITD796KVvG0FBQV3NlqUtzd8fodneD94PwPndTEa9WDJshTkFqvp2h4Zah8gYK9I+3sznoT
PaETslsfpZzZlRknwpIzR/UwS8JP3Jrw9GJidHBxoj+5tJ/qPL6wUxcD4RyUp4ZOafSxXgLShqGf
eUWUmGYGJAk4ciKEMBe1b109O+3KAlmg1kMCTw3OcmdnAi3lL3Bf95/mg0yKVpJ+dr67POgk9lZe
jB85664BENeDnTLBwF2MdMzAnBM5vpybfHHffIqE9p7uA4ekGX/mcsBCfXwepvNljDci7wdJIdwd
vy+c5/wQ3AmQsRZ1vDZCNVhBjgDOo+MrPFKOVZr46TJ+kJEqt7x3Mx9HgUqqmNV8b5mrle3kqDUB
8FpeK4rrXo+0V/UtMSTGMCn6c6a75pQyG1cuHXY/Qbj3XA0zxjQDWXXV7+K1bIBtBoGf6qBlcSoH
eRhAgrIy6fRnlO641AIfq8r41/IMnH3KIVb0k5Rs539quoJyVMOgeP3UJjR5rdAZfkoBPL/NVf/A
X3bd7qFTZVa0M9MN5PXms8XWj2Q+HWNrPAt6RXyQ8iXojC0oU+wrzFvbLwRVou3UP5yUACE6nZkJ
xs/XD/RsGBQ54CxfavoPnQrin/Tt8JQzB7cZSxPA78qVQ1nDq8601nQysuwosiE3wSOHRK6fwIvC
iuIISPbu5kePcWwNGwvJ/aryPZIUdC6FZFs3kViCUR5Hi2nsE9oF/O/IRs/tTyZ2B7eCL1MjCb2T
3TAopGGbSX6BmOPkpIzYrL+kX2toIWXvVW30XUEQIrNxpiKUqFRoXmYn9WhNkhixob6iISbYl5RC
4SDPfV/b91KYYs1uMrpxHn7UHsj+sJTkZe/QvsF9PDoMYj5xxFE1f2OyYmEsdN2506KLOQJEM96a
XFbhmiLKcebRHygSfhwvf1Rd9MDHhQEpHY8AATo7lhuzrCduiGLjlednApi+g6A9LkkqpOr9ylId
Y6TMf0PyPwxVS7RTkXiHM77E9QqFgDn4xTebLJCOz7ZU5w66kS+T6zLpQG8likMC9WlSU3uFwvuw
tPN7hr+z2PeoxiEirD1rB194VrDPU/9gDP+5bCEyIynNKJFZFsfbGPpxgU5J9sEr1YXlrz5R+y7V
HbJCwf2M5XUpwP4cydDQjjRiSK0pQ0Uva/aCYHJaKiQ0yhWFc8hqqUJ9Dv9BHMLcmtZ2hk+fV0SF
6rgWTJII1usxm7vBBu2TPXvgIzCSgnQr+x0JLshS0Jae/RHz4ZC0JrNkgzuFkoTXp0R8hrRwVkUd
OcffIAYudP/tkUpIJH2Zs5G0UW5QmQj4JJIeNmjAtfb9DfkVwr18DnHlkFBS88/1ZAqPT58K2uEC
CtGzAcPVLB6q4q65bBLSSyo7tEDW6C9nln6Sr6q1sCK1G9Hb27VlPTZxVWu6QInsX5oNtaRU9Bl6
oMYUQ+397/lToxNCnVE7sj4IdU5V0MKMA/yabBAgXOk90covqUEKl6N4VAIjiIoyjM0X64tLvHcJ
kvTUKlTvo8qqeN62lSgOoVrSi1EnHtpuebK64d55DJXvZAbT29UId/8QraOHq/d8BAi7KiPvEWyo
B2hiDcfldxynD6eBqq42una+tq1ZVmNJktwnIbSA78sYAyTTTIZNDYGTPWNZe0sGGZIcCLRj+7IF
PxK/rr4bWhtl+X4Jr5bfokatmXJuhqxnYkTsNDCOLQxW3hhQMmOv1zLEFMLyYMKBxUSlK9sig17e
hkZWfu/fIN6Jydu9DRhVxjama1GXQG9pro+mmOLtU91GfzExFf6oyNSnGIXAbDZiUhx355uFErAB
0L93NCBJeZaLjnFfQRQFE47aLLDJFgX6XBitjTwsbTb+SFYW4J5OFKorbWo/ot9PWiieh8OV82Oo
6rckNoVdTsPjMPMkZQAZP9gqx58+gqHkCzTJSTvgx9KB+s3+1tqPstWudCWRb6lhssyMr3p8gvv1
lWKsetFbTgYfjJTk2xPcp3SSMx6+mCxzfjaP2TQtRkHR0nbfY2WXypivyuhTZy2f1lKAFtIBUcqJ
+oi9qrxLr9u2oS99JLNdH8DQP4IyGne3Cgv1rf8+iiG8aSmr46g1Vnu4VvUrMsI3pc7vEz1pbM1m
ZPs6vOlv4/mOzov0QgKFOQ/3b57ZkPp+dqv4sUQSoFML+cDoFU/EEyH3m2tYUGMXF39dJlRObA4u
98xalGuMcTJ9Qom7y1yvWfggCjNgk8qD647cigUVc2PsPVb0K9s7IxdWRpc9zBp7kt8qp8IPxZol
J8XlbKkIpLjBGD3V8dsMIo3TS4XQ6dmpRYrJA4lf8/A0R5nLPCRbfCEEYEFku8jiUVuy/qwy9tht
UxuWibX8/80DWGfLSTFA155X2K4jyH73d4RsTdFgS8TuYNnHudj0xJbmLnnpzeCS3bVFMMCEnAsX
w7O26MGTEqhnn7wTohB1w5E9G3xQY/uM2VxYbeElaoI0HFFYes/deRgQCE4XMxTFqMzvZB0BNX2d
kwP3f9LdtbpkXnFStZOoQRBHfsJEF8IJEKjUMc4WGyhechhsXy6FMaDtTR8EVwBDa4UkqCWnd252
Fd8Guo0Sc+WRLQpOs0c4w9aiegADum6SpJKb/QM+7EAL2kUCiZTtzuQYbHcgsZVvhjugZ3Iw5zxD
9KBm/6geuovHokze1EgxCxRED9z0b9J8wLO8OcWAKwO+QPYsT5weZyG3J/STqVE+/nn/aiERwqes
PyUGwBq7b+UXIMbb3QcP7JwVajkYLgeKvOFZ45S/NkRe2MvGhHbipg/BSPtVDxqfkdipto3ohzuc
xyuvBUn4pSBnHghvHFINpkC+w9GBM+rzC8JOUU7Y6WV/iS1B1HAOCWbfAY/1Vb75DNn7/U7rMQv4
BcfEqg36MRX+czT2bOEQKOzKtOWkCLVLODcWxJiWoJnSYjOfG3Zu7tcV4HvhYTQ60mCFcVhXHZl0
vTZ+ltqbAdmyeBN2QBnt4AFQCnpqFaEqE2K/JZWztlxVv5VF/sMEC8n1J3OX69Ytfiq/6RWJhdXK
Q9l8EQ9uW5VWQV1CvLu7/9cwHegFNANMy1U+B6uYDWRTRJW87amSBkUcFtobmmv08gGEs4dcZCIj
ukvig+H0sfdfeMUxGQXPXzclftIZJ4AVsF7C938QXPxGDxERrgjlTM+FT2rmBA1wgCFs0HgDpChR
vFrHLZmuvnHAGz6BhtzuGVzppuEAVBD6UitSKRU8ljlIVpv6Vk46M56zv9N9VW7IWYzGZ5rT67k4
vv2mddjbLVugcOlO816L8aB3UCF/r1ed0WfJ7VLCxurGzxWT5kZ9uqySPDEDHr2q3H4CFV6Hv+IP
BE5tiEvFn0/tNoMUZhmekxaCOcZpERt7vJQEZ22zHcz1A+ulCj4XnP38hlBbGZwRJpliGFuRITOa
vIxrA5UCmFdOJGYpZM/59BdQzJ6h6Glguzn/GSSekhhziqJhOyZ/N42neP4Za3FxCHHLSJ9dbEqb
wEEAXetnBcKSNNv2uRRQr+bAZA++/hzpWMua3KefX3zfj/B7s8jxCQXNOqC3KYqsk7ORjLS39vpd
Sj71YO8ycbBhS0ue4pvgrdpEQ7WwVRnL0qUwf05HFJ3fr0FIAh8cv9e3M2f35DKzasi5UdlXjqdN
m2WifHMeIAi41guxp7gBhxZKmUMXZmVVVN8Ym3HkUuNXEGICV7w3dbd8Y65o+jHZcb5BkMSA1n15
VPggGX9+JWMcRx22J2JjblASCw7F8Qr5n8aXG5WeWZcRkXDiORWDXNOcx4PtWWblbUdaVvTlSvwg
rp9hl+G/r2j8db6jJ8miUsilQr72vQzWVZXTaZE/nzFGAXoR1tBnfR9P3aZyplnMO5oG2px5en/M
FtiwoHJoiW1hFsWkvQZgqSPR6M+22Ca4rIw9cqi0nwltVXqR9tGQVUmlauDZbagsC63qklsOQauR
maELWa+8MJ0ys4AF5FrqWs8L67S89RO/tO3ACsGb5XXjTSHEwgMsdoWGL5972ln+x87PUPtCDwuf
ElSIHESbibqMK8TuDFjBOog0nAlZnQ4YxpJyinP5C128czTTc27jBNo5+mk/aQlDePcaTUW5ssXB
gPEv8So6gK4oKVhSn09UNjLicWOPYHDmb7VA0bBID5SHs5LcXPNM/b0WUXn/DK0MoxKFreq+bLOo
GbQuMjgv2iA5GoS8Wv4ud9nEnpou121gK9RKY3euR9Zg1ljYKR5VHmccGIF4fIRrY2aqsRSFBfPl
3OygnX1pHe6aFpgA4RwtdvevNCVsZnPk52220l3EbSeJwYYrRKIL9NAKhji4HoghoTvMUWkdp26Y
BwZUA8oZQGESw/nkELc/jow87JOjfOpME5AMTtF6cJhwMQuEkGSkZx5q0CU49uL8o/K84uWrLwvH
PDJqxRNfUcxkrRyV2y9qgL8hXex3Pjy6CIASsA9nw5pNAbAMdRwUpeENUNGo4YRka7GOjEQoqha/
KyGuaJCe6we+N5vw7nnYrj5Wat41NeNhOLltzCHdvqXA8Z8OOKffTiSU1DkT0BmVvoAFpW3v+eev
izaqiPZVlTpZWg6fVVs+QLU/nepb3i0b5xt9FbkMDN4aStmhkeN/hl30zN31h+OmMKOS8WDOl7+A
G1/6i+jLa+jrxK8lTUWR8BQNjb7vlwWQ0s/O28SAFcru1k50Ac2PVXpMQtNGxxWyBhkvY1A4I+10
N568e6zYnWqf6NJ0f23YPnetMxRrfXqIsOjZH1OqS+D12vg6VlEI9dEt+y0Qvb/q9x4/xSo2fPsR
Ah13wRqtRw6tq86Ok/WXZfYPODTBjP7ldibrLtwThS8WVUSHTLbCc78/HRvUJjh0+3taNX1Egu6q
xdYhGWJeIIDG2j73WhSQtmc9AkdsYGird9IMaT6Odyp62tuEwaWczI6KsgZPTeUuhowZm9W5KEcD
Pf0YtXGSVcsGekPkJP/X3hWNvflTpFK4pZlZN2nS0Z5UedBs0iiE24ineAwKBZbx1g98C5dqxoSn
TFx40xQijkIaGfl8REL2iNcKzm47A3+egRjOTCzRoFQIkE7lnCIuGo+0X2lVtVaAlvsFk3PVkLP6
w46ASGUUWE8rHMQ1QUv5+rG1qdtVBQ/6sV1xFch3q9/KAsoUXlM2bgxAyCwGIYr/nE/GySB3D7Ua
RkXafhqzq4cz7E62tygLML/+fSXwc8sL20n+0QBAEoIpHQgJtk1lfORAZ2kbTmLnCMJIuzZOpFcM
dJUihAJ4MeHeKGgbjzUr0+03xYbUj4pGvqhL+Iz64mlO3DNAL6RGYcmonfdBhuPKv4Y+DwyVFzCl
3k5BWEWodwvC0UbqjMYMC85PiL3LQom+Jy6e7Jo8Pc00K4sawVv7gGtP0KmaUfcJ7u1QKuUxAwph
gVIY6UkOk8gjKrSkeumYoUZAQswcsuZaArAZZUtcTV7k0RmdTQ/gJ8DkeKuTan0bxplvMsdnpDZO
y+OfXF+ks04K+cB5t/0m7iO0EKXGAtDqFHPGlBmkzD9eiR36RC37MQFREA1bxy61vv25LpLVywbo
V6/enDEj6LmKunqzfZNEm/HQxTMJCfP2L7Km57JkUa72fnSwtbFeph43PVm512OZQ4Rq+HaDxQQ8
oDaSrqRHGILzIO7liXW6NbJEDAjLbFJ4yMv5EQave1E+BbM7k361lkUglYx+vRPKnXvAnQCVwpID
f3lpBVqSEtf/guMLUodl/ZW7v4tO9uTA1x8nMsrz90ZYdGx0vFw/X6ZSceRR5rHROnLoAwaZjssq
gByfqSDFJpZKDMdD45ctnDJiyldl9RIgbiPts6jEmWilS1k2BeaLlLZ4w3PHftGGqgXmxYKtrzLm
8+LKPLkNdYAvLdRMQI1EbQhWHC77ssM7h9/FD5MoP1qA+Bdadbto54U7uH0kSbnEBkGM0wL7B8rf
XqlQpYwZDIrWKhzFCaDl2GL9YH1M1b/ZhWdy3sMMQTTeOHRL2/Wjmr+9W94x6qMLgJdRdZGNIYvr
7VUT5UvfrGAS0sIgIqXIAjEgYShGycgH7TM/cVdeUCpGuEBE2M8QgnHJvu/S4OpEHUCfR5/Pe8pf
v/CAACjz5nBk+WDeHCK6a0sx8Oj05IuxCR7iX3KHiwutB2v1ph2BeDhDuXvq7jqd0uFevOlmAUji
gd1dXvFw56l49WCtkUVntR3+WX8SFXj6kmahm1kdPmQnrAEzm3rZXCRAvYnjfFYlU2b9iMbL3vBs
VLOeKU/yNr3y4ZjUeKU0bVAfNN3d+55SeTpojYKG3LKD6W9rgi4ZUjlgzG5g+USeJxc1l5S2u06o
ZSYsiYZPWARsqxF8KtsTkQ2kQIF3Qn24l9zU/HHUSgKCkfiZO5OiBpOYGWSqBCZkohZuWZMY709u
kGiI7uYbbmZW7BcjJ3guE1j4MYkEflOVdTBwz4BXQ7cFPN0KTMaMy4z5091DiYwq43AcatoyEeHx
M2GOk1B4EMXTyGhtP1jHAiv2X6c2llmvSECMnfGwdSsreaW2v4wMllQIaK3Nv7meynpY3g2FOmOz
HUGJBAj45LZ336hii17mO4Q4rK3SJBqOfWHeGZLAU25iEIl4eGVYzOq7TbVuwVeG+wRiJtKDfj3D
pq8qtkx9Zqv5UxXCqMySyWNHibIlBoqUTbZAOyygSCxwVobIxGQzEQ8edQF85YHrsQzaJscrDvle
thMtxYznNrnH4ztmpYfK+PZRMAc+8vYwDx81/8oMlDtgwXcjGnk48kT1t87DIZCIzBaBAvENrWGm
Qij2Zc/rkMObVsa6dWP1V2ywM1BHnOsMJw3RmwVZSeRfIZ+syZ96KATyZFu8sAV2xPH+HH+VyHPp
Z+uXY0YxJWI5sAlH2dX+FFUX4kj+GgpXw5ZJ2kGgbJXOhOfIxN6IvT5qvPDtidVIqo3lqI2Fq0p/
sF5fht19RmHkbU9CTvDbrqauJqiGh+PhVylC6qyPMc2LuzrAKYEm4nrVgioFm7l6rwgNQxpaZVd3
Fxj3ZF32JY1vY24ZXjz/65xcwimpeivMmylcuYj48lFqck7t3XoRLnN/Jd3IUicsV6IL/Ciw1k+F
7SGiWEl7Ffzz+/ko8gu/Y3RBTT/nzEa56/J0K2Xtq+/MYiX06dKgvtj9xHOVSwu+I0dK+/Ij+gGU
piI/rRrVqWlplLTGum4Aa3xq7jWZ2HHwt8jl8Wv1M4JtVsenJya/T6UJb5v4OZCK1UJSzLzwBMcy
KtY3lAUFjyhseyB1lVHSeAEHg7AkgFwBxjWDS6I0gVupllrehHq3QRQ2HX/rt/UdaO804xc9M/sf
dDq2HqvRyWm/aDr1ts8l+CZ7jlzYiegQ2oWoGSUsNOvks4XVldSycFxCemuwGePWVSWXz7zakkGE
8tjYF7zTNlB70pD2FIgQo4VIpvw0Fb549ouK/VDBqxamVaWXOj7RgsFkENZVxp6LH2/LDiNyTWHQ
FoeiAXeM6MWEJg7i+mAhLGz55fMNlP4zFwR9VolUkxti2OYRqtkNHkXgw0IE9sOorhu6eyaJCj6z
uIWo2TyBQoP6m9QdqIAXNP3fdJ1U2TgVgUNOT1wuZJ51kuWp61SigAyz7AT6sdyCkst8vyyNCjgK
kg2eSvBqJbTilaq9j4sjQxhfC+Qn5erUsxNGTnP0oytL31kYSIeVADtkboHgtszCRBcVzrOmAE+x
njyDR9pnQHxkh48S8owXNmYtSRk+jATTq1L4vUPorn+DYdKZuhi9eO8gnVj8trbO/8gJxjP5ZhPS
ROH8HoTLrJOgBrKrYIYQhmA2HWH+CeiLVxgBf+vCdgdlnGNBy1Yy+p0MkZJI6Ow8clcZmdKChR8J
TEqOKGqjkVSyNL5qIj0Me1U+2Oxovoayg7q31PSW3+aRAGDU4VvHURq0O6BxlR++cCOt84PWdQmv
x1tULEpmFWOlXqT7Wu0eeG00HF2HOKdNZvtMmPFALeMnoJMgvCiciIS1Nfsqq5ZynLlgY+3u9AjP
jab1EGxg8xnFY/yA96q8U1IMPCfnvU//y0wvH6DOxFvnKt2Sm6QeMlbxugkr5T8x1Cw9tGq6jTzb
QzWmjLdO/n2BRUHVPrSysmzwRU8How1fxMwg0m9X18o0//tQZ6wrBJqDpUFHLOuzovpKSOavrFm7
xfyyPujRsIx6AinhK9NeWWYgKb5NB+xv25nSf75+NmyUqABrhfb6ZZf6CbVfl+6JsyC+d5tRZyQb
3Y3Pa2rZeEbxVh1aKUaI8awcJl2O7KOKs07etzbXfj7k+FPZCIYwg4xaHSNlO7OKZRZvUbwCuRxa
JMWDbVOsoU5IGnA6JbnngoRJ0cLgrxqxKtiXge/CmMnZa84ksVKg1GxEOBji2XMsTbLNChBIvU8X
kutKGG+CD9WmU9TvO7rLVH0I12Tz+n6x++qe71HpMO/x5dYJdjnOcAyIhOoA7NnKEKhzQz8lTBkY
tiZjpVqCqwCkzJsqLQNbyKusx9V7OKgD8gqlAfPggIZIgQ43WCm3i4dlVoP2lCEm4T+LKOi5s62M
K7aJ5HFaI/GoIhehvkrZKokF3cLAA5zE75fGTxu4g/5MDDbXnCZQygz3A4Y2T6kxCxBstEQcp5B+
zFyPnGBFPfHPbwDghJLb3x68kWlhxXELvrmRSbGTSJuy6DV9AJ9DbQBYwQRoLdjtnj1UDXDp6fuv
LhteENAe+cCaAD6pHwqnpQ5rb4m9YO9TxHFLqA1j22o57aJSBoGw/NImMO22djg5zAlxwkiwXayv
oY8DP/Jd1/6TJ7IeQhOD+cRWfIiXbzHU2IpFXIbjOLU5cTHm6spp9xXhOEzkACiW9xfIOQN7ZFr6
tO30c49PLLtovX+fjd5xqeza7ycLl0eIy/Ki2fWIBQy0+qEp66rj7a3lAjbvkqpJRx6QYLK+HmxI
xZbqNasYDrSD3jgofIwnwk6PZK6hSpHRAjT334m+G86Ohaj5h8+ka0zVJxVV1Y9Ju6wBe5yioQu9
4+m5sYIY+nZFOOIRLIfIAACD5Z/CZiO9Ac1QQI0yvVf1bwAlD/0om5IWXa60l9nGfvko7AQibHR3
2DjAsO5sBi+pJ2p4D55Wjc2saEgGaEMUQWcQmEn7rTK9NDEmK94wdFHeeAjQkRdKpWAWtYDUWO8p
yo+RqbhxKe4rx/XQA4XgVCySCHG8OAWewy7xLkOGBtVc/1OYUpdvR9lTx3Zoor0F98tTpaIXtVc6
P+W/dBOS3/yTa2PhBvJptnukv7mT/AkzRvzh9Gnh9Nb4B+q9WuoLnYt4bsGPZAgj38c8JmfUQ0ql
qtdvwUYhqF/sIwwnUO1jR7H+Ty1JE1fkCGNc0zNbNa2OncjKgGO6jB1HKqucQva5zCmN1t21ger6
PmbvqoxsPjTFh8RJI4LXrfX++CtKkZpQ/QIzXvKzzdNxh6tUE/im3M95fnonFP+TjOfoPVzVvNfo
5p9KtJA+/+p94vwVKFOv7xy63QovgNJUqA9Kr8Nn/+XjQZIUH80BtdZct0dW58+m31CeHJGSaex1
3WaNwXDrRnMrV1pO+q/ss88L7V+tGqNyLqpq1MOj7/v0myRaJ+n8rgzYWhMVdtSijfNYQSh72nWP
fzgk6013jdy/F6e2Z5TQn6s7jjlkchec1hdW2EAFWtI5jS0US8bEGDcWRmwjt/skIMFjuOAkQSdz
ZzZUTnKPZ1uVzdSW9PXPldwuWr7kNO8jJbTrrLB4yDHdmQ8jQESXPkYRihNa91O317W2IgQa+zow
W43epmheDkP27a5oAuSwfWv8+zmauiFLjNB3iBiP+QSXMpUngrOMSuObTsCRK7QQXRw+lYDToLw7
64EzD0tE+EjWMwR7Lac5+b2P2NUrc07InBhE+3mOk84KQrUBaMu5NCK4k9UDQPa5f2gHQvIpYAwv
Zzlb3Lxb8rsHkVozQy27XS6TM2ZEeaVJdYjWtTQcxmbvR+InQ8EY555A/i2ZxZ4Ilz3eQ5DAGFLR
ul7LQzYFKuhAcw2obOexQY+uDvS5r0tgTXNVCPoTal/SeKMPpf1m4i09sMqhJlIPX6UX19fqUg7U
o+Cy5hOUHZd7WkOieJEvX42M7QgdTnjaXInhykX9igulgNlWs6O4ZeemP3WJiq+ZmOTixLlVe8dr
xDX7B17AtKHrs1mP1aXxzL2L1pNvTxLuwvme72XYrD8o7wb9skaogxmcnp5T5mt+9PeAVqHan4He
YEEZfdMn05PHfrQzP34i/FevAEG41BgCApnVtf8gqRjIPkjrGC/peoDWRTtQRQbsc5RYPuyqNGDh
4B5KqmVExsTX8jP+NY7kUYu/3Z1R/mo8YxrOnarMxZh9vnUv8Q9QoBPazPD61m0WS2oCWhZ4QCvb
BcOMgYvWWyOcWtJ7IbqbwId5ZeIOO8gGG+9xnLhskQS5H1cXfvj9IeXgeTd5ISiiI0Ox2SgHmzTs
V+juF6w2/pzeKrsl8m6RonWYdLy6cSnNgahrH8Q0VP6KrJnnwv0aA64LiqJ9QVd8Yu+GNitM1UeN
rBzWQ36G9Zjg6fM2eOpt/aITwWugWJwcoTcz1MRt8iOHCxmdjL1yQe6k5n5Obr8eI4PS8x5owmNE
3edLlqXhGZ7ANkgPS4i67jb9Mxwkrh0R8aVnOJYlDXZnFL407qVpvuHgRDK0Wmcs90IdGoB1Ekir
7vRcEw9VoTMMY+l3pndYL7SGgHB5S+IIyoN3zCiyTWfFFlFmmKRo1LDrTnfybMU3yss0Gq+8LwHI
x3LbY9fucYrl2gH18q/u6UA+Ky8edO7Tna+r1xxATeYO+eUtVSjTfVDL1wcIU+qJMoyYXk7HfFmD
JjnqeIdH0y38BqImqV/ugIWkN4EtwVXr+yWwBwPdZLPzPbiG005ykIq/9VCTmoPqf2sP8V2M5KBF
1GIk5JPU6Hya8ltprkxAc5Md7JVK9OpnkmsBPUZCgh0i/33wfRe4c83toDTGItbPBIYA/6Hl0HjB
0gy2ssIpk+P3oFlsfEtSvzkjgtHdHbTbXrKordTyqMNINQJzDm0sL9vJQixHyvxX6O9xe7lEHnxH
K1a6G4tOvMcIi+ksUhRdUV754koeyPMAII9RWuXTF9iLcuasuKT/eiGwknpFXK8jxFW414MfDt9n
Bt+82oXG/Eb0tUfGpde1QjcWpDjNV8w3G4o2mVWscOdV+qS6jnoXJrqKQ5+9S/F9mn9Sxuy4DDRf
bkByJW7PT8CaT0Es2Z70+MYNPmEonQabu05laVEw3KW4yzRS4dCeQvemWvJQg2w+C0EwIcjZVW+s
Y2CbxeCWxHQINGdL/EgQ2SYwYvr8AslOnW6r82gFFoUKft6i+EdDdzfYxpIXErUFRP81vvFVGrlT
PYKtoPgheRcuRO/zGPqu1Np7/nVUilwBOYpvkyYZX0D/+b8bflBvUnVm2gJf3ArVMKJuR+7shdZm
30XBGuS6VCBkNV6W6RS/NGC7dPLz+u84qZ26AQL5HAd/utvG8Ys873C5xIWCUd+BbQk2fgjO7VZW
EJxM3Wqxg/uBVwE1AS00ulGz331lTDW/cw2fhOOCT6CJUEK5XNnEhpxiWRRP6oG0kB6F8KuaXFtm
XX2nRBrhs7OWwi9WAC6VOY09xyn/t10+shvJZxy5nokDHHfp1TZdxeDFDd2p/Y7jiQBH5NiP73nK
PS5AK5/24DstE9ixpZzvxTL8XgAm4pv9kBE+1niEval+5jWO+W5+WU5WZJyoSlcNT6GN9kgeQW3f
dnWKTBDnK+pkGRv2cXTV00fhTcWz5PMXIgim2zO7xJxaGm3ylcc7xQ8IwiQmTjyt6bIc3HcLbE8r
hL+yBYZ09Lcuy6oC3p2Ij45fugiToxqWN2MEkJpn+PkqZkm7Sjo14cT2XkkDN2udKgYNQBAOfBLH
GDuYUenQt8yZCPrB49EsgDmR23N4Suty7xIpbhTyGF6VosQytVXm9De/XrZ/PCf/Nd98mvwNPLi3
bWcALqfXslYlXbchCLiGjjuH3GNuew4NadK0wYOkVOYfGMLPUqzJNg6NNCy6qkI/5flLvmADWkTa
GVRRJMMWg59iw7v2EKwxf7tkdb12DkhczB7CvnC7FhQ2SZxSrSb10VYoiBw7lwDlE0F4kxGUnbby
ltSmZF9TJvs+TUwDm7W4jo7M1TICtvD4mVkbKEM6LvFQGKEaHDQpC8l+jFX+Ob9CVrTEM9fYLjh1
Rlp5tRkOt7H2Qaf0CI2MvAZmO7KdnuIMKMBnVezidjDXRpL0eWqnwqPlUH5Lfb/km0o5kVYntct7
Z5yBGTMypflVv5rqDDEmPza4FJPtLVvVH/dHxUaBTv1YD4G60x/Es4G0XhB0PhFKlQN8imkcGhM5
b17sN4uYGEMtb+7JUdoA61kmll4A7y5Zs/kyt9RK6X+H8Y4eD54mwbmTEsGMWXZTQnld4n6Pm5O/
HJm30p1rbE3L4pbMJGwJxCNSR5qnwXoqOkjdMlRzjlmg9zzif+k03rsNJDB3fOA3+RyJFRodZ+db
GjQAv8MMLADDP/10Rr58rxi6RLFohC7vikFSIlA6kGMveRDzY9l0iwQVdXlG+kmbE54Po2moBCZU
EBnce+jE/0Smz5rys/Upeq0W1ZzyDwsFgiUz1sqRl1XlIZmZM/aSjNpOgaAgaauZTbsntt8rTsnn
6o+q0KBPxNaGomwsdF/yQ8/o7ITecHDuLS3GB2DCNmJjXG4puQaDlcu0QwXUICSr6CNm/Pw7af4k
fqukZh+PywZuIm2tEyktcrjBvYfW8TibY+/XQw55DSWaUm29DLLKosWAJ9xo0cH1/7FXDfP2w0nr
vYx0zoRXxRXRqrTOGaDGtOeJ2UIo+nzUnmSI1LWD/LFnlq/n/msa+uPXVKKOvGN42+czu6kQiq6t
vcoSUgb/6ajbCrxpiCPd/mQDk1e5imI3zmjZLwaFeJMzEe3ioMGNICY8McVANyo2WRs4TnNT5YR7
1Gfnv3OCO3QaYCiAwJ6ozWiDf2A7WUrHXRSvFW7IBJwz5CjqYbg4KoZ1UO5hcQ99oS/gc6h1+Qvf
JSSExb/8hwNiYa84t8/knIgIhOfb76GTfadDob3qhxSQ4b6ujjVjUxF8W8/RrYTWPQ+g4JlsrDDr
GDUp9IlS2GNaDsCvdE1aCB3SYdwSLUQF0xx5Oim1T1cOXUDnQFVpfbS7Ux1t7Zan2CXA0ol0rMzl
GdWbaz2wm8w5ZC+Ny7d75xrhVRwRqx1ePHP80p9Dxc7TgP/cjcRkcQ/ddwrxoIGTipJwIxrs1x3D
7hmIq3KkP2tZtpi7e9lLRQBht63k4gaiqSJsx6wBjsI+HpkOXXtpPzzvYcRlhXJb36tLqEIh6/MZ
8P9eJW15YvpO5XuEL9K9bIHf/s7adp9r0wkuhdhhSnS3fWFQcyxh31T28bW1m39tG3ceOiHVJ8MU
XAHjLCxY0nErxB8VKn8nnBXqD0HrfoCCCqeHSD4z587pRg1WPjEI3b1rkUsMQ7Fz6O12EQ76GstS
34R9H4PVMyX0UjbDlB4iMvRAyjkZVyfGq/tEWYrPyoPPS2geRh7zEy/pT8d3gWqe7C2WAotkDXal
mExWy9DWF5ofSVmbfK/rTBPBJjhHpcZH7c7ohDB2hqpW9g77tG9LGbJDf5tGW/6nwYd2m3PVtU/b
LZ8QsB9YelWZcvKTJBOSKJnGeVEiOrn77seqKVsDU+V7Fgr1nyV26QiXQn+z8NmOs45ob0ofBAaT
7U9Yxwv+aZHuhe/UOkAt9TTdyzw8kwdvs8bnwqLAwOQb0SegZqyalcWZxqqiIqucfUgGOeFBvbqe
7oTLE/8x09oRE3O8wo+jFwNv5o+RE5KWCIuCVsXZsIc7OCP5FA+z5qOXjhnEI2b22F05vMy8ZTrn
y08wxyUw8WEWtWw06EefkZbtnl5MF8RPxVQ8h3yBQ3uwnT0oDJZRm74X908LlgpSBDBaK5Lb/XCE
cxfAQKaFXi6rwCIVjkFD26p3OK3YvCOzaHEqK9aTbYimHsnREWF5QtY0Bf2C7gNFpqYtveV60HGA
C772ZSWzVFaMwh6Q9jttYU1VHkCVQkDy6NsLI+ugmVceXk1qxN/jMvNSuLC1ShbElDaFWbx10aYk
M/9m0I5NTRySdvy9Lwk4mu1MbKaPqISwofFQTkfKjX/xSjfePmFBq2R0hoI/rmxwGFCJgXf5Yw2k
G5GhjkARNykUjyqQ0OgDi3KZWe7Ab+ULxXHemvBydllDWmogHOg6B8O6ahO5PwJk3Qof972wR2SP
xmSdV6O6Q0YTe1FgNDamT04+tBRHgLJ+KwnvI+C8wpGgZ/fnFcKpO5HRbRj5RAMjrhjuZCSVicw4
plNYyWzT5rnvAM4r25qd8PJaY5sPKBPiltxxVfVIIbX/dvgNlyxlZ7CQAMjpuKOheYpKHk0tQBNk
tlO0as4dqvF8MeVe1LqUMhUo7plsy/UveybBrp//7WXP6/j5gl5bSZCj+UsVk4upG7VQ1gdRFjHj
Oq+tyU4CmFrenF2owUnXSxinXAm1Fx7X2kvtQYs3tMRYHl9HhG3nIaoHREgGOjNgKdbdNG9PHN/C
RaxeL5x7O+9k5Lke0d7FX50WSZRGZcL8bKdMnT/M9RXoAR9Ci+mPke4/hGwvcUw/4txHdUUzV34/
3DnkD5AuBB7rFEq2HzI2rUpXFGa/ll+lXD5CohXTN97kkiXYvRmD9omePcbR1azklEL7NJs7zjYj
VaNKOfWIw8ZTvA9mzuiDT6XIAIfyLUn+sn9bUYULFbtKOdNlSvqRi6Bo56/nTm89HzGJCkUtXvqS
2r/UkM0y+9uFStfFKky/AkDyCqvzpHodSTmb3Yf2cQyyLs0wtHnUDLL5hoX5q7O32ZHcordrnhYg
UU4nl90sIKULwt7xNIJ6K7T4evX7B54PlzqwwQKA+8+zeI5XoYAjrmqo1VhsyhT5YgHkw8/wrVyu
TDjTWLEFBdkoclJzHiXRTB1MQyTWmhYSwlG2AP06QFU4NOLR60/77cnkJX3oZt+fq1kh7BiZh/Cp
UpNxmZp1zG7vVrfb+YXZ/AfOJysuAUeb67M2EsUGHfM4m3nov+6gIGiEwR4WTTweJhBCM40lXOcL
/ppJSeYGL8QK3ritZtH1GZhR53fU7kfWGx9Q3FdQMDkUyidU/d6JNNYlYJY4JyqXFRmCwZ5g88gy
dbKiXzq6wKD4r7zEbHXXL44uvrjdDadwljUTW+M1P0I+FnGOcfkESDq9nyBDPkZJSUkyid6ij+R2
NrHQvbf6iEGClu91ktkNiqPmzDrcw/6pGGmLAd5uqdxfFveaq1toFLxnkq4UACNGxTDPrdVqYfkX
nMZ9wGsyYFtvdRxl8UquT6YKHW7ikRvL8tzG9rGw5/AmKIPVDBX/lcc2/Wj5qNd43FpRFOcIPIIH
rAFSJ2oXsnY+tjjRUum7JknAXXPx0oN1oPmraRqeYuIZg6z/DR8HyMAoLb6dby2P7pdYYwP5izUi
AEn4F5yDWY/sZXmER+SCEXYSiUurcWHfKj35pxzadLlA882HLpUYzVVIwPpOqK+jIZGpScJZjAqA
L5CMneQPV9LyXqJFDtc1B02NdG6fbqEZ4uccjVrw3zy8Qd7gpT9SoQpZt0eZeLzWpD/5ncs8LoCy
tOHRKyYmapiVR7AQDmxniQusxd5vrg+erLstt5jN6XGZzycCms4mqzTt5iC0A3PYGnZnmNd9pf6a
sya3/7tCbv+EdPFvbT/v1p+giwNOuIabeyrTm42uN31yV1SKgMinlT15yJX7itp1xvgH+81Ej1CL
f4GKBoZCjECxNGaGsUzT4NsqOiTzNm2cJ5Bvx6IvKcobF9xu56EOysLD/7hSIm6CmWhY27H9anRm
Uz0h9k+ZdhIPIH89TVIZKUHNHKiBHcMUhDECPVKRrqg8pSe7c0yIZx+EgwvdQtXAjfHy83xeAasL
lHq/EgktLYQJO2+sjL6AS95fBh2opSJv6haWiWIF7iLblStuYtY2+SaRnMBfoJU0HLMy99NYWDrI
vAmdlF1RKe4en/Id9wbHS03uLce3uC/rtFxA/M0VFd5huKQeTt42AXP7mDCWRQmbUnlYPA2wJ88W
iJzfvAT2pJQr9qjtcIFyGPIMh0JkWgMRhUVpYZRR+JmObK/fDOsKMKCXuJ4xFX1BLXX+DvXMAtRh
U9gFlJP1t+IO+iO+0Sumh1UihCkfGGF/q3MxsdR72Q0nuGQN4iJ5aastrlK+FkeGn5o/5xs6bncI
jRZTO/hhQeWJffz40S7YYGmVFCqknYqxmL6+JqQkXWpi/9T8sgfIAR00j8IJubUvz+BxrxUn3J+k
okssizSCsxLBqyQ6zzoZKuRgxWFktJqu9xh+jK+t5koXb31zL36OylOgkgfd9vAGeGmcfs0t0Rdr
bb8qP49EV1LkWHKA8gt+f+11p57O7QTA4BIi+2Z5EHs+0BNI+LfHktLd3bib4H/ZLHaNCm6Bt7Cn
hhAcPokrZ/CXjlOhUlOO4FpsjYGF24CWU9GbfeCluQnaSukO5zPu6BfZ61SNn6QgS6G7uYm8gqcj
ZPKiKFiecA8H29TWpWfYlEv3AOT05MrpchODhr9HuDY4kFK7x9Q927+B9fVbXKUbEQfsktswfd33
i4AFKi/hZ04dWUSwfjDA1yFCpscSgW8gGYeZWZu7HD/GXmSAlj62OeNmFGtqzhG0+z8VdFx6W4VP
Jy1td0dBrw3VI3Qxi+RQC2NITHLk/l6NOBTQ1vE91yZzXioKxTFmyQArlF4yuDdLXhbgdZRmNX1k
auuC/DBbmPaqhGh9fC0j3VbIEMEgGQJqiYaWJ+nabCCyEztnQ4455MHKoBi5NkAPU6s2EAyfY+dl
hNtneUA7bw9xOMopfWVbCaAowHYjI7Ul2lZCopOamMdt41jktxu/MHREQ4RBUJuELJqnxW4ETgbH
jr8M1KTg4CRre+YGiRVxqb8WJPq1B7ZRbIAjJz7mgd2TA4DR99ca3EknqoTn81brd//dZgwS24qL
y2jMyGnsOwLr536T0kPN5eGzDTq8scm2gdl4KhQyQ+8eo9vR1e3ggjQst5yCmg7z/pWMfZmYJk5U
8KS3iff+MjD0sY6anaDMrKeH7hwyNU3n1sVOEURrekAbQjvtAxvfEAYQmhgcBrmR1WYr5V8iU/Lf
zHEtaCtCL4In1KyUEa5qT6pYUfn0pNnO7JTFegnxdsUJi8KUHVR1a3Fmf5WShHn9oR+Du1wsBGBV
A2mhyxTo9LCb6WQ/MnJkr1zBmqN0Ai+ZJtiy+lwSQ2BOabR6i/Iz/E26LQYpwGyni936QpG+a5IW
raNSNjvr7p34KMmwqAx+DR/qtYSApc3x6FpC8ELwKqUUi7Tb1AyQBu3XVGVgRspAbfE0afZpSidq
JDv0lJtH7BmX/YDr9wMc/x03A9XWAhP1WyfjHpFy38AvP74k9nzC+Ftx0jG0gDSM/v65bxnjlx4F
fqQn4kyrQT0yjsd1WY6ArMelvxTttvnD86jTr3gzQfjcDaiMFsXiVnLADTwMtouTgQE3X6rkpx+G
7xwRjIy2FfBal67/PoC6GmKHoMy/FiHQbIzQPdPiik6rmX2Y+m2xsulRMtwmFU6pbdQAFFqPhBLi
jDiuOGavovAwpw3EewzETZzTWnmMaXWDOjXZ8z03D7kL4x1tJLI33oO9JuV5DyVXvmSxaZsflSLo
suiEscIHeatyTDlXagUFMEzL+fwdbldYiKNk5UZG4KXroMVoUm4QLsB7+gw66Rfts6o20w2L80PA
Pjr3XTQk9+Ec8H8mGdkzz8Y5wYNEcB4L2gf/2lG4UFnWdLElhBzLHLDNk55ngMVoZcHZSFIQFBJu
cAtaQmWSnQxltgbRSVxg4SzI1+9PXSV7vNow8dVJDS3n5p1jruemkQUIiS3ZF4hZ8dBkPsnyO2WK
scBb4cR0RJ1dIi5HZV3OLr1nyPZoPKexyxM67sWYmHogaRsdfCu8xSZcRl0QtOucbVh6gFwqUcQv
me0HLoX1VgVA8/E4EmJhi1jypkCPMr7crXk8mJ/Izk2zNJ8UhSkn4XQPM4171sTT1JNokMP+3BwD
YhFIeQm2MuRf1j2L5ryI1eCmhOMtw0m4b5p/We38heaGFr2CwCEgL6Prxaj5ox7U2MEP1oJSh6DG
aqSvGSD6Gs/hhEXmc2fWjhKQRQJXNMPMV93IWQxb740xvEOv8keb5Ej94uT14OsMYqWK2139FSQI
ekkJuYSKv2KzRMyyvrS6UTZ34Qfg+T30flfSRKaF2H7YyxhSNVm4rVxeSMmYqv+a9OXfDS41nXty
coT1ZyKgzumDphdrkQF/aLoUxlJwWVuaKvAn//nFk8yzrHI3rxa/K9BQITQa7ywqvYpSw7h4gIYW
z2WyvL8HPy4sEhSnjiQKHziOzTM77OE2/+zEBXhfNn6Z7HFWp0skVRX+HhtsJNIBPqRC5f5QQwpO
UUBguyqMNjdnCsI5tPlgOnPEiywlr0GPbmpXB89hhOCaTUFkG9f6XN9dOffq7t2zEqwuycpkeCWV
loJO+TQjMsODvUwhfCiw1L10i0dsw7z3wYFxvgVxHDGzP1RYgfE0sfm0oqeNzc4albzhIQ6dpaUU
Soaiiy0Nx9uVOWYh6kkfYFZwDFBEJjajTdZ17dxwO/Qb2RKHHhaDW3ELr8QM+SfeCB6a8QGVMG1S
1flmPs1pq+Ez4CT7lzsj6muK8oT5QD/QWmUQULYV972bzbFGapNR8jieKkEBMEHedWRdvRJcWjRg
wE1+dQZ3T9iFGIZ7X1Af6xw9l380mRU7xsEbAwTEB2i5gecKQ0GVJFyIFJ2L9Gg8fBHkAbg8S3yz
1nY6ZMt9Dj1uWFjLek4DounY7y7IEEqil5gbPRyAm36rxM/lhvCWe/yQc1jJf/K8k3/WjFN4rrlg
Gv3/RGO7ELRF14255Fp+2nYVAz0EICfdh6dH+wkdL4h9HsrRSpJ7VRN7qxtmUGZSSEir+0XdVcgk
smjl1+R7qrvYIjSwIzX9Q8qaCCtiDPZQ0rdFDfe89HkpI411UzedHrToy2vqA9M+nIfa32dOYKdW
DgoZGemTi6OLA4vDW0pZW6CMMC3LxhPFK8umC3oclAIv74PSytajYBXo6teIVuqgJaAPBLIyIeYg
Yfl7zmj+pRWx8Ntge+koPu8QfYbIQo9Ien6I0ktr+aLbOIbD+6kQ/8mD3FaL+EorFW3a6ZUhjH35
ilUIppzu8g80+afh/TpZtSJz31MdBnlmXDkze99m5siAbvWWV36i7PA1AG4K6pskgQYzjq48mjFI
mxv1NNEcm4fKqi8hrr6ifGIG9uOOt6XPHVs3juSW8z6mTnXq8uRtufWLNkriW9BUQ7jLavOv85N+
xJzM28zPSuTX/JJ1Gaw5pJ7WR4J4oIKk1ihlXQJTM2e8LYHIcj5yn4okIhL5EUSlXndKhd8Q5lZF
q/W47bcGNrdTpTYxrp5Vr8ysjjBhB+YBE26xd2FjrgT7Y3xosBQpx2l1BA4V1B9a+Xd0Z/0BdESh
F7od3fevMDc58cS08ZqxH7BaJH1zVpQpB0hzLqvENrlZDNPA2BbXnQ4bjkdd44iOfMoQ/EWVyOyI
z1mHk2Aq3MX395opV1o6EfF0f7SjbN4Ho3NsXdFafTt/jQpxQY5I5IcvhrbEDiD5RsVVKKwGHqbN
+Xszm06ULUzmDPtTdoB22WRO8LCRP8pYki5Qr5iDHnyTxo58zrG/dH0rtdx+1w61617lr/g01Xqy
0VzdFW0XmSzaBybSgQyOLcg2AzTi/CzGYmmVc2LIrMeLvwzTS9bvmOgCQNlHXemvxD8tykVJz5TY
yeetBKSjj1HKTGHB5x/V+rEZb7nkK2XZEDVi3PDhScfItJ7oqqs+viQCn68vPd7jt5RlRicPA6Su
1yNKePlNRbPhC29KU9hIFussGXF70QToQ2hdR0e4rWvRiLDcq62kh2EhDQ1xItuoDmwJf74nahDA
PcmgoMnPxwQebqeWJQY+Rd162r4TX9NaRJmWUTEy2nTpVgm9FXQpTf7tav+BLizKCvsF/B+iWC8o
aIeeFW3jJOmNDjYMDqlZuY8Y1AeeX34yEIopr2t6ZNiPYjFfb17VKaG7jkPK0LpfPN+YlT618BLl
PtjcsxnDgNDAlRrAegi6wt4VLLXorwzlhJ1z15DuKj3Vu/2xaTLmrLRiNd8uLj2M+sPGvR0lmXJW
cvwWwHG4/mcFK3Uqq5eHRvp82IUxYJFX2abYlpsFb9vSzgtuYNUtJS1TO2TJo3PGFyLr9DN7qlws
LzHgaAbFLOMs8q+UtekMt1+WOkIt6uNPIDoOGBGf1z4yrZnsf36okU4uB1OU3azSUkwq6zAVNezT
nXG7N5LnV+93eHxJ2C+twiCV3M5rAbPvK2JLMLrLL4Pa76kQX1B6yF78xcwZWO83Z6ihu3qPGwNK
8/P/Wc9SbsPLrJIQ9Pmp338Y4LUyDPy27r7vD8Yg9cmSCfyoFlD+fGNjUpVz1e+JLHc2k5BUMGYI
s5TMpYshEzpwGVawOTXaW9+QHo2gyv0SstNJ2N3G52cj70rjuEv6APNfnN5lT41sa3Lczi2rWbT/
QKbqPZQApmCXtzVdWRWan3povKNN33C+xcFPxqnjb6Lu0dPBoau8hB9ccPIBqYT+DYURe+AhKgQW
b8IilY68J1ZNPL4lu2ggZEycvwRPLlyw9qeyxE126Wp8/tQ3np4XU2sn1imIYmvMQOrBPI+A3yDO
xYYh5StiibozRdpo4jIIAe6Kb6Ccuwk4du2rAx5kaqKyuZxoLB+bk1c7KrC/rsnSDbT9w9nVJt5X
8GC7tcY6QhIPg7NViT/AAh4imwYEi5Rz8fpG0gJuse8cq9qVcc6OzuGjVvUXmKEH9tiLWR0lcrLV
/HFZAsRbhfL3hkM6cGQEjKkMyfZYavT66P0bvNpipqsY7Z1dqcA2cg9vAol815gjiXLCdl0d74DU
eTkUAyeCjcssFIfHsRu9lub/jgdwJhVoG6nrnnU7wF12dupjoo6meQH8VABDM24FZUkTMJH8AgAW
uij14+aDc1qfxPf89r4DnDt2u/yx4ZkGKqjyGECPgaRczcoEQ69Y2e7ODj3h9XQ5h+jQFvURY8N/
oTysQHT2QY8yBA+vCgE8EgDvtMBlMs4S1VKyvJIv93wHyAwQ5n5GyuHWY7sD9mN0MGAObbl9Q6tD
dsigtQOZAzWq+GuNuyQJF6ypwTFLHjvMbFxUXLlpTSVY1feYnrat9dXkmV3SHgmKdMZk4rHEnKYH
y5/5mDOTwksBMDVHgI51L4PHB6nBgHuXxJoD75bm4v1PByq5qrEKeU9747V5qM9mGHA8kym2lgic
onTqdhJtna7nRQEfCewCrKOEsV+hxh0fJ1RkXsGfNZuiJ9KZCP2DBM8z/ZSZncR+bdf87cwQAxyX
aWC1oSpwJVAv8388MrIe4pxuhsXZAa9hubpsWk2f4Niz/NYMnrTlGs5P6oICZeaUK7apGlzQ1Na+
Kud2D64qv0uq8Nzpti8e+PbkvM5C9G3IzjUaJ27F3lKCzODNr8gU1z7bpcyXbxgpa0KZT29cA2uX
UF7MTOsrU6vuZyOebJm9Q8uu73AoLgDkRmlxRhTWG5Yw8e7O9Ft1//Z02bfJhq5SN6LBPTzgziT5
9X9Uxbo59xmEdTuOL7z0ym0mJRMCVxgsfKgfCdjSjyZFSNZJDuUfEe8v4GzRQ3bYMyDrcly2W3Am
9xInJWO31OoNASWemk4DYGrW/l/Q8sOyrV8cESSQB5zpfJlHUHeO5bVj5YrYE3NbO0QjaDQvE17T
9+ZYWtS/MA63PmkGxzieLkYcdA/xnfEtTOVgQejDhd0DBvFI3H9QgxeRhpfI4igcQ0k9T2O7rFuG
B3x2z8taQY4XBj5Vruwn6/jlkzyNS0whxsFezcaBzJJU6ziwDPOX5oorlEQ7KiildZ/s7E/j8TYD
HHNeOki5b0QXh6ozPnc+YBGTjr/wOMgDicib4ImJawibg0mX1uARLWQAqGrNVvPYra0oLM1KkWlb
2PsfKm2nfaL1zJ62UstblQK7QdGmKD5HcU5hSZliqE6KP13OPMddG8Jfa73XPKhezkE0gpIYY3db
giEr0MEs6evKfCITho2ubzTEeJhy7gBkL4srOgLV/UGafz2rRrGVU3qJc1hv5dqFROJIlBEnZHpO
GDGDOwUvag7GEb8ttWQjAHwRnsdbH0EtjdU6SuO/GBpmfK9fbaMDRsJHESQck+xF/3Phz9wXxCQW
1um3/8ExtRD9BCjFxmwJae5rTz9pMK66qbkJIRYHs9ncwj3eakMrdo7RmX0Y0/WvVuQiCm/kGxwK
N7hMhIlGKJ/+9OdbSH0dDuNtUlsgAa1jC/786ZTHVZi/9lYWZc7w8/g4DvI733oNe8bNjoHA9kIn
QMfVvPhmvMKTRUp///YCNkQ/7osR1TVSF3kBbugc5bEDsoL69v6wXajY70VMdlOgknb0jvN++qNB
gaZ5cT+P7M8Q8t7zXyW4f89zmyZQm4f4h9T6ebhmPsMMQzZ7q9kGavqV10NlzQw7jgbF/Dw1/PhD
Dz0ZAwz4dJ3w+hjbcHk+dyGAEhkNfErUZD0fSpGP+DxkvF2NlZBKKEO31SAM0zcZEygQDK8mSIoy
NfqsX36MIPOUFhxmruzhNncq618kOyV8VtOMWqPdh4NBa/lg67d+4l9baVD6o+hzdVfr9hEUaYrx
iXTm53Gvbd94UgUAOYy14yY31sCEXm+EC2i21hX0d4o14/O38a3rUIzXdI/8PLDXR6l5SkhcO6Vy
bLuRffZhhQDB6ToUVtktQBvQsMcmwhxniFHjuL4tIrXWdrHwQnXuqkQOmZ4HPYLAY0DBYbjdDZsc
kGT86GnWPNAkBjpxhLGwinu7fi5UrSYlp7ORKUbzyxAxDnriXxaQR7Zlm1M288mhzk8Ec8aoOvZm
+d7FvfEGE7UgDuyXJvDfv221lsLGue4/0m1l01YD+8a7+XaSndESn3QOzCReyMkssd2IqB98az6w
rmpS5tc82jPMJayLdSVJKpfdeWyKciRGaFV3/vp6Lk4BhC7Kkte/9pJ1DlPZYtycnU2juRwM/dJT
z7icQwkU2S9hElcFR8ej4wQjlfuPiyiggL4BqKsfm9kRqQOg8CF9EEUJdqbPCnHcDEJ8cozc67Sb
EauILpMvDKrG7yFyoZA4nZT0fWBrUI9k++IKres0vlKMKg9JcL+UhpEhwHRHZqhNP6DSrvds16R9
Dtm/72ebco6cRUI8AuYISq6YuTUONDpBBaZEtoz96ktGHdWeEzOiCVf/kYktUo0qXGTKkZkAdBrU
Rv3zcRQXGtW0R/M8gheJZhwqDVQbhXPeUiTrkHNcUv9ptWKJ/XT5IWbrzqiVvH2uFZWt02/9qA7Y
3URaBB+FbBSYsf3q2mX0gAs+0Gp3lOxv9pns2sRBQv+m35LtmAu1hu2pYIF0MM0HhUCdRDEjEHaC
xqVH74iIfe+dz6sYOBqY6miMrF8auBLYVY0ayrggCw2JAhaJcAgLZzaXNJ86JUsn5I+BdjfDKOZn
Qmzxv3jKGLi4gsiBiprKsTpu6hLwVbcnyweO0Xib8d2o3AQ5WjkvP98UVDaGqs87cs06o58PLiP6
zG1IKYYlqXBn1Xs4+QhdOyOpuTr2GSmEiVc2jqTJiG86KJS41/tnAzzYcSr8UihjTkixRd0lj1KA
gtHcyqwp9S6FWj/lpiZMlkEoysw8R85rMSIE6TSNNtVowzjA5yLSgmxicAAoX6Y8GhNqSzrvnxCW
XAh7K1vPqp+5KwoLcQR+SeummeAaRu3pDvUUivox5YDVopkxNutCatRvpySfcDpm8Mn81mvCJ+YI
xH/ubPxDxU4dWoZ4Vyp40CHcuL4gyBuVh2sDAbtVGnQgeAJzRitAv0kOqppiL5DVoYZhWhKQcX+y
LLAwT5ErtR1X8GUAbnXQS5DwTy91JV4uNNSRJnds0mf/nBvN7UyLHD2lTmA4U/7h3yEaatvxM4/c
nw67lQv5cKbgAc9b2XJPOqlljO+duWR0wSb69/ajCj8NAQUrOmYy0SuL8kCSLdqoS3zZO7+VEbcC
7887o616z5OQWMplVPFN/JVmOlitSTVyQo6Od90UL0W4dCRejlXT9VcTLND/X3i5B/8vH0ubkUk2
Idhg6PF7X1CGvfJLXorMnh2ylVT3R//sdQn0EyfIVhtVH9vi+toxlUDvvugnybj0gmSwS8AvcJc+
UoXx5MSbCtbONPiuWLKQf1cgapr+9mizHqCVHjc2fhmpwrpqnBJDxhWs+TGCcqRFSNkCzRMblpOD
7N42ImTjEvdaKk0O0+gQF1+HZNErRB9G+SLq952pBjBtKt/G9koYw46b6GOaVXzMZIYW0y7mDil/
hVhFwHdUlO1fMPktq7T5N8e9FaXMW4EvlNH7OWa5vpBooJnUFJTa3ztYSC/Y9Zu6H8wGWvetAhOc
/ZZ7wlrNJwr0NBrBWE7ugrwHB631n93LR353CVdlu7Z5pH+HD7YuIw14QUvk5a3O5Wfar3DzKGGf
ngvPswfCU3ZyWq+IO6NfqjtyyPZSRkmcouOGhsSUP3IrKbr8lgQMcVzX2nOYiMXCI1ZZqRZGQiaJ
pOp+uholo9P0C6oRTOHilShjaiRFA90ifTI3YKsDkW6frv7SUi7sJ77ieAaKKzKajuqJWY40CTVJ
eUXV3NFaZj/y2CfetDa/UT6mtHWhWlWlTHrjZaPgglAL2le4MmyfHtF2B6ELawSWXosbgkAWoG41
tWAT5hcKQ/Irxs+5ansTc/X7makTHK7BHQ0/yuMwCH9+DtjGTT17Qi9l9nJ8Qj3zWpbIJWXIS51b
NbULlYPOgBtBaTm3GrTwe9+BHhASs+aUnojImbhagy+SbYhdCLAnM4BCQ1w85YbSfOtKVoiEdD8/
5PQ8dP+algWip0D70UhAQoLtmDxclsrUN1WjL5EN7KhXguYivGJZDoQC+CPueetnkEnykkDW2Sr+
yBowOku6l2Zj1o6bHkjIf+xZgazpU2wiW1dvJnRAP0ExFcoI/68IY4BLkvgjb3AhClffSiJGYksX
naZAeeAXjVlHO3I6Zjf0S4aY5QFOPORX7GpPB/x3VkAGurQ+25O6Abkn94tFHQg255xHeVTXnEZV
V0KEBUJe7T58Pu19CnS3JQOjtVYsIypKYy8wu/ilAjMUJ6XIJAP2f6IoeRVrf2MNU5Xoows48VL4
JJljP82Zlg84ASUFijBO03ck+ElVkUCgT+FB8lBZkKEzUNdVkcVdTG1N/5tY8gwh1KpYICRUMN32
SleEyZpau8m2Q7ZHEANUSU+uodCUwrxBWBufkvIjaXMWX9Ly/qyrmlUbZgGiXKobwRNnJqQH7FFs
AHoHnI6DiNfWmE1xE0A5DqOkXgkMnkEhFEeDdG+Z2BDJGW6KGjUgCu+lcVWIsmMpJLoNHu7WJBrn
j5KU7ejDfQZZb/uEPDKOPEazD6zWw6fVsAsPD4ePn3EKkbXSKwi09n1YAzs3R7fsqbIUBtxXDHft
dAqmiZOuiErDFRf/7A3UQIJw49cnXCWydHan7YGJXGGwGnGv633OtcQ5vhd1VBCAwNPdZdEItdi0
5ohGjtez3pRVf4RL3Qxm2TtyjRYTrcIvGnmo2WPr/6YTdNiqMsCDip5vCZHEnkqaJ92qLkXFPPkE
LsHE2bJ8LxvBspxuL0SaG2s34xNTR0A02mA6jxs22lWRNbli88SysCGgkbM7+OnGVuGC32lZaxLT
cmR+30zItoRjzFRb++ibYmhmQHcWbcpKPHtBSulQYm86ED/7RLnmtgOWEIGZUJMMzRTxw0K1+7KD
I94c8jiOMsm37WzWEi9CrD6E2ctzkkvCTbA4P/ziv9l0D/NgMR7aO86FZ4ZTrOSOXWW0oRSzk3eo
QpkOOvH12KHfEDex02rBUqGgMde5Im3Ksad4gi3GgefhKEdJn5INOMJz0+qcBy0AF5RzgpeK+8jT
shuPAgCUpVU/1fKcCBPCkGGD+PlMCpzXmrMJw3hZAxi7qIq+aO/uVtTM2sifvXdWvbLJd+HNmhjO
iYi/9OVAh90V7R2fmFNAoPFAAiEmQ+y7+BG5PXU8W2DQfa4lNlCWauM5e6C8Uf3oeuzQsHzmmVZo
aYYg1SmUsCqL/9z6Iq3bCHgOvb4THVuk6auXC+Mu+is+G3MLEb4j2Bnyd1oS2YmrzO0gYzIkDE5C
y3zMgUQXyIGMUGhfCbeRjTQzkFh9XVQUDMfmJLIjBWcaadbGeLHPnFaWZ/k0AhCY21/gSCSavwkm
myZq9mKSFaub75LoR8VfdrBzyLp1UxOoFn3ABuqGj4g5qIoptly1kaGhFFQPk67JQaSbc/L+Vzww
C8cJg4rnAxNAQnHXG6H1WZOpXMtcHOY0tBD6a0dbMylqcljAOtCN7WOqn5OP8bSSRZ3al3NSU+TB
/lQs2D2b9RnSueboilo90gqGAs75RWhwahOfIz3Sz1ecJ2k1YrzCk4dPqlDuo4dLJ/yLlH6yq1PR
5nxkYQt9sRNwxlngGbi9dAaMAhJ78D0zC3eowTB/ZO1zKQldR8/aDcP7+AU2X0vpBUboJ9IW3avg
fa72KfFBa3B/Qx9SnDSn6dSnew348v4KINg8F5/lDYy1fZTNzg09IYH90kOxKB8wpi+LkFRhhgSW
gs299YqMdtdrlvQAsxymuyNgJNZbEfVOMTFdLBfHQey08GZxt0CA+h11qwaafshmnAgCEpyKkzfP
sSxOMvAeUvcx8BoA48m+Z5Hl2+ewwf6EZ0MTSxUt6CsUY8a70eN9tvydIvwiyaJVwbk1uBPfKww8
pmdtFq0SF94qCIlwYIXu2FFLVkBk1hDvo0o5vRbVk2Mz1Tl2+wfGNb+FPPkvP5KTsuoSbnuP+ey4
fwvw5kKu8DVm+7hnuy335vRNuiChbVrxrfm6XQQs1snuGPoDVq+XU6xYzH/hjeUUYN8yxY0cNhZe
s47O6/IIJPewBSUZkMiTrY8dbeDISWzHWkThcjZcvvx68S4WGeWdRZUlIVOd2nelWF8A7iqTaY92
QHZZcWAcAIR9Y/bDZnGJ+wtamGySn4Br+KUnvW+JKYQ2enXMtVLtBLt+L7LlB4zkqGZA6K692rFh
4mwOLHLJ2OkDg/RJYNjGE1pjdD8SJpx+LZ31+n7Ays1rskoNrhFzOz97lX3dUZQ5cdWhAKurIqa+
dKVnrBZKrUHmHUyUES8PUD2BuvFnSj0f2Hv/1GPylYzotLrIbQItSbs2h1e2AW9HAZD7V+D18EJz
xlPmjhH/DZrXUw2KrrtkMYTt1PfQVrE5vTK8qynZ4aRrwJDK9TswIQfQUeaUiWzTYKY95x4ARqx3
lK4KUzstR4GzW8/xrfGz08P5j8NjsEdazC9GTDVyX0r4BkXzPw8mWBNUyjqEZ8HebZv4Qj4EyUNS
gY7KBEamVvsUUwg+fT8egP2ySOxXJv6HdBe3eK0CG/W5ZNYyorkwt7OVUI3ILfYAwicpOeTMTLeT
cEibuRORYwpMm7z0HDZCTqJ4c8AvnFYYtkQHIbZpO/kZgRksDrin+szSNeoBxsHpd1o7q73Ya6zU
C27iRK7gLuOWT9jhJH1bMUp4SGMCLuR7J7XsB0GpRNDmWQ2zjwClPJpaGNEHKnk64Xvi1IQUaGhL
rtvHwp54DZWUaiGJdsrj4+5p+9ZihBeQg1G3ep0VdEfsMKqrJxtvkBxxujO0uLBmB7nKukLzB32N
Qp+aNo62Pbl4ND2H9+p9L/gvrPQ+9ja8hJLtONbwTwykMXiguCiiumaAvdnr4b2yIaHDiIa1qipr
7/La7eO468OpPKaskbHsqMQAFnB7YRpFSXnSR/jx78bp+v/S2LCKXQIy5LYdv/0GBOtKnCfzfG8+
UwIGvXnIt8Vbc43v2FcN26GbXMLGxGsqPNmJ2uZd54PCxEB/wvIve3o2AwHkmP9DhQPbym7C1ndn
tEcJnoaxd6uNQD6iNRNCVhmdz0q19r92AcTi+mAWy5cLUgXCfpz/1rgErIHpvdwTE9WLY1hSlBc1
8QQ4X71b1Db8Y3VhyOsiN27QvB4O7OQjVcrFsoHP/LVkXzH9rE0e8kCKnp9ZcFXdF+rof8EIf4lr
RIujl+4oNTpCVFKFwsgEMopl8AUcElv4UVW1oVR6pg7MfgI6nUxLQVruWOkE9YNAlgVzTEMLhjsu
2dzhdRwpB2lZU//1Q59TzdWgeQmFsZqdR/anqKUOp0FCcGwi2gHjVOGOIyp6Maj9hSuWfxR3+KtP
NPM5xYsF6JcAadEHOA2vx34wC3DKd72ZUAOUl8NJ7Sq8V3JETpdh83ETtIX0qgtHrxvxAtO2FcMG
SKyv7slFOQNnouoact/n3QL4EhTwt41Van7Y/A4pIr8uhf5+c24BvrgAoi+ESWbwd6TatVr6/Eyv
jyyFroRPRnCUIDaDd3lBGGvcSw01woo2RpuhgXxnkPAlT25QOLSFZ0Ps0Qq3d+fkH1kkv26f31iZ
3mmo7F1vTbpk8UhR0dmmJO5S0cztYSmf/dFyKBbm4wZy3FPleAKnKCtbapSPtChgNCQm/49CjMJi
6D0HPDZKUM6glIYkM6YV35MPxGN7UvmP1HJaP0EA/VNZs463uV0S7vsB7wKIBDZtEBHWZthhyR4P
gDFJsqaEsTMfsuz+IU41wlcBQkXsjOlmf+kBkUFguUK8U9Be/Ri6mwqNoNx4ZTxpMq2wsNCjemRE
sHX0jbUHdoavic/MSQEJ1cQkBj5QvWz/k9bVyG2uWiYJ+4Nv6xIQJode4m1XVzVgqXG8Q+EOTJx5
l+8V4ChE6JTrxkNRxUebxCGTW0SkSJbt/KwYvT1Ao7boAJK+cI8V8tiUrVdKNTQj+BD83xdKawcw
zczQNWckrxb1jQ7A/nEKayDoVlU+/KB7hggq3+zcosqHkFxmHbMeObuNTXA3HVrVXH48Y+YQKwHf
N2A6azjUVz1gXdjUGEDRPbVku0GJV1uZHNwTBDQqll20dQkhIyO4TYRq3od1IA62+h5ZfvdmSG1t
T45wbWM3aoj2x957iYYGnZ9fJuZWm5SAmF1+Egr0zusnws1ohGD9DjclM67Uqo021rqNPEQKB062
LH7++mIJonz6ueRdc1Mj7SlnOJD7IrkCLhj3aTcPuuv9xx2WEu6YQ4doTgmfy2p2RnQKXxBhbDdu
ZEAOxzMaeZ6C/K0+NUSWqAB1DkSX73nuSaaF0XV8b983s2hPRrYSSzfaR5UVk89xBlb22PRpbok3
4pJeEl4gaGJ16va/Nk5tGtN04cUFrGTXt6jiwiU15J1+naZgL4fl21p6AkpY+dto71GGdXhjCtAM
5jEiK7uRaSpBgr7sS39h59stVv2QO7ms6o/6pXVwSiq2KZKyM18JN/cCD1eN+h7brmbCM5ue2rWD
Yp/BLB19cilX3N1fg/+Ua94ZcQXEfnGpZrTltMw0CxHDj2EDzfo0gPngch/rjRCACXHxwkisum1f
RhFZdqj6ITPsQ2DVFlYj5a2vm9+pVGpoMY40FFpA78cZ9Uf5HhoGmmDpN9v+fAWp/gZZzI0wLQrh
LKnB4HmY85VrHBXwzRnrawwwUf6XAuGfrwdAwReVnw6tO1SWd/RK0m4/RMP8xYB2RLQcb0hs1sGt
BUnPFMF0R7mkTvjdYtH9qcJ9oFI7kVdVchIZ1XAAhPczhl9GpZ5aBveLdK5mlzclMsWOy/XM2XkB
u9fQwpWh3pBQYMnQpQAsqLt+J6GV7yMh0Ma0HwAJS1m43+7BTA/5QVzFL5zrAbyPCHjmgVIFQs8J
DgT3W1F1EyjCia6LC0pQfRiULz9+4Xo9qnfJvsRBoquiF1sTA1jBdAd22Mf7g0xGQyl0N8zqbVjs
mz28cf9tkadUdtShgU1Ni8v0eGgmOpgOcJQgjfvYeyoqVCNOLlRBtJ4DnQ0D6jpuLZN31ZxNFIH3
wAfQFMrxebWvuD2GEcB2IZj8T7uC2wkuHkEhm/djJUFvJtjV2/YpD9AkQkMKdEthTS8k5DVHthRH
/FAnuWB7/2iYSRGY8CKB+2oryCEGaS3mS64dbjaUN6UAHGSm3UMU57DnkeTRJvkSRyivZHXcLUSD
ogsqt4jXIe6bZvBJsL2e8iDP1aZ8SzXKfOxs2tIXaOorAuE8M+xEUl8JQcFKUYd6bjg7kFTg0kcY
G/kso6gQIVAbYYhCdSO26/NQ0JSten/5NdNseX8bTWRuu5ZkM2XbVBv1VTpfbNUQXPE/hc8rZnc+
3gP2AhC0uGlcF9m6t/nBncys9C4AlkFzI6q5haX3p2KSEzIZWLHpMFQaE7hkCPL71tehX3Me5LOB
TxHWBRReSUa8QGCh7lUZ8TFym5P8t0QaeBmXuMG4dfY+KzchgYDcftfvgK9JMnNkLv6LljtKmFK/
S8N56cH1jaKJZLyhA7EzLApGLtf4msXZzh7+HP4B2cZHc7nh2omNypUkYBO4WU2cMOXbwNnRaLN3
QeJSZqyCekCCE1vNL5KYd3Fl93AdEAZXWy2Crs5iZ0NYxZhyTzTHevYyugnbaetXMjPYNJ6gLOXZ
ChTNYlaqDL6ucTxu/4xViBMvp0SsIFOON131yUgLY2Ss2OXkizV8A+tOGYj//OIZ3Hf2oTiFck6p
qMMsNSjLgbT4hyhwU4mjizR/8I+u18lDAiPtbMVatfAj/uu7YTESLx+KEQs5v4DIzLMIY46MaWQa
AxmtK30g6qFCk+Zehg4j7esWgZ9OLsIqVwxVNEd31U+5KGtMy9J9C2aXbY+2wpxMdWrFB9zvuPQr
+wI703DDXNgpGAhbdku6bXQ54pBNSuJiedlVKXyyEuJwtKo3a0Nll7DDplfNLs/Qc6qRdKBpH7OK
SQMD0QErcIJwEEkEBIg04/dY0AQZedkr894/+ldS8IustRkxgws0BpHTyLTDw2/Q746qrywEoX/e
hjEWlVePhpag21w/S2wMMpMybW61v48Gf00CeIYLMvwuKrDBSU09z6pZ+8lSO0E53cQ8Fjyw5rQW
CiL7C1RCLi3JPF5XnMvVSsOP8oMrUeILVnpW7BsjDfI8Sr4KZVMjEV/XxVE4ewENLn0sEZ5ulxD+
YLEoSF0leNtb9BJk6STjZ3JYWEdTt6E+X3znnic9Fbmmw/2IwGckVK2GoSvn/cd54HJZbNk7piZo
9tpxWQ5ICYPQw73TN0gycYuK8SdMux6rLDT/FWXphuzJVfI6IEOhhlHZvMRwWjLOLL0fdQA1yLIw
moPbalFs+TQ/y3ST9rT6fS+vBT9tV/y0Pv+akLum1d8s0NGT9bUreMNUB680otQWgs32LqrXS8Ih
HgPNI7qvub9kJSNTzXnNf+AW0ybrZnpYC8somhihC+XUEQXv/z0mrcTZFSMQPnnXQdIoKYzdfyww
QRHtGuXGXfddqKBmsV7FEQBkZRPN40JWGBR+GzyJga1YKt9dVkLJTDHQhHoUgY/lnVeIh0OEJUJn
HNgVTtOzcLE0uSokOV7HWnGNZKMs5/i13WWFyXwo6tD6T2Lr0rDw9XIu2GMjE4QgY6kj2au7N8tV
Gerh1cEuUIkd8vRyh2FksN+X3Niozf/8YZPyc+6IrZG7ArZaNuHdq+IpLx0ZxU/UNsZg1IJRIKLR
2YPQb8LnDC7BBl6TuM35XMa7EFzsSbizit7I4Qm5iK+18KV/2xObK1p2G7BpgmwSfL+yMfMAP/1j
4sjB8KsLXu1xuAQzhCPtSjT91IeC48RSNMptFFUn9UV8XiJKZG+7mPHmrOhT/H2dhkH3BvDmsphw
/ZNx74GHyCtYy/YhPI7fPCVfRYu4bVcFyUzeZeXtAWqQlpy5k5zjYtvgL7ldNPVBC48kJ5s6j1Rz
CWCh7mfqZjf4wae7s/h+bph1v5mzLY9sQAQW3xKxsv1ToZJaWZLxQ2ItTWV0hH6+LwSUJqfogHSc
6y7js3Av3QWGYXT2IDNKWnlthUNn6PDBp5S5DhEN+UoAjT/4T7pdI/JbaY03GXh64cnjDxv0yyxN
wkeRPdMzktWcOAAiu0EX9LcmgAYgCLkIPEpvCxSP2nhuuGwQ6o75OHyAxjnbsE6jUm6SiIXPu7BM
CaxIVB3PU0CPmVH/siLi/tFbA5DT5ySzXV/AmIdrfSiAktQ7+WSs+X1gydV9Co3i91uQBXrooTYm
4+sFbQdi26fkImM1pcs8o71D4duxT5wdSc9DJG7OqPVr65j2X8Pc8qYojvoGs9jHTfzgzHWQ8Vvd
d9P1ikn5iYqz28uIW3E8h8Cnvs2KcsVs3nnQRjEyqgstxugYsNfAkuS/egWRT9E/474ojrmrSEho
8NWy0+7UQFPFRMZaX9zMnEFBldULN8rmE1UdaTvtNJnkeZaRrPww2liVj9NCUuTZqWbHfXj5HDk3
GeW5yXvG9Jf2FRgYavvk4hCO8ZT7n6RpX540S8WAsO4osfZRUDPpyAeRbfr25LFgamCa/JlsHweQ
whTBr2Lxf782iH0pKX/EJHWM0eHf3Oo9PNdszNPoaRB1bnv0OSyT/R10y3hxhR2k5KPu3/GLYqKg
UIkVTEM9Wb9pDwqqM53Bpw28sGG0t8pcoIU/qxts77/8BpR5G7oZgOhsElmmY5x6xTp9Goq0iVaq
9AMrO3hD/4byGP3HqXLo0Fm09tCtx51216s0i2Su9PXBX7gfWEX3Lm7U/uuP7ALAWJPPB08E6RzM
ROS63FoMM7Iva9VEF26CrFXrO8SP4eW9YHAW4E9knO9evYvqVe2gFMdbLDV++Z2HTy4qPMn+2WKA
4uVxSYctbHwG3RWLHODjCgDlFAPeA946y4YfbBNc7lalSPmg6KymNY345bn5zEY/Pt1kgU/reA7H
F6qe9ybTvaW4XZt1JMiioLRGHWvfAiT7VqQqvNu4KDjsqYr9RbO0TqyGjRgdmfhipGXSaGJlVovK
zcpHYVeT+egeO5Uw5M05Z2VwVU7z36duyW+O8J1gJ15j2/BLgiIU0pooEPmSUozTjNeCnKNMIGpG
pSn2uB1OiD3Cf0izoI6BRL0cgQvRbtfFcLbzVy+ry3AV7GTPUORfJJXO5qtqLWD+yurred/L+qij
BACkj+3M961AyHhseAQzh52MafizCClrI2zpXd+bTrDsHoYE2ut0aKrDroZ24GEX4O9CkbgxcrjO
z4RQbIGmMm7JnBXqAX65sywEP1Vlx3jJe2enq/0HrNC6VQtQy4bDrN4flnPT5bwX1HCZI2RGzMnZ
g1Z2KVb6yRw+rMB2PrYJqVXB/bZBURlSpq9XKrqLvFbeN55jPYvXFw6uJUgcuc85LvkL3hDfoJok
Z2xQJ64kBcmb2kH/jT0o345nm5nNVKfvPjW6vbVoPqngsia+sMlIrqHMzVcDUDZ7ErClVYDumfXt
BDApD0J0zbuRLBlSkX9NlhUROciL+uB8CVjJcG5Bf5UcT6nkeBHfg2z7RLnxNCG961gnwLjBb5nx
ynAXsXSgGA4RuxHGUMprEfv2vu5E6W/t+vzRyyu0e48iX6IzMALJHCkR2vuVavjgLS+XooRuVX20
UhZfToEBeAkyHAlJyEeYBJ6LTrcFe/tkcISP2OSGCxeqDWWccCUQYQRUJFjgs7EbVzluioWopOVq
uqTYlaHy/4N+/njhQYujY0lDbX+FDRdf3amHBL7qMqJ5hf6M7I2DFtSJBrmSxEW45gXnGrsASplT
WCJ5Msi1u4mAsEH/O01dY2rgukpZl9KHUKbdZQ2uVRRVG6L5phlUq5AXRk3pD3IyaPSPNWaX0xYL
2Kd5KLCRTyfH/78QELfK8UAMTjk8Pd0nLJ+95aNvl346yrftQBgWwGMYdoU+VhBNsFivE9TfNfCC
9TY+gOXeVdrSbJAJn5/vGhIQluzSmSjGBy1vYFvY8T3Wpiry7MriMLFWKS4G8+WRwktn1XVr3m6u
P5LGDhJmGrgSoLUrBNwSJk94p60IsWft6z06Ktx0Z2NTuHK5WsBOY08tFVTVYl9fYjUcT6hBpXOg
z1V4akvkZYVTVZOfh2qbiisliwviwbpy44zP9S4kwJAYpEXhhVoYQxxMlDyPIH6k0sYyL3yWkXNz
j9lNuOvVRMSS2U7z9P7o0FIY/QPK6zvlbIjNqdSGMwT5hXjhPV/1b9EJZHaW+FIYtffB1GZ/vu+v
9/CaayYta4Qniqlb0Yoc4rMh9isaLHQ+pCG1mQ1Rqtwg65Qk5UhFNqzS5MrFLIe50qpAQxnB2Aoq
2H36yuIv7/nNI6JajfUeR///4RvDzvfIhrcoQvH89ZsCAV5kyhC84vz+GxQ17Py8rAEBpLvAXwny
kmiesZmQRCWpbQwVlLNnDz1gnynazyuBGPo4dMglgdHwKw/+RQB50KNYHpok5cg92/lJHfLvnJF9
EKUgnHY7M30QYJBIS4QwmanPNxmYboEBuiGrqaTs2dDwHiWxZQrPE0IgAo7U9DBPDiKOwMi2dlUt
srRZmueQUp4y4URDHH8q3MQAS1T1dvFO9/+NnJvrQa6f5BWtrEzd/UYvhi/apxMbTy3Gdx+7ijjJ
/oH5TZq9r1YVvl+0ktR9IhW/E2LS6PNS/C5v3pO7Kk70XpJd3EOnmXy8UJFJRpmmcfizV5GiGfsc
/pT3C7pRlO0ljDZaD6QJDYB9JdlPMwdLrINwEBXeqNsEYwjGJm09tj6G338OQcOOYC+szdrdW7Uc
Cd2n/L68aKRUYY/tvSkb4tutEsl/avkzwIvhDJEphIBcrOx5NTF3QQ0DZ7N/P68eElPC9DLhFDcd
t4SJpyg+JDPoKHfsPhuoyoI4bNllCHQRO4G3omohG/SmIrh3uHjlMdkLaxd4ajvIuAl7iRM8rz0E
VecqWp3QB+xAg86feMsNFbOhANOP5QIFf89UotiHVZLadG8siv4GyTRYVYm/5ER40uqDgU2cruDe
n86R5NBm53UGWMrGHlKerMyuBIS4HFLOQm5LEcZyj8+WU43GRkHHrAmQW8fmUp21Jae3iMAM7c6U
YH0pFY0aZ6TChuP4cDpARs2QzZkB3BNSfkYQbL48BCUqavKu6zPAxWcTUEtTnCEhZLxj+j3hQyZd
yAuuvyCWMHXyZ6V+ThM5O5QMzCJtzRxRCmHly982uRwFXTHaHYCdZr8NTK3RzQ71zCVrtxfOm2Af
7eXuhaVplirP+8/TUdKHsC+N5aVpyLTMf4wGHSFMxUAJLjCI83NI+qhh/L98KwimYEADOBTM5/R/
llIyfKrcRxJW95M1KyiX6S7xTkNoUMgnHT38M1/DQqKiQXmGWOhzLMatuIww9ra8tOkhKyCcPLLS
gm26VxxW9oB/ZUDFYCTs8Rk9RPyBu71P3JPNUh7IWTvup2HumXO+zxqnSnDMhbHm0unPosWYzn81
9AY0MaUjpg7ZUpkhOH96/im7P/6hD7MXOKtqZlfeCftRsgOWEQfCMOo7pCG9KrDKVXjc5LuJNEUp
5DskvlzoVxffLshSCoSZrGnyisWWVaxejupKJHqDJLIhK9z/ayUbIlMjdBYd73Wsv6v0WNloJF4S
4cDBYdlDcjuDaK0nGr8SF8ovYSWPZS/tfoU24Sg0vbBvc/yWS67Lz73pxmMMPet7wJuFq1ioit+E
FDnBeUheq20EKkWDrjAMDa/pqW1DUcMUW0LMz7lFbmKKd9Lq8vjJVd5xlBth7sOw04wmEr9blyYd
CugNK/HCFZ32gJ02D7wGK4TJ4tJu29LBajw+jYk2hTeI8jEgMivXp7ucY0U066ov8ehd+tR+bbis
yDSX8cbcdUPBoHKHhwS5ijcLGbsSl9RD3fq6FHAycwPFm1xre2tRRLPzcodBCj7ECVosvpsHSVV6
MY2jhgGQG++oaZiUhsQ+n311ucKYwpKljXQhjC/3g49vqBxPDSyYjojy18Cbw6YUK3Uhs/STrKMp
1IdyPgTooXII+lLFgFESY11hMRic/D+/anZu1jhMWo+YQZ386yaihMozkJMqukIa2nkgnjzqYw0i
7RUn0rtOgMk5FosNOlaKXu2fnlbtAdVfAxDwuPAFZBgtjp81DodkoP9vzOSZi95mpR822hgGSfd6
F/+JOVH8oF5wf35O482IVZ68iEEdz5679+zWtGDlCqOWN/aCnBW1PnVyJBZq/ObiOkO7LhZeVmtg
PDGfqOsoRkBkZxlQY/28EgR7GWUsk9i92oojj0SS07/iM/JmXCMTsHsJ4pDj4UurIrRaa6bghsU6
g7fOaRuJX6LHHXEHcE0O0FrTW1Wq6gmHcd2Djq2zBtEXqmJQXV5albvFuCtFsr63dqkPkdZO2qEi
lCPIHSs71BTv0yHZ74/UpFW2c/cVFawPZs9yZz1Vv4uwLASMnlI0K2Icr6wLwEqQL7unm+W5m1Lj
jUQHblCmhme8IhDCcb3oeN1R6q+8KLNKooZ1M93+0meEBA5WWz0vckzTGhkejLdwm3KU6Lt23QU3
tVICNCBff7IcgnKX3GeJPJAeEOj/D8VuCAuLUX4hmI3Ys/n1bsWMyglFpfETQQhLXVUkapE4TRjh
bUQlb0iujGdORd1UNVj/boU3prJYfBsKrHMIJQa75Dxkn2oY8TqOWluj8VfIff9O7eMkP3j9q5lu
k7/dAFhLNbQYQdRlQo9hBmI6EQS0QPwn4N0PC6PMIxLidSers8+egdMtqTORlrTCuET7a4TYJVRK
qo4CBXIlEdJnDHayR+kaboGOon/4/WT0auPzSrVvdrgRjXD7VLHEjpeuL/KhyYOIk8Lq46zX/qwJ
cv+v/54OmQyn4uof4gxgTtTxh3hs+BCBFnJCnX+cNKWYQnRGe4oHi+pX344vJUTQuxzb+BPyrJKH
/NDvKaW1M62lGPLJoIumlDQYq/IjQsmcwnDe5C2sjes5SvkCeL9yjLlvUbN6WULpEz9qm1RAq6Gn
QUWC1aH8h/NY7wULvGDFjh5DxSSXE13HmKpvIesUGhppo63EqLBkgj0g5hziDte8iv2o2KepwK8Y
it1k64q6OP6QPAiozglCGrEoCkwBQpHoHpxpLPyuR9E+OGyah0i8mcFo5gLaX81rEsz51nmJzxhC
h7rDXiN7qpIC5JshjJn9/xdWzCAGE6x6XvC13jUdsqlUU/jXqiF+6Tcd/03MZmzgDjIbpeOQ5rtU
6m8IS/9YLqmdyhienQgvIz7UuVUzYxNX3+kX3TsboS6juq33kN9WnNnRGcCWpqddKbvVYfyMCuSS
T0zB33jF1tdTZz4VAr5Fuak7lcxXvnvuUcYkW1/WgPkCt8V2K3LbTOv08A5h2dj+5fETNhXbx4Ug
ua60uoN3Lst5V/7J0VobBMT/epklpz0YsiL9kASbDHFLQik0jbEdgS39ZEdmY3N/lVB5Wj6DYWOE
S+kjHuX411j2yggxgf7S9OU0bisQtDIN/grrmgtAoz9wfjQpNwvUrM0QOLzpne3ginKNLTRYo/Q8
gHG2YMb4e//PCqwx+pgE/3gx6S/IBK47dRu61/N/lrETdaj3/+iSLEPffz7uCdmQkmIEh5XL14sH
cuNlDR2IjM9WuZ0O00IuY5rHmH/omqtKUzgkxHqeLU3r3TvsV3TuLxEgzYeNMg9xz5Aab0l2fxqr
zX3IrcVAVWxSxNGM2nNkJr5zuZNDlr0LNKtSiY7dzEiSjY7Ut2+n4OTvV7wQfOgpaszxDPcKjE+8
k7cHBH4Yrt70+o/1y//lM542e+6EGY1CSQn234crmNt6nrRL2PZX9id+iHyqjbPBS8dJr92ZrG4R
P9LqwJd91NeVLQOOuLK5AN0Zb0VRemAg+3JH05w3tOQ5z1wYrYxuumlQ4KNffpqBJtqTvvZtC54Y
lHzMBaEGaQveO3VpLS99vltd8Pw8EPWr9KLw5C1j+JqPzC7tNxECcyG4zIdQXVo52YS4evSUkgH7
ru1MSDuZ6UvZN9n27ON3yJ22s+KuSS6yl3kkPeL+YqULV8UYX69awD8Dgdl1v+8TCwQutUdjDvG2
xII7O3B8o2jS/0J3ocT4spsZ72chjJAc1MQGozb2Vm5J4feU+5t1dxLBHYaaq8I5Nt4aVIt73O5t
prGfpEJrRBBFuFP4UmpPIb2KTkfDyxHqSrMxuc3/7R7PAbzICT9OEpeXksgoZrN/80zNF5SP3XCr
HKc4YV8C2VQlc2LrPk00zheY8b8zRvU8S/UGvKwU77OEENrtSgBeCCn80ChQs54eI1MDnt3EuSDT
KdHUnb5sZykrKnJglTyDl/ma3YJsKz537cWps/HgLsoFgyFIXhTDwqqFEFgPahlCzHVaHdW9gaV9
ZPGJjKOmD6MuNIt/yA7uzcmXi6j8aMLuTZjBMpL0ZlRSgzvuhl4n5SdoqVCNUxL/rJ+Ag5sMbDt7
BQHzrWJFkY4n2GQXDD0lJYv33hFtc6dan9if7idODaoRQwE3BS3HlymgqBiJtLYWDmEMA5ORkLnw
FqmW5SOm8oOsMP9uU6ooB/4L9Te6obZTY6t6IsK42D6jel7UPAUk3v2TW1SNoO33kXYz0fj2KXPf
mlFlT3e/b6iuVuMhH7lPA24aNRSmd6rH41uZk0F9A4jX5gWaVXSmcsXChSRSYDbQEKTxPpe5rqSI
dMt1T3a873trp6X3OdDkM1LFHhHWEBIF4qOr1bcBptLPftZemy7fPT26KJaU6agnxyJApZ1Knqpo
qpMpon09+TCtWnYrgkTohpQqCxEKC3VOlTzJPfsVqHnXHNuFepTGMJhFIYCNEbxGj3AlD+D4+Vk0
HCKNh6ByXPNOGlDEazGEDyG6LGLVmv4TSgGA4yX41ociSMyUitt0ecnN9RTyTHiwP2ptx1idLbSM
NztAx0HlFpCF0fMlynYfaE+L5Wi3nw3kGJ2dODqvaL2kEJ3E3KZB9Af465JfNg5WRf5eXIxvQk8k
t+/yOBIDo+GOeGJ60q1PYAcFqe/eFWCAzGRYVbM6Zdhua23dYdS1Co5tN4yGofXbG+lxufHd0kkW
Ll8xdxOMR1nX0DDnpYo1InKjoNxMaJ6uho3PV+PVaN5EOfL2AKz5G3VMrwFdRW3I5TB4kzWcyqSG
AP9FuOXwty7uBOC+++e+ZezoP9naKpgrptPep1qPRutvKdZWTFexNo88b+CuzrC0/tQvzgyWuaKx
YE7q+kFTaA2e6i2InHLZe7alUWu5plHv+1cq9Vppz6jxw455hlqkRs9FteUNyU1p78zmrzpAqhXZ
LdVMcIBTS0B13NJ7YjhFwy3gpOGSWmzyOumyEYnUmIYg1rZpJe6jpPckRfmRcZZ4SKVWU5bwreS/
5PU8YEvZNIeWPV/Xz9NVRBZSU4nRj7sUnK9EUx6okxkfw4ZAQNSgB7b7yGFuBiv0o+4oS9oBFvce
wDwZWh6ID52e4SsBnFL/vZOooeBBIi4aGzlfjipzTbDBB5PKk/ZfrnV9eADrvzueDU9I15LMDcCH
I6dnrPDDg9U4rKtN+MqaaxmyZ8D+/d8x2LeogVUErKco7VLwHsNKK3u7YrTr0zzJor0wFbNCTmo9
3VyYLhZfpPakgxRYFZWZhFlGHgqBp2RBblC36WTpUcZNzc0vj6l8i/CW9SfMYP0YDS1AjnmWkyB6
W/yMlNHhZd4iS/OD0vhcv8aisanJ+ggMb8Nt9y8gtGXGmZT3T5c5ALtKBUfjOP/qijAe2z3vjP9s
P4XQfZolciuiqd5HkPoSs3AOGbI4xkKBn8A4g/7UanpKStjmgh5sFXJj6+jXd21jqgeLkIVf5quI
fwOouSzhHIrmMq9CZUrIxocvYBeC+ML9mvqHcGc9w/bwn07WNn8UYIn0Pf3+4IUNG2aaXtSvPnnM
4N3KO2MGr1VSMtFcr63ZdYvqhKt/Kge7zjp7WS9qCeno3x2tvi+MshPrgl5HeN+Zvkn9GjQlPCWg
7d/DFwlva7KacPKwj6PMpB1+WdQ+AhDoktBBZIyj24J6Zdq2Yrkauq3j4rRm8xOFGpX1LLN0pD+k
08mFRDZUMJe1u6pkJfEc+pClqmD4hHLIYcnReYwOBv4poo7HvHXcPFIUgLx3JzVt91EXBEAdvuRi
db4q4JGAe+LtjXf8pO/NmzSBDL4SH4Od7mG991dGaOUL33acy7Mqvf+bD4fq+CbrrcA3pAvo3cPL
we0t7ObVSwSq1s275fPzizxtURI7++IFb/9XEZqXl0+tE7typbrVJTtmDIVtko19PK941lFZ0E0x
TF9T/0QhLnPdsstfVZF6s3cCuatAKxk5JTu6CbQGR15WGKCtviYpTYRzEaLpM5V2PQpPYwlEjYkc
H08xiYCLgo2zBTaS+PbwH6h6gkYdmcElCeh9xlzpAaEhvJERsg1/t/sb4ZTFW0fDwNaIqCLhbSjt
6WkNO2walKC1jN1XBjXAhZ++sBI8GSFIJqoPfZzn7Y2q++NevjMaXGCf8ASAmW46w7al4XpEnKPC
StyCuu0crq2rf8dHYAcce4AIY1RpVSDHExes/eMF8x+m4VxmUtwNGhWqNvQeCxqXMNFIYxSR497y
s744U7d5EXl92IBzRPJpYDCp5/Mi7O45RVOKjpa8NStucFSf1PqPBagAaoqf8e6Wp1Q91scf3aKd
dwo28V+ZGQ7TRR8LBhXIcC5iKorLUVtoZZPchDaczqwCEIz/E9BVKkix/QyWXNJP8AcQ/x9umr2z
Djq5+g4pmjK0pUV45P4aZlKyOziUaknpXLQw1wPEVEESjmVNmrHlmdToW+2nwyDbJ56/zqn7Tdna
PdX4V4wbakvDeqzYjFGlXnFe5mJnjCkSF0AaAWKbuBAJM2Xc840LzDmQmAS5PivJCT4x7frISYPH
yOgEsK6fWAZOjECnHPnLYoKybmmf7b/1KtDGyjRU5tf1Aw9zL1v+UXjULqwUwQNBD8mZ5+Tm9imj
OMMShj3aTp8YSb1nNOf4RUGE2yl1pcouYlzVAsIa7b1s35hQ5DctaPxE0x0sQNkrLhuTtIsBKkpV
mXreJcWHG6yEwW1ziXd7YkiU71WxVyIq2+Vgiblgmr1GTG9mYey8NCs9YM7QguFLlZFw2LmxdBlE
U+fTw6pQZOoEi991PAl5MQQGu8II886P+7dhcXuiIxn9KCXD8OJnj0Njo3rJQLPT667WOh38DetG
JoqdsuwDgp1qcAYEom9IlW+Nsc4YFX8qByFXZNXFPEgsURDL8qi79gk0NnK9F3Ws4mii8+khs/v3
cJNsQklkuYFNOkk9Bajwp1HDUNu3gcOSVnWhwvjGG8u7IiE6IgWg3/3xi1gfXTndm0knVUB36/UL
yo6k3DtyzXhDz8seKHTUM562y6fArvDrtz24D73IauxQdxJ95hdszsUfj13MQ9VGfIw/v25O/NVK
p7dgyLGlfOw4C61oK5VU6SHK2pln6vrKd43YeG09rCp7OCdNh6tP+c4klor2hHkYzGEcJeLdAhjQ
zEYXg+Zfl8G52FzwMre+6Ob+D0pKjRydf282cyDOA/xOz7ugO1JCXPSOwbX8PBa1Q4/KboRY4PY2
BBRzBu2i5k9/4Zq9g+wkDKOmG7wRBC78+LghPnmbyVZXgNwpMptZ2KIyEVbhazoUg2mtb+aekOSm
r5dUJRrEc5f7COu/SQt55MgSHzLI0lD3r9OjAW/g09Z+kuF78M0SytwPtfj/VDkCyYtW8C8wSogB
l+lDB2lDIqbaK3lQfy0Gab3xsQ+ugMlzi7mUPLjRgZFgjpH+eWKWoPtpSaHFiS9PLvt3C8VT+rPj
aFU96Sr8zDYaFMY35d1c7UYxL9bNFFmQg03pQRrvukXZQvRB3DcIftUCiiDY0D/bgWDAgCXUEdin
uZDlI1hFc19neobISnly9mFHq19AMcCDnE4iqkaXHF7cNYyyRtdev3HzZlsx2I83zouH2+LXWXNk
arh9CLjN3R3gA4bwgrDEUsBof7CG9SVMWy1S309/GaxgingO06EAhJeeFFi5QpUQNEWPMrAE0CRZ
RvNpoTA9x5IEyq9Yx+C8FN4h0Z3FDHhoHrscDlU0GkdOjC86jsbCLUvfPpGIFVOuPXIyQjbAdHVT
jql9VlZpsGWixLUTluBgUWZP+1NsWapUpfGKPgwx5nftLxtsd6LjpqFev0w3j7sM6u+R/OXLI/Rp
budil584R3JFpm3SxZT0XeVt2Sz74StekeYm1BLTOtImWO+yjHk8pb4doAzc6hL68uSQbi4OzpRJ
2BdwSBtf9KgB4JTnYNkScf+kPvwfj3hu8tuXBBSXzIS3qBvSvkf4kfF2GIO6683DZT2BOChVlhzs
1kUh3gvM5hEVjAbUwDAl88hoUAxmPAAQWWtDkZ8TAzPWIB4ib1KoOEafH+P2X8x/zniTdvn+qjUc
llFBxU9qk9htJKzjoDwvLPFL7pSWa3WWqvrapSv/5U987WPNhtz3U91vRcTwopcLRAImZ/xjlciQ
RRV3M1FWwfJsWIGnXZD2Gt3jTlzjN0MXx9lVxMgS5d8m3yEROEE3htu9uc9CysWMBM4+6mvn2+vl
sc2QpaM4xqPiT+XPTlz+holpdqG/HfSMLNYV46rGrt5m+Ll9qs44dAguXeMKDQhHxRLd42vCGd8N
rLaf4DOnb4B3a9hnsVW8EhQCz6e61i00Ovjjlw1Kgabfzd6MIWCPI/8FzwRWRMRzTH3NTiq7DNFn
A4co72wz0rSHLrAMpyl1y1c2C+Xu8HcHYLmqbU+9L++c3zOssfrAM/xXXVW5JZxJ3s5kpm/zxsxi
c2OXLUcTO5kYmz8mZNOIElcZLuQoIiH5BSfNzKvHArK9APqUR6Scxe9l4YD4P+dXvUdlmr+JSQr1
gwSJEr6XXJO4deHMSYq276jg8b8HvZnQcNaY4Ap/vYZDjykFgMflKq8dXLvknqeQqs6uvG8o+5L/
HSNdFIolV4zou39DGLvBrMwWOHurUTlvNcZUAthz07g1bLAfi1S43gHFsZs7r2+l10Y7XkqR7nUC
K3pgFcw2fQrtWwJwnIm6YGFaiwaZQYoLPfWmugqIAbQ+mvYdDFvOaLjgZatF/njenNoVEOrJO1aI
OcfeDI2RiGAHkbypNFvNd+EEfDOkvEGUXlmZUefSU6nWiICqTBuzD6xORoj/WfaoapJuGDuus0MN
w0D/uqUsSq65+uBd1RiLWcC4XILdJ4vqtNNY0CpMqZtgIn2h1gCp+4lM4u0h/Oah5YIJ0WYkQHrG
favNhOLrOMdKoAihwk1FchWtuQvJ/WRYlG5t7P/2kSYq9+SIo3dC3ZCCw62xAzT+QYrxNcPXm+pB
ptNzOqzTzpDqA30Fd+9CndS16p8T2ffeVREKBhGhibIbTTo4ytn9DFCQwddo0J04QfuUwvFALifT
ENFYKk96x5ribonOCkrOw6+mVFvwqoKNUORSba8X5oEGkhKhcOSQzAnIos2OZTUh6KIswtB4f4sN
I7OWLm4ypWqWf/cEmLqj/Dk3QNO2l+/84wnbiQw8KLr8TUsBFgorFD1LIArlk3+J5Oyz9S7UFksS
S/mRKVNsC65X+kxUXGBkPblg4xkPAIbAhJeepgkHj369VubKRpVQOi9oaheAm39LTbTzbcPjb7W+
+qX4IiTgt9f5HNQQ4E3JccfOvYKyITtWEKAizeH7vrHDC+y18sqeAnJYZLf3s8KUePGXzVFyBwGu
oIbi4vqQYbtj7efoXeM5BmuuNSnnR2RoSNnFIS6wrvOKNCAZFkKnFsAsVr6jiqjpqK9Vf+KkT1hw
8piI0PE5z2JFhWryAc4PjOBiBPiTKXhYLjg/ccSc+Y1Ogjj/XR3fZjPgbMMAMlGfN8Z+l/VEorXf
ZUARV/vw0dzm4ZxqUB6LaKc4IsXA0e7kl8RtCAHaCdC7Nk4e5wY/knvL3kftr2MAO80tSSNvRm12
tzXB/3qq77h8INCL4r5BAlE+ZbM6iQKwKqfN+tFhwQkKb9jkV0vGFbsxIqsOfv0/UoDFTkw7tQF4
+GkIZSHlS5YUXHCgvn+dalOqCYD39d4KObH7nD43hPcCGH/U1h2THATP6l2iZ4oj9E3k6PLCB8L7
zSV5zDOsFq0gd2vnJQ6psKJKRmHbYdUX64VLUNXhHy2DMhKRp9EBn+RYkZszwgIWezWBAIYdprlI
x9I2WDaMWrcZY+1s7pHrrnJiASRYHflcb995Cuhvw0ukiX+a6vSg1I2spzamy5GhMZyeJ3ksV956
ndAGWYPs5x/a7CSBPrUTLk1YFJztXwX8ZI3cPSFYnm5IPaCpwwPVxzHZ/a5/ZH7N7aAWoT/EKYBA
0pcQ6Huov6tvrpit+5jk/mD1ATb9W4K7rj5ure0PpaJPtoxKAPj35sAPf7b/HCtSp7ld1Czc0T4O
iJRAn5Iqb77raGBUmrpjDlO8Q7mmfQGn5gT8EySzd0Y3Qw9yaOukzMQ51P5CC2WxEAx8JqoBtiH0
WgbPNZARjlIvwv1HsjxQbgfegEzNRX9thD7iKsqy5ifKFuY75qwffJoZ4q6EpG47LTefUc+dNHnS
XDL/YnmHzRNAd7po8RTInKlAJipD8MEKaX5xq1s4CKjgpWWMMBiWpwE+4CMPfTO1A5JFTlgSFqXH
S9xrPI1JuL1lIDFKqcM+NEc9rzaT5fNyEnFRXuPr+olOsl0jk094WEaWZiqWdh5rZlADzSrrBYRr
nJtM7vwOHJ7czDpeBt/WVStS3R8sf+o62JXH7Uj9gduUkSjaT3q49veYAyZwLNIh50sr11s/fjDL
txpMMzTl7KHEcsdRW4RTMxNENbhy1ACpIwQdG8S1TUZFVuPY/A7mSKtqjZgJRDVGZ+TI/m6BjNcv
bSvyNwhQAD8CHhGy2zT39axVyIDG+06Mgx0J8/vEeYBDkkOVrilICfctyqkjiu2s+v9e7WIYgeKi
lx4PVNQkGP0LQHsKaf52CS68q8V42PQGR9xMt3+l47/igR6RnjljDmpiOFsvT/wCsAbV063AydLi
MbdovfR15JVKevJS7ctvHLqjd/Fdb6meW7nNVsQL435HzF2U14UmnDS4XJYwIP+hIhVCcXBr6MsS
j6fvk2yKCOY7VcmyDUmQgI+tGd3cxIezV54k9sKQCVdvPzFN+qSmR5fUoLazsw2LWA2FlZyiXPnR
ZIFXjyn3LByw5HprH2WLvOLz71kCMs2McmSgBpoHZJiC5TNXru/AHW/9TTFVTLisgOoI0NZz/MeX
a7n6Roz5uYLF8RdHlSYWDhPu41snx8wrkBMbBJpZs8VBhtnGZbhsPYlxzQvpd8gBg/6s1Cf+Eek6
g/noHd3b+KqlRikJWyXWdSRq8debfGMetxCYZhHvEYvm8UBqzluVBHUWnxhyzGJ+4pUbsmDYDl9i
daEX3TcSMcUfkonUTMp/TlSnxKD1p+cYFOhjXlM0gvHbu34qaQfCqpy9x2n04GQSwutpvSdBlsVa
2Wgo4cBVHStzmY0NZxZKWWnlF7PiHq8f7nWYMVQIB7Gm/V68tRRJabE03WcOZDjlJuuMGeH/MOMM
m4Kkpcrmz/ets+/4ubFDZdiQbeOZHpOPBQR7huz9UyH8WDb+qe2Qi4JzXb74ZqndU/udUPFQwwNH
lcQL7tDlhxRUSX5kYTKpAaktFkkjw+mlLOHoa2XM2EjE1BLJ9tesPomiFRH3t+siLjvob1hIDmwB
zUfzVOFrZY8bi3Sx515K7m4I54sINfCMkAsM0qRBExXXffBqnHGRnCCDfyfCW3CwHwhPBkxAEJbV
Gm6HyVLOt7nuJC0uIT5ewMzyDKjkabubqT5kaDDea9byAZgO5KCmtaf5EpPTA8wPFzBrbMIk4Vgd
XAANWKGDMAI5+AoHMfhmTnUvANpXSILAUCBwaMmLhYx5HrFt7ADUPJuG9TDw3JKSr7IvCDjhqZcs
WOaaNtd97vs6pLHFIDZK9pV6N+/P4nqIi1qQc4QRR3G4hSuT3LYPgp4iptgsK3Tp7kZbYGxO1jPR
ha6bdXcM9ubIV24/K5OoxHoXwls1fYbaa1S28iFj5o4nPWg7Zj7L1Vaq1+DChPHdoOyWWRkwhlD5
G1r+jc+8d9Ln+/YF8+KIhK6ucwYd9tsvwcJfvHwin4+Qt5cADKRVhGA14Mece/EDcD3K/Wfy9B76
v3MGa0dNWtX+wQeNp1XZl/28O+zTX0c7RyLZA7eRE9pGlxied1YS8agSGAxA+iXoJETRT47sUkie
UHW0utiipq7DjorDgZg9ltqnHSv6dBcC2aqn+9KbtDUnOQ4WBVTs/NFk8SEOyk3whJy+v+h02diN
6MzPEPoz7rUsARJyCF6WPV8CsRTHGQMNMuQZfNICdW8kFHuh59AgtGYC6nLNBbRF8tFSDziAHEpe
yYwE6LPdCL+okzlXde632B6b/cEAQPd4luHoTDOyDlkfokp3pEnZCFhvUZoLQjw2mPJZCCRK9YYU
vC44zKtD5nBthlTMIq3TmCHxxP1em8ipnGyfDWim0+DwyptYSs1rq3F7EPn/g2VlGsHDj9FKb1EG
u9tTlKrlHKR0hKP4jUpXQ9KkymgitBSGHGt02tJCJymzgjlnLsCjHEaFzRJ6nRH7/36/zcQSZua6
RWwUJhJ+gHb89CNUhMh6OLd0zbJ9GYYio8AleHyVQXAUEAi4Rjt039WkxM8LjMyXV7LXW0UT8MTy
a6CWaskUuSBvHq0c06adIYoLGm23IhmSpGAzA1Ygy6x3KaVzwp/Jy828forzruEt0z3HNdfmOpAl
Vq4Aor7kaMLiUpC33fY/nqtLyU46OobINA4L1xt4+qCgI1ZWyruAscJTg20YkPZGRt8Fb1Xq2zFm
w1q5RWP/nR/Wkmglm3CvwKSBCEd9VKolmFiPW2oamvwQRAi6yEYXzcCYgMYG7/YvJXW5sDAJGpb6
N2C77k3sqQulNcgnD/4cctZqoJQFjpyjLerlUaTh0jFcOQxWUN+06H6diYGMWpsTSUcaXGwqWT0h
cQa2oMqOeDHcVn2QLtnelaeAX95z1sQa5V1yoB+tSTZPRMbxA26IS382Um60eX7PYhRNRSRJaIwx
Z0RXV2RRB/fvBD2id2sMcpZQyWhJ80uD3kCULAGykey2wdw6TKMbfzdIWW0WqQLwbg6Nxg9iB7QK
bAJQH3RTQiyCN2vrmZH1OFWJuq8jBVS/lpL/xVqBZo73lDZf2WJDQvk7eXi6mvRJrQWSDJP1EzTr
QoY4umgzckv3FRmi43HNTgJEaaFhMHggxe1HHqh4mmGzS5kgA9oVMNiVP1KmXPe/WGVeL443oWCM
jGxIk08dbTQskiLBlPjW15IG9wpdYOHxHyxxnQiVHER3vs3+P1G1TBX+jFC/PTbw/AXfyQQC6WEl
HnVYyutbk+uB0SmiTcw+7Vc2wzCt3k2x2OqFuMagoOQUUDoaM1bubzDC47YJAIgvxZFcEgfT/X6P
vH79cJKi7wHQ6jyGzZ1jYqobT2cyNwrsvC5cpX2wIKDKmG9f9XfJBisVF74Z8q9Rwb3b/imcLu+r
6BD94yUrerlrmxptNIkt9C+Db0qI/Rvajsa9vFUaJsAOZ8+gRE3d3SCx/tva8EYFFT4oeQ60/pAT
1U9JEw7g2X+2XjVgs+j41ftIYhMg5hg+YopTtCu90FKY35s2kL5HMLeTqejXI/llqZZILdgJ/W0G
cFqsX6sl6HG0o1nFSpb1fLi9A401736MXs8xq1/T2yJ8yfKjyxDi+Y+vJ/Zz+iP0SjeryRXK5VM+
PaCZzgCbQ93GOna6nx2GImy90ybuQbeVHPVoTqsoiVVfyGyBFaO2t4meIhbQN0bTug3/5/eGT0V5
asx1AqwUzYWRIHC8UhfwFYPx0Zqqm+yXHqzkXu10+B9jizxfpT8idkz3oDDqcEcqM+sxOoRRurLH
wJVEpNGy5E0J4dZDxj8iuG2NfTmZj/LAbz901uWgqjcAJ23G2WyPFNpmO2EswoT7cZN51e62XhAR
3ew6GHmujF0Gh/zZtgqVUsj5dBBC0XJ5DUw2UIFFKBpHSSKnfNIUOmKxRMZIlKICy4F5Yn9uMLkz
Dbz9zGGyQ6ggdT5Jq/cZOgs/FcLlOQoBuETA29KEq14fEkPEocmwKij7E+AN5fRjPWLocWZsdhpr
gcpHSP5WX8VrA9d0X2ThfexXWEVa9x7PYwYlT4ZwypKKt4KGJsI3/LDSSJTvNtXJlwkzXtw6fNxN
v1OKT7taOB+4D6W+d1YCvIPRUb4eQscoxNCPiWaZqv2SU4a504WYIeh9fB1sOkBlr8ImmN4xd68K
zL/aA/MZD22YTMNj2xJNmp7mw2rY4P4ZfUDZpPvpoWFa1rygdVzbxpOMX48jIyrXfub32a+vb0my
r74Pr3zrw4rJUdbGQ8ahQQkbnZUk/zNYP3k6fQrdw/QdIr/ZGTh4uj56TEJFAxtjNV3s0nVB9VBG
bhjBX8yLo5otveJqan2NHbcBTAf4zFJRc1eCRHoz94v5OL1Y+lwIB2BiYWfuJEqP/0ErHfhwUUxU
TxA2NVthZgIBSdzMTb0IGQgPI6xc/IbxWV6BAfDX9sZiIxK3JRE05tdq3JNyoRijZK5Xu7DH3Goe
gNRbRTdj700QB1v7Cu84JAu3MRr32O+78+VZLmXlfWF2ry1CEcmXLkSYf8jQ5sk8jnku7IGJYpKa
T25akGvNKbW4i3qOwSYTVcZhStoTXAJojZlHBGOr+5+q8eXt7NxMDuhV8eScPx5gco+xw5kso3sG
uENlCHnZ03YFOuUSySDxO2IQovymq7iGug4Wf4MbbXor2mJvdnhbWoyoIvegcXFntv2+COutOLzL
ysVF+aAlW0Tf2Nu6ShLKDcSh9ZxfhwguFqpsQGpzuAxZyONHUO+mlByjMhXHCBCrL+F6UwXqEvf/
KCnH61rch240pTHkAr42lzukGxBm5k/faenIbejUNHk4m0mPXr2Pb5dN1qMy6sUe6IXXjr6hOolU
N5WeYLkuyPuFmNnpdLB4uxBNxlDH66YyiicFMy3BS4979YQI7MsZuT/AkzhT/77fAS2VZ8qvbh7Z
xm1RGNsPvrvU7oUIXkwYe5hh6or6TuOjeckegCcQPAiAk8j+uUMGtYN/E3xvMojYtNEfKzt+sB7R
SrfSjbdGxuapwDMBQ8aKFAPFacOE5AZlTweOZE48qTv595UOneaVT8bE+pujXs+5OotLZey4lHhx
BKiZW5aoIG0JeJixSKruqQWza2AEO+TLdACmDg5hBVZ127D89/gx5V2e7s/RaiAITAK3RzX9Av5j
mXk2B1vgmkrzvNbNM1ErAC7XUaqc+qeYSpN8edhNTa5kSJ77SGtVdGGbQ2MQkr3xcjqYYAPVyr5x
3hHSfjHJa78128d4KtmOSNOyHcCBL0JB/GjE1CxG7JbH3qQCiL8wwrTus0i4H03xsQBlusGHqZba
HodAUq24e7S2F2rsfKrbnvnfPLBVIOAJl4QXhpkpRBJ9tHijBzQ70MhQFLgR14kL0Z++hbOao18e
K656q0O2S2oMFNsqQQ50bJUD6WHDPydQqOrGY1dbwLloP1bzl+t5p8EJLVPXgPCIC7p9cj7Cr0K7
iQ9fbD+/BrIRWVlkrsh4NwGzZI101IPgiSQgDvAqzEWXbbVauf8nJNx3dykN3pzB5afUjTjNXdAn
xheRVhsBzbdDGD8sfHKDcPg/3MPLF1CPFxuhDRzzqZFjfx614ffrmmHBtcC5bTd6/Jjpw/jp4dUu
bun67xfw3FP9C3H3ak3RvTwkfXZz/3jxdyhNvqaXdKuUSAt8CdEsIm0zMxcITCAvll18SxUFLg/h
G1G8/Znxa0/F+beJajAl2wyJarGhPY/xCH/uuINNsz6lGbto1KeG7zmdq7kF3VFx1iIdZED0VPgo
Wcve4/WKpRWs8t4o5Rcr0Trk0iTszOKUWWLLTAYxSOMBrmfTjO6Wvpo0/kkQ+jUFV8tw56ADaRJW
YcbK6rgu9pyhc1oewY33TwyuRTaeX0mHI8xm0tS4Jwue2Xen+lL6VPjZ4fe6RRkxnKOis8z/345p
bMudLwVOzoQgwTWwct21uR5TIyRaO3R8xfb+6C654SLUT0GYmni9oQPdmMTGtIxBPuXrcNzEIWkJ
udusxO7IGzQEYBxOm3/WsY4wnaSMlBGe+Xmoof1BjHog2VrJkmo90fQeuhI4SGhEgqVz/8Etxphq
6CHA0hNTuC3JOVY1hGKGxo4xam8dvcBzus6eXfsoDh+T2R0OZ0kc4KwEB0wYmOywe2Fe5oBNzywp
BmbB6xrF+117lh3yAIo1EndEKamb+EV3TWR5E6p5zQ+3M5c9qJywImbqa8Wii3Le8QWa1Bt64jfO
04fpf05pQ0Qs+o0xOGkddjZpKDXFaqrVQJ2sdgrU9630HIG4xVofox0rhRnlqG3M1/KZ8j/riKtF
uukG6Bkqq85bxFV/L3Tgyq7uyBBKvo79AHrely6XQAUURiWmqBRMWPVqMR1cNIdUdEChptLyxBFF
V6iw+nY93nHSnliTCjCvDJJSTMjWTIS+L4B3PZ1O9gkwQEvneFdx38ScMR2uQ44q0oIE6HsV71c4
fpiAiYzgPKa9Ab4HGu3E7CfdzcYiH09BuBSBQy+QfGwYOOhs+AtEE3zQH/mVXsc+giUgesA94ClW
ADARQ4W7Az9CUHIHdan5PB4C7dCq3YKTCSzPdxH5xKT4YO/KtySPlcy3ADsBgnIUB1pawuX7Oyt1
RMxaFPfl1E0gNODn08rmRfsxd5PJofe3/MESSnqOi7/Yv74OzvR15Ce4mB+YleEjIm0kOJNQI3jf
klofk/zyfLNbc7/us220UGZ0FgwmFDGCroHk6iKEDwyBg5jsgXlGFJBrZhXPh689zlGeVdL/XLvY
tgUzJlOLc5RcxCFSOva0gllwCI7Yr97eAeiq6u9r90OIpvt7+rLsmv6fsPiBNUo1Muhz+a0BESZK
ID4ljnUwV5Lt76WcKPSxN7zPzojXMBWRMk6GfHlGI8JZ1STFrbZgckU5r0Wg0sGJ2m/aCHhfD5M8
9fyPadbDm15fhm4ZkAjrICE06UGRoFwTbyvOCYVfD1Dt/qnlaasw9T69SEceMRlbmwwbptQ8jhK/
Pn5IicKVfEOhRCj0tgz3r6v3OICOpdWhwYwzgv0T98lPp0YJC1EG6MS1+DxfNv+/UQTy9Iw60CX6
vyIebfWy/rWsKTfLd39FiPnQQmZjwXBSUK0G50DJQ7GySb0EZ9WVtyDZCC7zDKaiS5YgOpTj9hAq
RqewJln702M7YAn9BN5j5vI31MPTPqWQzR2IVeO9fQfnM5MEhuztlVj3Biel4NhartACXorK8DUH
IYySVjpIKWR9M4uPZ+opHDAz9zuwwcFpXfh+Q8ruVxjJ1W4eo7UdevOBviAUfxwik+FUX14mjLde
G3dsoTuxEqpS6RX908LYbo9vB9w7MiXEWskL6P3pHUzQmRCE4qU2l9Slbh1+XP6fhCyZWGkCY2ZU
1pUvd2iCa8+XHTd/WGtiVCLhw2bR1+jNZi1YuC3pUyeZdRQLQ6y8SbUCsjDJD8HjvEGrcUH/DYIP
T3wv2oeQMaJDeFsg9OvA5E7sbIGlRO9y6owhzZ4n7nJnz0qcdJ97aBU11DJ9HjeLdVUao00G1gcO
qr4T1A2sRla4WFgqqFBEqMCubw4rek+3LQk2sTIym3QYVtRuNjn3fTbbyogblLiczHdeoxowGUFr
0iiQw1afc7Z3QLfFeACyHmxWMMRVIkRVMcrflaV8RvrQm19R8O91EE842yWgQ0POqANOwQ+rEogW
TP5SxYzbpw6Sv/QCJ1tUxuYqHrXPmIaESiO7aer/p3ktUyVptroLF2ukPh0gKyJN3j3P5aq5a4sw
qMoic09rfEJwllaprs/qe9v7O8t7S13/vBkxH9BG2dZxYT9Zr5ILPoOJw7RgJoaCCxaUqysICUBb
bvXTAJb4I7NvWtJCBYajn6Gyzbfuw3yWUVsbU7cnv/7j1KgsPZvOQO1xwNKQlZqThpXNnh+5P1D1
aUpuy+NuET1l1JU6VapIdJPfx6L7E4idRHxxOT4BFEXKVXibMi9QrxRh/xnHkG22NKpw9dqrtbPQ
8GohQd9PbvEHcuJVSgHHiLaB/c+2Y5ksPJl+IUg0tQ/0AuE4ty8MhF1QyZh45W/ae3lHerwlPhNq
hCMeGD5rkEZCxsPiSer9USciVvWBh8QNILBfvuV4bg08M3xf+1sP3NUj1m2sjzNG5TrBRJ6pLYce
Z3xsXfNFwZnB62TGn1oN9BnngEyQ6sN0eCDkghOx/oS100XGcpB8lX7hCavkNd3ar/pKrDevyjaA
stNOgUhoPU1WfuC7pmo96mz1YBK3Y8966FOOImOVnWBYh8ljIRDgZCZEXjObGv3uGVOgJafea7W1
Sq4J1QBgzjJW4viSku0uT0BBfqP1ebfdcoj9RSJVYGh7AXRTXsqXMzLZRWC0KtRLDkP3xd0ozFcI
VW87hY6SEcK0pxv5ve1bp2Iry2X1TQJhs6l6GNWNJw9v2qL8TWwPA7WkNcmMd1F76cYXDa1SKaLH
lVnfR6sbikM0QQVFJKWgo8ppAq00xkxMayzChnGbkZsHj7nM3hl2gz26fpkEijfVJSOQGo5EIPkV
V+pgSoFknyG9XAvkg8/dWf5zKkSsmmpW27ggcf8UkJCDG6BXeLnIdSuAz5U5q9NOxzKSse6NN0ex
LhQwHyFedDr9Os/cEwMYxXNX5dvflwjfkL56vN2kzb1qkecu84UlV/6yOr6fXVoSXIxfYc1uc9Qa
8Pa06ZeKKNRhloMVdvnOgS/+7+7zQL90EfBM85fEXf6TwGLW0OH0TLw/CPrg8PvCGHUfj6OrreZa
19c30Kx2cSEQ+Y7hPFU7k9wFtL/I8VNZl8P4LCBAEHk4JOKHjdeiets57JzmRCRLcBboPa62+l2Y
dncRWk0J5/Wy19RVP/SMoobFBW/SnXU6bxiKTIBvynJkQEolD5f5wnCTx8kUkAPxBHC0swHayCOQ
K9ecy90bRGCnnNzTT3dVBf73ht2zhK2TuA+ezXVTaLxI1yzKW5XjiZ4M7BG6VEVQorWIDX3+6yER
LIlAd9CwfPEar/Dek0Fh7wen1IeZuHdBP0qRP+dK3O5AMe4LLK41XQpzXaGgBGSuxHLJuJeSZtWR
wn0kObsJOMjjpP84Vurug4ceIY5BCJJMxahxDffXGpovrXN5n4qRpP5QaW0vLnfAL7PWpn6jWGCc
gf+VOoauxesm5ouSvHRFukH00KtdrIvkGQd4pxxFsjpupNU8ozJOM+InJRQjRRBog6Zi2XyiztKm
IsAoqhzHSjupAinfj/Omn+4Ld2LepEeLMCnvbLod01Q4HyaUdn9l/DfVfjJ012zBLwDd+VXsttbo
t1po1jzKsNxCLK+E4sKzVWuVuBiljvGjvn8BryevnIwJGHupcw+9KgBGiZMQ2HfPuho0N+JpBSuC
i4iSArCRGQMNhYuDhX2jd5DWftEt/b4vexSQsXWlK/sPy7lioUXHajsAMy8KEYpWLlyU1/oVYMbD
WKj7JGtBrT/dVmUxMJGVK3ZB/WOoNHMH4w/4Z43cTcIz7pugTvPpbmrRb5hNxIjWjLSyE87xKYyc
wUtfVQssgJ9I6J+VdtS2MkuyWI9zeF/je9YIjMO2ckirhtQntQKPze6O5CYuVlITssRNEW89dH6u
376CoPUg1RPJGKutXJQDsEQq47wH76elGDlq1wXPZVZ7afpMM+DHA6Jy0/eWcilKFYLOVNDaJsmD
/22k7sBKTYjA8j/YBHu7ngzaAB0a1Ur0brXYMII/InpTaaKwjjQLCQrlko1diSnK1WUaeJWhaxOq
SbuYSBKSW7hTaG5UlE/wxmeOuXbU0S7g/A2lCSDr3nBjDSwYx+9qvlrXgwwoRKHkzr75RX9879Mo
yTqu193q2LwyMakuPIgRtJoPAJdP38nqo+eYc9NZ86T7Dgz+jMBUi2eYqiS0IKWMR+pcEUeIiOBH
vpwDWBzDWPiUBlsSaBxeP+EidclCV6OBwKNZIbCcVnblIt/nJl2b5oxsVjrS9HZwzXWWKKSC6gWH
YGlCzwS7R/R6f2pVMGUC0DVT1A5fRial4kWIpTTB10YB8e1U+tQoa759lc+TEDTzKCVhGG2p1GEG
oNacJTGsOSs3wPpYutIseP5wRjV6SrOxCLu4/IWWWZ8CjeqFVHTn3crFgjMiJgoQ1lJBqlQG/KB1
3Nda1fTP6UgEEvoKteDbTBBfjiPpjRfC2NiSzc9UkbcWIx75xf9cuhIuA9YypDgwyr3rsuEcs070
94F6R02BjEmwkfHdgXTO95gk4BKe0fjNPXz/fScA8+L/Q+0p96CXh2UJ8Roe1q4GIl5jn0k3qTl6
x35h3fNXKULH2FVDH/PZRSMpiPErl9ZTe2Cre1RvrViePM4oO0Borwk5HKIejeppq5bPxVCbtSTq
qDF5E1yWixOaKOaL4CNJ6NftDvgk4FHfZYp1zo/yN7VOB+Zx+TmcPhpCWqPAv1Hv1dlHg5TU2z04
bdFd6rXCH8xKNXl9NTQqKDwZ06lYBoMvbDwP8pIv2SCc5QCp1eermps73futU/K2k9A3N06HjB5J
nxEytFpgYYKX2MPtQgnx1OLLBpPjbiejNzCNkrtuztfslK1ct//FNNPvpRgbL9ccMCRhzYVkI3vJ
R1mt1cYl7Kl5Hnw9rpnpTbXfuXL2KPYMefIAbLRiQtG1xgArGFICKPnw5VGDmahHrpjcGkP8wZDl
atRV2Nn5vp9krL9uiSYFvBD02yQd/aUUujR7hHPEMZ9Xd4Bm19Ma/ynsRq7QZAlTvf4bpyzZ3tVk
JwXuk222Cx00YyNbe6/C+mIGDjY8b4842hNXLz74OSqrxsZOo9qMHI5VfTK8bk6df/dYkApp5X5d
GpMWrI9KDzRieSoEoouS81Z0Qp/M6e/fMC5zA369IgIw51rDOaK299hsgdAc4i9kCWB7qWn7rOGI
lNiaLKTptVjeWINvwp2TQJpLoA+RuLOMUSZWyQU+w2vzaJlaRLNIIiVqDF/Ais6ym7GCoZNeJieR
GMo7ZtMhtmPW0FqV6RaanmzT3NAqX/+OdwaFP1J8U5o8wBxwZ3yWvFZycvmbJhTmWsp8Mb1dzWgb
uN+igZKRi9Dg2y95Ie07zts19I8IxN8li9kmQ4Ov6O869Yhr4vNOJSSkQlU0Il9ShL4MqdI6Jx5Q
pnJqUrSp7mb67BTAzjAuZ0ubij/tGmdoO6aNYf8NGAYUA8l0y7tX7czt4AK2g8IhUWXj1lUb0Q7b
u08e8GAbkebIA2YrCwSPh/syfZcAzFxbs9hNvHDX+skhSrefH8fDCwqj2IBDJ+uA7g/vOwfTOzTg
LuhYnRZZTyX7UxxaJLPMMbwduEkMxY+GfOjakKOwVmBvIrnRSZUrb3mZF52VfQemeqtoGU5i1QXi
EQWsNkZjRTVPknQ6s+wb5WOxzIsYoHSl7r1aGJ6Qk+D8OH2Px5Hqzd7c4R2nlnoL9WF4Bt2ta1KD
6+SX5MKNf5wFCtJTSKCq4meUxl+ijc/ZWZ1MblnFnmEnMIVg0Uw0qSazg9SCvuNJhUrmhi7XsxDU
juEu/7Ns1R0iTQ6xU+hJ3XSEyrgQ9gjqdPCCgpb49lGJ25sP8UPHBGIrrhaZAop4U+XrCJ65/PQv
H+I30APGfzxSx144RnvRuSEs3bswKRlRTmzAHNCzYADtIKZ/QtLJMbe4RSsnxC/CX1ynPTGNPWH0
OwtklFJWroUvrM8++8XJrrXogeIcuwVx1dPWnu38DKOe85O7Qz15uazXzQp8ojcUTQkNjtwiDL9O
soz3EPALDvjdNhkGjHLKeVYC1LwCxRPKm/yBYznpQViMpONGIdhef3ycxl5a+mKWhZDm1nrNxlnT
8tlAci3GlWqyLqwZmm+e92TCKwCsMKwJAapyFtcE0OZw2M4pSmIyNu2qBF5xEgSAHnQviiXrYaD5
LAMMP8WVi7VzOlXfEjpFKWPihlqDgRWAw5tOXeQykHZXVZwPN5TH+OdtB7hwtksLVhqBYsTYQ+vl
lY6qXYB8WHau98vryKOfb7jxfu/RcXpZ4ueo4N6urUCXF2yahRdl9MHRtcRnu1phg5ey+I2gQfr2
zvYh5anKiPkKRbi0MM4zAp4P5NvuRTDxxL+lMtoA4BsKT4y6qJuND8AS3mi0h1xATKYSFUd0TvNm
x7KHJAUK9sSm998+BQI9OkZuQm0o3x0ptANFsVgfqOajtDzGFYHKUd2zCFFxeHaykWSS7/UvkkQ/
K+V6q4T5ed1Ou0WzxpPPW2HBOOB4zNR36Tr86H/y+cjQI3ZoRT4R8aZsVctTpN2Xg0ts47KJsKdY
VBSUMmE3sAe35f1WAeuDDVKcrExUQBECrbGalQuBwNe9SesekTc1yrY9qOXMHHCowOK9L1sOkaNB
wXnqQg0zJBVnIcMkW1NZ1GzgqECrXQlQ3WAIbtqRcfG7GuMMKKueNd/9znBG2VQOh/9OWalA8aUX
4/W7RT4nMLz41YGBt0jbGvIo4N4zrHswFw5syHF/tn+gmvzp4rI4XOz8XF+/n9LKRRWq6uzUotMR
Af4j58490pfPPVVJrfx5C1Ed3RItlFeLasDIsLieSqyjkZU2hBvdHesFQK/8c34ayuq74kkGxYH1
qb95t2l3QYjtJwAmBV0EOdgNphXxza4Fk9YnFiU4YqWWLxj83hL2VlZ6SSRmv1WUfP8lCo9UbV+5
DUY3pCxPqyqZs9vyYbvGSeD/q8Nc8KnlafReOwBAb2ZfMiTWW2EyVRD+40MyIkcpDK73gAH416ay
JYcajxJXrc5i3gvr9cFXSoZm/D5dLHs/mSglvf/Wy8YqLJvA/i3UcwIUbArZ/ba2CIolBreKOB0P
bDqv4vMEbKmsuS0DLlYlMNSgqT7ZQ9Yy+NpF1hsFdSgmr6Z0efVweC5PPsmEi0mQtuIP/B7rYS+j
o9028gBjZ3MWLZ6Qd7DYPwvkKOwJc4/2oDUH6/XOtQ/Qs13q3s07Wy4dJW6hsa5OXAHOPSYpEANI
AS2U77qKVz853CI2MRV9BR8HhY0vpm1p+TVR1ILF3ToAexL2o/PWZSA/DjGGNOrbawrN7GEC+Cg2
Pm6NDhMWM3VNRKpzqUmPcrHSxrlpyjbvUSU79dWXsWeatbIKn88qQD2FRKi+azioveT304Y7pEDA
Ou6+VVef4+3QeXk+PactvcwyPMIs6YurLvPE6T61hCyfDEpio6B8ToDGG0R6LmNCK1id6eytZeEj
JmiNOaU6KKuzb/XIrBEAmyTT2pjJ1G90/gtlmSD7IrHB2DWo5Yz45lSVIlyI3dvFlHkKIRCnmPyA
CGrhK806o4HMQ4YnHTj2rEzfFHyna/iX5VdX988xHRGNHjFHm/cEKVYxJlZOZGBsgsqKfPt8nftA
qmskClOvVQ87yoItEevs26Op0hwaCB23Qm6cI/4uQxyq7dUpDElt7lo7KD9wzsu71sJ2xmKr/Q1K
ONixTWwWpTpKY8uIs1MwAt6MDzOhcY+6MKsOJrH1QnWNT4iO+LjFkGGPI+rav9/Bj9Uwz3+EbOhE
OLJ3+IYaUH5Ff9aGYInKsgV6iuUhWhfOh1Z8ciy7m9SxP2zkH3UgXigDL0aj4Wdyeh9eZgvl0XM9
GkqkQnQ5jrtSWBPX7V6LvNose/Bq66SoIkevOkEYYB4/uOGACibTl7Bxfd8C5V6wgjSMokB5rJV9
w0ask6i+zZuaUIN1e0QFZsPRjQdG/T4Jj6gp68MUyXTcicYJhJ8P5AgTfu65HZSiwIsXvsYzZwzT
5PdgQAafiluk8jzZ25UdCwOKcgsbcrmlgfUGvD/GGSHzGTZkbnB9GfeKVmaNwlmSvzap8GR556CX
ij1Jidr1LEWSVuUMOnsumD5cNeJvabEFXDRiRVEM14qT5EYex9jOtG87a/TnP1TeBV2dgQVs6LWs
fBwrAG5PVRMg2A3FsxXC72QUQuW7yO3tD6KELkcKyisOVpPewyLGWrKwYKSgft5pkSqvzUt00Ujp
yM0NAY2EnWgt/EbBdQBTJzxAYsXlsBTh3Ss1UUqUc1x6taVnLU5Vlo5X0izn2fyJMinJ+idlucKS
VK0mtrYF2BUObf9kpfXQpxjNB6c79DOc2jezWKZf/R7ilVT/Q2omaO8uhgUbvrq4Vdw03K7BiDfp
Etw+J8qoHxcg6d8Qdd3XsENGZxuXJUfWtyPoWZk1AZ9K11PgTPuIQqhUW/m9AP9D1Ktoihz+G6pL
BM1zCm9aJfOyYWYDUBBqZwQK5qIYGrtyAuZzNa1JZhfd33Xurqvq4g3AZV8HhRmTceAjQAHSYjUU
QbZZyEW4GR/kpGDxcI2MXwNmh7Qx+w+Y8LoQcc2xHUwnQflHA+y4ldUU5Mg555bq5B5Fx4hAlaLh
zXxgUEvuTx8RE7pSPpVJ5QGEyLMhd2mfk+sDCt/7EKZCzvUhc4S05rHVGxKX+5p+pFHY32hl3rng
K2gNX7PeUacKY4IonM3cvMuXidomYywfms+QnMWQdwUlMytjDKT1+UoH+GnsSWQn41dTLE/pGH/v
BA7aEZWqToSBa9P0M2LAdcyd7x+SoU/ZxiZ5PcEfilvT/Edg8jLeb3qZs6/hZqudi73kHSH3SkmT
sAObk/3VYqq4je/VaMs98Pdw7ug8Hox3SGN6uUtGMwUE/4OHscWiUhzuM11TuSrd+QVF0OUOePSd
YomGMXvjjJeMWRQrYu65tHxKmEsStA1EOoGE9NKJnAxB1nJGelYHEHnObUsEm/5cbfvjNsYonZO8
vHK0gBEyRFzfchVswh3gT9pvAnkL0bLmlNyKgfvbXYs33+YDCf0VzW9z6z4Yjc9PsIH/v0HvY1VN
oU5/BGgIs4G8oCl9HM9x+r4ktaY8awoLE3VClem5h2YmQJSWVfjjW918mhXDic/Kjj56C7EdXSQG
3YdUEFLm3cBCjnw0SXciy10P8jPQMuKlcLRdhQ0DhnfTL0IMz2d1fEQUAKT7regyvjQnR+Ej7mi3
Tnu/QlDa1JNNJWQHhCalbA3TEZj7pUePGwo13jrhYsA/TLXdbZmZnYmNhCn1bX021TKvXGU0aaT4
KZUujAZ3aImCuuDaG8rCZnmdjKP2gDidFg0Q5DA5PdstVwJMz8Cr+W6RTa/fhtDrQ+Dir2xCVnAU
ptoPWF275r2Hi5cp58J2UqaaO20BWZp//6fxhLDKN7k/rqCEhJH/a/ftNV7G170A+a2HtvEZSTmP
6cvcxEzR0NTrijbhMP37530JcsFEQuwE7jfJV07iKVRcr3vXTr5v6hVgaqWiUIkAlnTYs/WDwftO
nFeb2jHHzLQtngwtg/IfHajtekOFF2cvdUOL3+qpH8RoMBQK2wt+xmVJQDCn+5nAjMhG0Djm/G75
zEIIYMU8zq4wgI1+l68YEz7UfRlmfkRCzFpLTombb18ts0pTEnp3tQVVRTRXq+qNPSeAyEdCdaR5
lURbril2CK0viYsQpJlWIYp0dd9XBnxwTy5nzGUdDZGxGpAoFTupbzeCyDDf0l7fHMb8/bcwtdRf
lmGFtQKvSfzNCaS/OqMjPXmvXEyMgUFRz2r/0bnd+iwY2c46ga6PCwJDsv2Oz07VmrKmCczX0Eyz
bzDL44tIjy2es/77z+aRURuiWqk/gnjFd9xaNe2E1kckxtNaiNLxnojml79wYNg4XpoMdc3+754L
TQLOUIi9AjwF8nflDIkWNl/QpAUAacbgAxYWPShANCMSjEd1AWFgnhdzsF9jA0znG3qDThaOgwVz
R/LzvPgEdmJZbrihZHUAybafX49MI045/uThjc5+pssiEaCPnMlSuU27+NUEYYif8I7NGto42dSX
GvClGgtyUvBpQoNnL95ilSEpmJixO+Riszg1TNI//WswoavmudvXvl63ymXxvV70n0n8DkXhzwuT
u0CD82ok4dPcCTtMO0f46tB5rcdLMc32uQCIGdxj9ujragJAhMh3yqzAyvIV3pmf7yg3h/nuW8d7
mmMUCmmh5Txo24qVo126HzRVOhIFH+PoQXDwq4RdRVXQXTnHXgVfmnH8UCJOEgzmI6uJigESTZJQ
AJhcLodWrGmLOXDz2QLTxw3TJVcchboqy4E8QZJ3WFFWp8Xgv2QQH1YcDVtcV1g+SFDzrFmP01Tr
38dc5mZWgHWYa7PMGcXdGsEiGvYygtWWA+xZh+nPrw9qsaKQj967uTs3ElfZTAF29k4mg5YCcw/d
JMnwaASPTQ89Vfo7s0vy0NhLptwX47e1VqHnI6yDrdgx9bWUILnWKD5jF+0FFvQrfcZeBJHT521+
D+cJiknnni1DgBazKQ0OU0fMFACjpKobhW9Oqyt1xjOZN4/zgibUZ28k2enaFvS25UInJR3ePETz
cp9fX5SxwUGXZ64QM4e6maQYh7afrPnKjRNXPaBTYbYTRDPRt4hITy5P2LqFPQ0i4hdBHy9zer/E
o56Ejl/PUzewqYRd6kceuFsjfuviHJfG6DbjMNEl+0QuFQvSP3Akjz+LMXGGwqVgQv/xviCcxISl
kY6vcv+x4jh+9wQ+iCchMFkFzj/ftKh0DtA10Cty8EBKvmrObPKd8Qxwv00N95LBiS1fVyVs/p5D
cj7CXgTtXZ10SSsLI6MbcTGFcbNXo5dN+G+EjpfQx7EP3AwrRcvlu/pO4w7K2hZ+RYeHGuyD/sfC
fBi4DeDyEDAf6eVwor6Ce2CH59kzOq7QrrijC5JuUsiZ1cjnoCQpwxAeQ4fygSl16XnnZPNGy0Yr
Rhc9U7qRln9BMe5n//njiOJFwgBlvnMdOzPCw9Y3KPmH2eBmt3da9Pze/fs8WYuXUNj2VJ5sS2+K
husILYgkhqRYrzJhwe/XAdqCpt6OeREp0zcNPb14P96PEihrEDeES05ZzlS0p6uipB0GCmton2es
InS0FuVXGyivmMz8I/la6AF0vmQfLzJJepbEGLwrBC4df7aRb8f24jYj5D66wwbuE+gB2Ja+CFhr
lRLwDaqb7Oip8h/Lee8Q77iJVZ6wgu6bNVJyoX5767lDLLc0W4ZRBAMBjlIZ8zkhTmasF/SGYbOG
tBkOaXOMEvsKmKGYEfyqeRmdn9EI26o2YVEh1rZaSOrgs882XoiMeqOqmhVZ0LjXpSwgXJavMe5Z
nUQqX3YLXpEO/GCPC7FiCU3tb8hCEiO6N1nPTWuuKfjQFyuIi3+2l9edIlqyAs0qEi+vbXr2Rnma
RP3WKMc6eQFjNft89K1N/cLjcoNw84PMbXmwjCWAWtXJOZm/3bLAYPIIqMm/EBIhAfVTn389lofA
m0LLzlWn/THYh+Bpyh/3mfEM6aNyNIiFY9KKeoD58MNX1knhlC006VlyT4L5t0LC3rKiVYoeD3WO
ov9PlThpOHxN1R1oxTX3+igPu5zTPoNJAXvAUOFT7hoWtZkgch//Sw7Sw6CIfctiOt7sdAjQHWuf
mDkBrDGRG/q4yZK4eko4hLjuJnnS2PYXRyVfR/Naw5yCTdze27FuB/zYvLK1JgKdFBjDCr5EnfTh
HV4SyX4vhI8rWgQK1lqrAMBczOPKZM48DMxlYMAUCeLLl6EkOLwb19fry2HkM/xysmDJWUXTAxOL
KQ8tI4GZVgFRt7y+3TrieyQGsPl8YQ3nFscB6ud9JibgRG/0GNHA/rBqCuX66Nc/+T/hP5XNAyBY
SlJCs+LNSxXUusmKLe0pkuv3Brh+LE150kpc17FoPbC43sztFTFoV94Kcsshh1VcrEfKKzkmt9dM
ek0ppiq7+pfjEcn1cUpJ3GrpzXjJiONmcQL94a1qWHFoPYQw865UY31O6w6YRIeqU4JcnkgPrdqm
YGJumFlwA3Qtv/eZI6jocDPLCrxjuCm48+1Dsq3g6vsoefSEcnI4uZpi6UplzGYXQPbmDxSdrxXv
RsHqV+5Z3+LSDLO8egurJl9KcE+Oxkg9MWP28Nji012ktNbIcl08g83orzFpvvnrLe4MgJDjRGci
0EsbcAgsszSCWuew5EOb/IWs0SrArutuQYKWdfZrVeELCXarK+NtZBwY0zVkj06YQqfovgPktyC4
5k9BKowDwJ1VrR3eR42gsGhyRU9DvqTaJXXx+Uzhp41Eib5G7Dq4sHMRFZxD+pLa3Ukl23BayNFX
1DxCUdBLQaNDKhRqo0wdY0XUSoB1CWdQMaMjtdN0f1JZprQAuVj3/SCq9X7mNCgUFqjGNbwwDuQj
FMG3dGcHtjBArA59M6b8wnJiJgjalPwPNx6GV3D+3Tvsa613H6cXCJuqSdGwIbsj0p0nX4OBIo44
rVoyCF/b8L1fpEn25hR69X6Qtv7LzUWizcSVbfTIzu7GnRb1gAP04sHfHit3NqKqapfhbQEWNgwO
FS5ogY33/GHHg99aeiG4BIZ/qwPIcOMGJ4s0sc1+e1JFiNaLY5C78Arpg3nxz4wwTewDxtmzSou8
64efDa4G1uBqZz4T8LM4AVcu/Zvy8KHDeSoUBf7X+EPNYCuYJwxRA0CR2wcRUu9TIaIg0ZxvNarq
rXFHFx2NR5QcbwvQj0NtgIC5HeKhmOAvYYDD5inbWgL/eX+KXyYrLeRdohrBram/GdOVXZiAIU6x
mSRSqkr+FauLLTT3LFB1R6ykDgSfnWu6AeCL+djQBHAPVZZ9PqyA9qUxHf9L6B1zBOV8UDE28MYR
mvRnW7czCOSSLRLB+H2ixFmXUoAocfimCXDnm2Br8NDtuQLBQxZ+1PWCh48/vhNkCp5VTjNV6cFd
q7fu+q8P3A0+4a+t55FanAk77G0iuOgn5ITlYW6ECFMGeaJzr47J589ZUWgPUjZViHj/kCnRG0yV
5mYcv6TuYu1bl3nN4PRm1GShs2KfUfZ5szeqD5vlf3qh4BpQrtNCaqMCdORO8Ti1EVKZbRYP5oXy
r8XpH8kRLdUS/GGLh95Kmu3OMXxgYRImCddWq/USM9mDbN2zYS0NsK3vkVcQHV2QBEnFtoyU9saM
IuYUadIGZU+d9jGqbNCipi5DzZ3fl9JQagpzdG6XxBVH0czTiPDN5xKwgQehkf/bHUjpiyrqPNuy
EEMGKYCFx0XkLUDWPx29jWzogwNr0d4XcXri/4v406sg5s/V6Q/ZjMCGPfGxZGYjxRGy0ZKmdhYp
/nsrdmJHwIYvkbd8ikosEfB4MET0MwXFCj6EoURVl2bOYlDBez2apsbgPkVoQCWCRGe1YU+DSocB
GDQqVGIFMAI6FZbODf0XRb+0McsFFen5zNNHtAugRCLhscmaM7P+4TKGD/TPKDEVBVQDCxpRfG/u
ahl6BCd/0c2I55Ao9ykji7bTv6gp8SwikFz6hEHhkmyVxRdXS+BYhO9pIUNktVtsfKasIA3nsVM6
+6z6Ka6OjLebqnut3kKEhg9BI9oZLaD1uvaLXxhKtcda3uqsjPy8QNo4Y7OU5BywPEyv+AlGQ040
FjHO+MZ58O4SIolQuah14VbkJqEn+4YzgeYVAtMEnLa/aSEOdAWuLOtwBPHB99B5Ff1gC8o1kdAy
tQ4AS9qlDGo0whxHMwUUGUmWEBbYZFuSPgWRTgHhIYNSOtfDQvq1Yq2IoDuNjouKto1kC1BsI4V6
dhIisxrGKqz1mZBz6o5JPGB1qUX5SftK8Yg+cdUVy1NhKLLOicTZSaM17uZ6nvLK+S1HGl8p8nv7
vKWSE4wkjI0ZYgzWjh5qz/MkXehKd/YeiffjFImJUT9itsP2zhlYOz6j0XpaeLp45NixBtv8/FnP
XXSTOiMB+fVQt128uRcQKhxYtk9Ldi/ssg+ZCGq0mkH7Gp+yVqeV8WuppHhs8KmIB4DWJPMPnSYc
4rei+O7oK6eSODwr0RA4Ow8k0bWLEJ4jBekCv51cAWDW0eIzXhsnVV1CGW/O7XZZhbY/5Zz/Zsqv
fcpeitSvIcNq7q/XBa2T1xuwpEUIObPkIoMm+c78OqWVIXtMHF3UoQbeud0A6t41lE9t2tApuRNr
aI4H3NFGMzPbFsUfIfGPlGbqidNX1MZp4VNDpvov3gGsX1QZKIXW5aYoXUy9RYL68vj9cHRjHYLa
Q9MvdZ0B7A+muLyTsZJFImJiivL0pznjngUOrE2jx7j7cybW7Qz+DuxCoHCZ/Pi8ymTSVpEhOdRI
R+PrlG78Ax47TnffjUYZLugtWpH27cVie3qXX0rvJgBRva3JIthu2atDxATdYiMU8WsKlqV2pCX9
CoXtfJDaPJNMfdkOflkLWYLWCNARYquqxuRZmTrX/AFZFItdgxZBeMWDjk1/b4/M+wF+c7MTmrmJ
5er9BiT6DPQ3OkbX5pWYGydbh583MjeTaf9RsBPIR9QqO7lbdOAxOHOZIejIiMODwFarpwLsG+Ls
KDULalYIoAPg5JjbrPLiL4ESrl5ApI3XXnR0J7SxCCJo4KQpJ/iLCCunqns4x98tNpWq8c33Zdr6
/nnQBowneGRCUz+2uTvY/LUQ3odDpBYJNTIdEkbZ5MOflvlfElDjGgq3EfVTU5dCCJTcND884ls2
OZlImYmasqPKjxTY+7GW4SRcnk6esRyrMuGv36qLoA/agLhCk7bQXaDthbBvXgLQaW/etnWKjJS2
Nr0GPrqC6ywJ656s9kpbM6zz3YMIdVBZMgJObjbLt3hvagES8yW10IBFce7BoNkqjtPERH+ByTsP
WBB9LkT2fg1VJwNXaAlRV1c7If3mu4KpGgHz36iG8x4eBWGqTdcjjgWskK8n84RjE5S//an19w31
ZiTJBDRsN3CbnTtbbr3Gs03juJWSfTbE/pZVLRmAwCuZVU2YVB+NiIjFYZ4oIQW1qfpO1nDxsoM8
aLx2FCWqwbA0MAg6y/dXavOioe678+i1h9Cx/WC9FVmRi2hDSqMPcvnSKP0ejfbJsCkGBljwAus/
XARJswQUm/wKyCZiJzzD7f6i6aSW3A9yX2rfIDjUmELdvXSJpubCp1ez1bqK8QEs3acnLB8w/V0g
urj36A9mlT7M3r/A5Mje/z3D5yR1GQTJokXe0ZUYlaSogGcapME6VBqdn6budiFQMJ6r0AWRSSRH
odYoRz72cSfLsMQSazMpAUZA6Czon5U8yHWw27qLHNvuViYZEXDfFV/PVyONbokD4q+sqwqcyzJd
Fj+lCKVxPVys6nwdBLh3HGLm+sS2e6ZHY5ecObtZFjTa7rmmWm2CFiFIHDRbS7E1sZ21NJ94VRLk
TQh1v6nzQMjBtENiRQEiufmuuAv9fbpWNDsbSPxr89PzIW5qsDQ9XfqZBAJ6i1jsHYhMkRtytu1S
xoD4J/FkpJqtTgNRv+z9pvYcwWitM4kglSTaGuV2b+k6ydtzeQKecC/0M1IyWZPoeePJbu7pQITT
8Lcdgk8+AC4fJ/hT99FYdn+mvf1b9wYZZ96hCAFb8wzWQfP0Qkf4XAdtBcwRB9+IcJw6aURV9GRw
S+NSr+W9bcN/BNdLDk2aMWEPerGNRtZJFEfDvp3onNTY+SWqgwwGhUAJQmteTLDhIexiynETEcUm
i9MDqDNnb2u21fZmuRZaNossB1daRkexJF1IhU/PEr0e0zgmeUyWSzSDon0A9ulVfQuI2R8RGu8I
j826i/RmWLmIarvoG5UL8KUXq6s12BWfh/i6yxVuyjeVBDU57tIGbmGXmhKcsjg9crZmx7WpQzY8
ebq4yEWtr7FI4wZ0cV6B6CwFL5OUVH+CsksE2LGBrr6pronh7rgSvAj5mideVaty+f4HIFfh2D/B
KLqExEB0rAH2oXdLIdL/k0c1oeFSjcO3BW/HxRDq/dOkEe+XsM2tzwfmckXgPztmVOzJShIIqv10
jDHlwmPQNEHVYlxF9hCZUl98+kbAQMfB66khcAL8kbS6nz+aIvGYKE7PtENy0eMXurAt/719fd7H
leP28ENgXZcHgFJJ8fsWDM8iGFgogLz9uZybyaicxZPIEpXkw9YDqg7pLBfjwLEKuDqVp2t3/kCz
R1R0d4dOwI02ukW03Cge1b58vzteu6vuOElJZbaK63prMrs460qeVFGXOHSgTR9mtUeFCtPkk1lt
AU8BdVxIyzwEtM0DWKB7BGD1z5WSCGNx1n5V0SlKdtVOOjf3LlKsd7pp5tyQRE/EtDxlx+VGHv12
U1U47fpjqUzXZk+Ouv24N1raa0CUgO98J0QSFRjjbacK8rcPC3tYUI3XlIHypKrJB+3XSvtp3+c6
I5AJPW/Jq1csIKvpMJbvhiKauupVX55nqyN2kFl+sWNV9K68gXYJcLhDFkrFdOAHjOm9CH3fIo91
Xxn7UVMgVQ8saM8XBlM9+rfuTIfBD7GoXrop5LxhNawAl2OYFt24ZMUfaiCx+Aem4EB9otO69Asg
Co4QVZe9RuKiFrB9pVvm0auhps5FfYsCljgsCoc5APo8OJ+w/QSjCeqUsFKoq2hx7GaJ3SkdqMYC
soSPLud4efN/5+DJIuqO1CHJsAobYErM2uW6lKIsr8Tq3dwvgA9kAkF3Wun37Uvvxc/dOEwlBmbV
WGxgIEygi4P65wnc2VepUVQ8sVKoBBO1zEafej2fO2a+IFUTYH78pd6uC+RgFrzsocyokMpQgUfb
+WYAtAT8JNVuI72VYVyQHBqTI2R42Gl0lRN4o1ioZzpA/iiPKwOoqB48EIhMLT69RH45r5KypDMj
VawePgcRJ1aW3rTueBOJU3a0RBHIvQb+VBtgV/YP0xfjhx+lqT1e1sAccEFQmyfsAbdfW5BNRTdd
MWo668mGwV6ltazk9ZkIaTwauQPgJ7waEBFHQQaXyGSFd1mE1WevzB/0rpBIwVAbPxQ3SiJrdyA3
KZkbrsQljluIXT0A0iEdH4N82Z3nkLnSUqPgasbohUbnQHiSUfCR3ABITfxxD+LpmROOwEs5TUVG
vWhir7Mu8NWIiclaAg2ZB6rnFGNYfXPsdW0/2UPWVWzDkwQlpZvJHllMIhh11+nLpnQCzkk9rw9J
fkoYcFrYUBi3W2jzb6DxwOsqWqXQpZzL+nJeeVscXPbEY7/XCMA2v9qPEdjdSOcid4FY1dPzlwuD
G891fU7f4hYgdZZLR+HTmgpMKhIIihibBcJiXYXgzpmBHG9DFAWUCeEWdSJcrOkC/gpFkwjLUoAV
erEr/bvC1I5balDr27ZU4sCv2rz9lkZohaqCLdA+qk1WA21ojFnOI0yUUYNLRgkiVFaf0ADhRv+N
lbi7doCQLzbV63/29HDOMLP5Hcr8iFpuJX8D0XRdkQiRiVpuD9iF/6dYeX0AN3X64gCmInJv/GpN
OfYwcJxf+Up6S/bKm8V9FqIeiuS+6MoaBAyLxACJmNTkpoi4VJADA5sNDTJjo89ldpUs97NjoQ6M
ji+NUaj2z2rH7ap1EuKnMereUwf+8Hy5jKkDVWaLV5m+YDE2xhnYmW1iBcwmQoigFmA6EyTuxZ9P
87LrkLnaIu+Y3A1y0BJ3GpfxXMI/67c3W6W+mkCes9kFkQ/+Y+WJDX91s1tW+skl8JJXnhr2V53n
RIVH6n0zqx+JPY/16uLJr98h+y94kyP6dP119KL8f/VuRYy3kRAwiSCyVrv3fnr7MjvGGu0o1NpU
0kF3ono3MjjwImTeWPaVLYnwf1RJhq5+GsrfpWFVO/Fhprp49GUhlEDn+LDkKAeLWhy9JcwQAOIm
cFl9j3RKY2bxtNFyy9vxK51YDPIJFvQ6pglG7eCl9J0H5IcI+OsARUcTPzPDNMFWDj4jKl2ns5Ny
u7HVhZQ4mCmCHsoQQNouwthJmxHqFVirPWCzJLoUgrLVWi3AvXPx4ESaWKdy4PdFUuGR+fQBaeeO
hBG5T6oKk2pZ3n42Gamr1RKrpPWRBlhQfqvMN9Ih4QyASnhAqVW2B+Skg4eZTXimXLPyW1jNJaaH
mF/rUX1X8CWIjziKQX/UpxBNB6x2YNYWxMCYvjT2Po0AO1FHpldBmZLnTtt0cDh+eHG6VzkVjPqg
WRgh2Zs7UQ2Jl8VV9+EniBwuBu9emQOdvOWbYygBLvv98KYL8UHaedb7RoQXf+ngGpOLXmdOrNqL
MU3PvMqisfkMe9CbWH+gWPsN+fQlFBE61dC7V/MmWfLiHNrgiaoPR9Dj0oiBWYGe6cdzhds4lslo
jjV1QKNKLowdQjSZgwSPXqqbUpqiyMQc7VPdx3KTBrkLd4d2gpe23huXL4DBqxuR4iUlPuV1uLps
+PI++6EG2n9M6EqmxmIk495/1X4ucoumcSwbuWdYprzLikRlRS4E9BA3Gbj5VOPmvUhCUSyT9hDn
DNC+XC55p/6fv/WF4UpETjkMZhFLlyqRYpLIqZAMBr/OYCS+Tch+g9ntyFXdlxdbnfWAxE6NLnjK
xO/nz6FIsb5vdXD3PHjdVvdCeLrwn+Pz6f2JqtXZJC6KujAXBrI2sE5gUfCxxQYSO8DdeZUWp0OC
rZs5snYTM+Pv/tCHJNV21axhSAOjPcU1iwhbSFj35KOG4w1htu8HWs9pMMsVOgbqfmSJfGZDVkT9
wwQybi4+ZlHp3PpPPvgE+fiDBmmxtkM8hdADKOPchG9ennYqP70WYobFMApcRjC3rMns5qxoikqH
7tNP0swIoMvcr3U1OlgNe3LQ6GCV8/Leg4iXn8/u07YZ3szDUtotEPDc4EPCIbPvqmnhPtMBHyXd
b/3qg6SO5URWeGWlEGweQ1G5c2nhrnVFls1j1f4BqLT1EZ6bBU0e6rNNjmXbw0l00bh34LiZyUyI
YTJTLu3rYoDiyCILCormklMwB/BwFvt2h2lNrLI0XrWISNLamF/E189aolIQF8oG0F0yP6UYHmIl
GA9fO6DM4TAv2Cp4eNyBq9P5RLDH1uc7NYawtZToq1bKWj2iESaph1dxVfPgWVecFfmeeD5+7Gn6
VGwsCQn8c2HceeBOa1Ya1/M+GBrazhAITdS2VBdhhCVPM92YEDEseKPdTLAz3zfAi5ZVKwsVZ/uy
kr12VU1HALBTXdogy1jlBQJHal2P3vlrn2DDI3xcoorNvpcWWGlf7QtIJnz9S4gfi2y7qcuqBDi8
Id2UtT7ZbraU+JsxuUpDRzR6iXWQQ+s8HoV3jjUvFfYmt3DFhto6OlzaJZO8lhlzttaaFt0Qtf+e
AyO/fQ5J1GC13/weoCwm66hQYNeE3M1n+2D2R7DQcdHNrTZNUEvo/Q3UWfxhFBslLJDTRr74kyWn
k25fkwPUn2LDPEvIVE7N58LQzm8Xs/mgG1xvYxmrxkdKxlw0Lbt4tYE4bUAmvyDS4CL65SGs7exx
YIuR+R3vXnm081X/ciXxc8QhEfRuZ7kvsdKX+v2Aq6zRiWFUzQ17M/RSwgx2GJT07dCgR0sUnpPF
ljjmMCo7pf/FheBBdXOkryoSIgTxtbTFr0xMr5sZUaMAnslpSq5llYY3hjUMmx2GjjMceuhqiKRF
CE15Ga08V6XxRG9bdtqfVe3n8KKm8rs3wwa09BxMK5UQfnRvC0ffOmSJgyUt37BtxSqvysWWUd8w
kV4PXDxks5dH+ZCJUGpc+szHF0de+2gPeYpZnFW6g3mR7o1Ku+QEopiT5qJHzLXgJ7QezemyiRDL
iPDSVV8iJlBOMghoWSEKZrARUJmaJI1t56DlK51ZS4Y3QIe84AeWu4297PfaXbt52IpYKhy9Zcag
wHt/cyANg8fq8LlTJsSp0Zkvgg1UelVvSagg1mGMIxldSe8S/M0E9L8SmZkOZ786Uq9Gl8WYwkxN
bRSw3QLoW/lzHygApG8lcv4K0ZvDdySXRShI6RJX01eGZhkDDG4tPJwniFUaI7Nnq0Xxl7UUXq3l
b+rM6Ck3nUkn8nLK83+Hnke56LWM4hLb7hI+cGA41mUsYnswrd2owoJnLogKkNUXimrFtOMtGZ3V
8zTTskCjJ2ABzCSGIoS7bjOWy4l+v7O/lV2JAVrFE3jc88kqJC5SFOiUwrg938wx3XKVrlIs6Pvr
AgDfxm8DR/v3mPvGRd8lJ/O8Hodn9oDmJXEdQhbl1NHyHMmMDq0w0bG4Uj9htZxBxFwC54sCtUam
p/XtYDJjytmfEQR50FBjfZYeKa1FSv1QifY9LfQmcIAQk2ekZEuzOsKlpOor78KF9phy0vsKE8Mq
btY/yCOLTH0Aqv4ByA20IeMuanIGET3fy4paYTvwuFsyHvMH2jwSYGbZvZ3Pnnf3rlSQnBf67Sw7
nldWjHVfSxS7dKrDIzloC1ucDhCPJrm1aEex4R8uMZ2JSj/3llFx1TLCInWioTSB8pTiErmLO48P
qWa9qnj8IlyAIKoS0zvGw2e8qhAWfbGuMvFeaNfo+7GuWLyhJU+FTnRX3/ihlQIx+b8wsu4BJFaY
vLwDt77KApX1Tk1pWoj/+ijJROOTyK4ZM1BiKw0Xooq6b9dwumq70lQac180rQOhsHDiKyjtM6bh
dWHh+pt4T9Q+cbNSbiBeNHcuaM+Uy3P6WB7UI1nQrkD9BpMbg1PfvaGGa4CYWHVQXg1ZcBuFseqY
FH+cbbxaPxJlMU0hS0X5cr/ZTJK4/h12bgIqUuNNv5iPczIMmAwU8SqiYpGHnNTf0mYVbJrTFJn2
wpl2f/1q3k834xIgOlcMg8J/0bZMHimgQPfHGiQm/3Y6btjNJSqRM87u5Y7/5w8HgvWo9pF65oXp
lIM7XO2DO5IitGv1N80YcTI37jaCxOOZXTp89X7eZ/5fbrvAtmUAzSrxVfruLEjxnArA7mph5zLO
aFe20Ym3d8EAfGO9w0QXvTvEM75ZCAQCRpGMKyJ/LDUY6ute7c0SAXgC3cYafMFmY9r26zq7Yttv
mPBrksvGrY5DMvRJXDKAugYhb7SAt6zqvDQusn2ar8Q3hcx+Oq57Bwezf4La8HBUStFD1I+LJJ2j
InafdW976JI5Sx8gCz651z20bO6PwMxqDAr6hJmOEVIbb/srVpaV3riapsBmdhs91Pi9I2BgvHHD
Pr4FOXAwJq8hshKteYhON5oiAt5dk3hFSl970e5m+ekt5uswDEQk0kwk6xdaIUGdTM5WnGBGAUVF
EOLGlhfnZgxZWRhA+rFFdrOJbXm6k14fxJ1Lye4PnfvrmSNXiXd0ZYoZowBSLdtsGt/R82icbMLs
0uaHtHA6xHY3TSmnFgOLbn4OhiYpynggbuJYVfNF1E+PI/qzQw0PJsDHAqkpULoOb5e7LcM4Trae
gk2tVWcj9gGREDBrOEIKQxzBkUEGp/dOQpr2eKveReF1SbFoH0KTIngCoa6P2gy+IaUMERZc7RnV
/BckeL2PhtgBs1cw9dIuif/1UuQ3uY7XPebA0N1R9B+meD3Gp4gHlLQcavPd/FnbJCOputT4uQ0N
iLlI2bX12Jwrp0jRKM+hplmI7XOmKCzu+0cdQ903PYouD6qOI0ZKRfFIW5gZ2TYcJT9l+vlpGkR4
QNzzNEWopymzo4jBdTNWrzJkZqC+oh8d0KD+F/qtqnOO3fNV7QOWYRi3fkIpv9a70SQxKztI0RPP
tMjm/o8CWhg1aC3VF2yKq8CgNFITpwOQbgI4HsRtk/wSLXLAy+LL7aXkMM4a00i8Ep58yKQ22FPW
kLH8udQgZXbGlsWvikD8XmpE1FpE/HM9uDBK1Ry/xAbtUq8l0FM8nLOIHZNYl3fv7PuRagBrmk9n
t5yKKoV7gvvUiQ5AaesjOl1wQLSiWtzpdxUin486En2vXQLmwtsN8bBSGwwe0fgboMGkuU63PD5R
PDIqvgRQRSIB56+LIkLIycf14idtBQWAg1OihaxRMXaTLVAmIZcu4oiMqHg0B0d/aIfnhZsUqB/j
tekn/yJ0QN8WYh7c1V0SI52QEe/NmSbueB6D1dyBjF88BwbYpGcWzbu9rWFgzeAJJGGh8dZti9mD
pse9taaeeMJ9AvhkjeN7PL1sMWYI6VRIBWqFEvr5KqjVkHCJqXHyPdsp38HWG91WtHWa921C7gx/
xE0SIdiBMMqc4E6a8O9CdrIn34GyMWndEPFOotEUBuIHakfVGngfKi056wOX9vrNl3hfIenEJZUF
bHgoPxbI1cipO0VGObBQXGN48+b+Ii5WwPwn4JJHw0mqdjRbw/VKY6lcd42DLVo6c4kpL9kFPABI
ooFo0L/prldqoSyFLQ49vzysDm+bcJBA7TnMCTykXCc3ijMmA3/wOjku7+xtpDTTMkUDrgE+Mmd6
Z05NLjaq9IadIV+4G27dA+xP6GzU3bGDYM4wzD1e9h58aJRk8Z24Wc7akDSEteqtvS0Thzp6asKV
3JkhY7cbk/vGF0VU4JjPOb3xGrm8pbelNCJIbVGmW2socxQj03JTqXLUa5bcg7N+JoJ7xYZQY2cR
HDHIh5xuOrzkgaviWwJ3PzOQDLi5prwPCAeLX9m0lJjdqI2hKS0BGnbTCS4FG7qC8tYWMfcRWbUD
pVyHU2xBrf9eM1rT4s3wVte6++7qJtHFuPVr+ERIhCcaeGAfj+NNrexs2CFXlCNAEXh9QHy6pfrB
T/ujmcW3II4BOWPbKDesBlW6ECBn9vcV5GSnniOrhdfGuHnDWoFKyuwiMjeOO0Zhl0GRL0c74jd6
W7c7iDnHHfoAff9Ce78lYpGYeeRTkPtk+aAboSn+hy7oXZyNJMgP/XEWuxeXRY4bqpBoJKigO1CF
HoM4OtWdiHHOvaAWIlzyHfZC3j5vCe6n8g5GA9W37NyrP9aFAecRmrE1aYnxhdD8+g0UA/WvhftK
zgKMAcqXTCcjSOjz/sqZBIOgqwNlgxEWVRvqj4ZdPtCNa0o/aKd2/5Kglp6a8a4wrh7DJlea2mek
pxE9hG5KFQoC39pVcdPgO8rZp+fpxbkkbQNb/h3WBGAsz9ud/lYFVKwv2K0naFuaCNfGpIKJJcjW
+zyhKBcLD69thn3IcBKnrVT/ts/jCqSFCcHsRFed1FvdRI5nLJEN/0diCijFmhHsRDck/8arV0kq
unh84w7JfQIdlAOgx90vN9SZUHRiw72vSXoTznqjy0le2B2GPkH+bItQbfJUMLPoIl47f1oog+yr
sS4VNi7baa66V/CQEeLEyLDKDm+Avh24vJ6vNELP6vW5TUXwGEV4nj22LTRZQYOiPyB1ZypB8D8B
cnXHs1k5vTr5KBw2JSRYaSnWejuSw+mActn9rSLsOfOrAz2NJZojWqrQI3cvThEHJrWur8PjR1Rz
N/R4nT1NveISZ0chIojaEzu46GNcCB8mS9swjloia+TSmnu2qYPDg2Fk+OXWGdFD2mhBYnCkoRPX
2c3hV/OAaMzDuguMnbii/JcFIcxmOBrerKSkcTWGHMmodr2PkVjdCu55QNBRJNX8NQ+oiUb8CwW6
/pAvkVi2pszYWaJYC31IAq1ro4Y2VORpEmZpT61QpeCv9p0ELMxScJg37edmvKHlZ63siIt73Tf3
VQpdSAARj5X7GX3M+0xe2/iednt5/gfKPjK3a8b6+QLDyZdMNSIpjgBuBRZhDetXMp7NOhemmNsc
Z2m4fAw+gn4EsTZgupKPtoZt0JzUfHqQN+FFIj9C/g2m7aYo5olBtnNTrZhpbp7GlJRQ5LW6EXuH
8vIWYQDsgboMKVBuqg/lcX72pY0xHA3I4P9KER9Qhr3zIaYQbwFQkVIVLIixiVTylflLyeLEGs9/
QVN90ceuQ2y9uL8gdZ3ACVa8uVPvXy3odYfu6DrOHfsVpLwBdWSZ1OYKs/ZtSnAeWnzmmWsxzKlh
bOn8eG8ftsfeV+gd/kKkCHhfN5I+zwRn/fEt7Md9tqwc4U2TBAWb6N0pfoYHP33Dm4l5uvDPH4ua
hBGrZbPZYEMuRa5DUF6dt0krNkuN8ZD123qL3Wi4a27Nqi8dBSDJLXHsq5S+n1Eo0Gg+vt/RmNuP
dI9imb6Nzsy97N4W0AWOrg1tkoY7k6jmb9k6qGG3f8VzT/Wns5sE4Cs6M6/v56IGzx8gbsWnBZQE
DVVYL5Y8mb64oDWd0v5e/spf4V8PsRAysuBPeWtQUqNLo/vyN0wJ9O3GVpeEVZffRyJBal4nyKpX
qjCdMfQCYB37U510b6MQvBt/6KpAZQcNjglIKRNX/OyrnoJYIKo0+UL3Hje6odvTUq4fvqAS3XLr
Esyjjd8cebTgFM7eCUkdgsHVVSNN7OdXHPNfJfNNbjAeebgjvZEY76JvRJTRfW5CKeIixEAMghQO
xnc9zmccGOuKdk3KNEjFlZC17WFibONQKCSs7toND0/XISWvk4MFL1K5QTWVxH2gJNwfsLWCCrNC
2c3NPkSp/8H5eLdAd2J/PR6i1rVDTd87meBk0GEtR88O6YeUrUohFD2Ko5N/yR40q9Iz0+YaX0d7
FMOC/ZJPOrFpYbqDjMDCUM9dUNvLCXSsS+e1QrfXErhFK+RpPjQ6flnA2MSCKKCmpQfjLg9gQjGz
lu1UssBDG28tlBMz8j20SeK3pnQ/jF/IeDDcCymCaQh41myIK9vvX+8QFnbHZnWyUmRWMrFJxUZS
RllV1g0BelGt20l+eUllH8oT9PKhtgU+LIWmn6IWIHDnVACWu8xmzFDSARac1wU6wICBxrSxoo48
7Oj2ll7tyKjJ3swJPLPtOs7K+s03vygvxm3D8hdxhGFKSxcSGNGyPJk98zHyVDhGkJBHmGOxuVQM
BepdQufw+ZafKqzcDrsCqD28QD0C04ryA5uvs1nl027gtfg1L+7NVjZa1n4KHdO04/YAQ6+Azsat
xfCMl/4ejwk/riaazcFeIgVokkN0W5OC+4AYtSt4gRW0czblOv5TA01Kv2kxP2GeV+UFsP3JOjDi
7na/s/4PZA4WePlNcIsbEG21UQPCeTHyO3AlbV+UIA9b2lv7KSs+LmQb79Zs0E/hw0911BDASAYg
Wl8uvSs21Q41d/BVGPgdPR1X238ksLHVxd1tcd9LQUgsWwaNKpVFw7MlHgcrNoI7tw/FtzsG9O5t
okw07T1El+H+2CMjXTR1A62z1WFLLuQomHWhy12B5ex9yl1vGHGqbpMmSzr/4eom2+YVpV4p1odI
l7WGp95ErQPECTrROZ6VVOg4rFtVGISk+xPIWCu2XZODXwWa4D2gL5G/v3tbM21KJ/kvQ36ATeqS
cgdg633Hq9WvK3WGxwB05REeUDmWQzTDWD4RtYgJevvxJS6lmdY6XsUHYCkpmG9Fo8GhOYG9cdLG
DvuJ/wdXMs2XNgIysc+w5Toh0/8Ho2iZ6bPIsm0TnkaW3yMgJOcfUma90ECduRGYvm3oM9db9Uyz
YQ9IBxRjMgnN3gH6sjOy4wPUTkDfZqlLHYMguiD5M+ggyAKD5aAUpVIu1kIk0WxQui9UA+PWs8ci
tRgAYsYunl5CQr1RVEFLZFuGpB3fz1pclyxtwq9ByB/Q1xsTFRiJPnJu3GOjl5op2d4+kdtg0cel
iPc7T6mHidng03KoNI17pb/WsY5o8hglxTVdEwZfV4WnZHSQUKQqKoraAIQSshu7etAqUAK0UIKl
/QhbFLS71Xl+OYepb51R87HmYXgV3NwBj/2PjwpQaXnfY3xV1ELT17XYFxUFPzMeISJMxmgvy32r
s4n1M9giTLKRISML/MIPT1jkIqSDA73tiVls8waum2vGhJyEfBUwfVpOkCDShClcE0vuiLHGRwVW
G53PCeumq3L++/FyjRJlY6D0pwNInERUlCMwkRBbLnzg6DOfLP5CJJgXRNv950pl9pnd/N/WENwE
vdDoMthYIM7Cp6n8+V5L66W3nKRy84i7fs3LhnT+HQzZnIIa/LyCS26hN8eyu5R3dxkG8DLRX5Ua
kiO3zVcCAyPpAC2r1t35eoA3qXOyaFO+qlmCZHJexB62R82H+TieAvrvSAKvSPWFyjItfaZc2bBm
zo3qyy3bqnfB4xdUMMHoqZ00hjhCWqKJOtvlQseuO4sW1nhtTTo0jo1UjPrWAtn3TVuznBomhtgg
ZDEKs+ggF7WXw2uhRjZqXmdsRagBmCrf8NIOQ7mZeNU9B20Yd52NUxtn/qCtMR7wl2M5QBR1sxN6
8gc75a9eh2HSqZGoT1EXq58DET6Aeas9f0nqAd1KTR8ygEkMJT/X2zUqkbkDv8r9BvLg/P/5m6Yl
m9e3dZq0GvQ9LW7R76x/XMglQVVWZq3E5W7aDd83LvxTEU0smDIWzlHcLSXRWqAcjvwpUd1giEs6
gJmEo6j6wUc3+L16LPZxHq40EqNrHhYs/dIezx6RwtH75n7OwhXJCKSxrX8Cvv1q3oRQV2oYFnTs
sUk43pgrSx+AbgoLOgVQBuAxsuQF17kb7oklov+H6/0rdaUe0l5UmpFpkvL3FvU5SP+wWWUiNujw
aljGmLchlAULwwAeyaRgSu4L5KtLaW38QSMfACxvFd/aijwq7ctJrdPWyoomIlOxqUkcmJeASCzK
dRwUqinJ3g3j+d2+oPV5DoQZvWIVihlg0Gt8p+NFBlokDzfrqpDdbyh3e2gZc7eKEC0zC5+EBGG/
b7Tjo158Dchd6gRkw7KeK+B8RxS3dvI7pPET8qhKx/MjmC9to3Pi+5IcY55/6Cvn0WTxUCcjd2qG
XcdR19Dw9/F6iXWHpSs223LmveeziWJ6S82AdOhdGDUURtfOle+5dGd4UsATDoHD3OiSchfSdA7J
PBkaiO+MTQL6kN84T7V74ohMlTyLyeapk1chCn1oy9ZYFSnIFHCXD7F/hOH4/jKOGkhAK2OYQwtk
aRPI6VA1wBFVSUAY3SeVBhxqYeYmyVPOpAE/kD5T5iprTl0kLR7nFdUKhbhwH0S2kOrHPaM6K64k
NOpg0vDeSr4qDv2HbsASltMB7GWB0aNGjND4R8ggt0k2oWvlZO9fxO43MM0W4WtyBQmveTXJA+Pl
JHdSUk2ccVwZhNZ1LmHvuTQxh4R2SpCA0O/sSV24rXH42zaqTmyErXkSLzJc/sF1tkYBmFML1BTo
LwjhnlqgM6CO6SX2vCsRm1/4kCiiGC/RfuZizFplieQSmg86ccxPms7fAPyQ63UGLdeFQFKM5VvN
4quEWM+01Sy8BRZJ8GzFDkcJttvwjzRU5xj7ZDqPwXwJYC5RX5YXpT3uedU1W+fskU/1PyBTprq6
/4N1eTTBRyp/DV2bfXxavuVY15JFaDpxYokROHhIgxI6//dSp9F9ERjaUyL26nYOnsD5SGTY23yV
gUigoA2HJEu/GKlhTnEXeV2iEve/t6i8A4Lub/yphLlIyQcWQ/D/UNtGaC2f7Xl38q0Q2u6CluQY
ufQSoVI6wtAQvf08GNoNRf49H1lqAeVqXO4X3j8FmQdJW5MMhPT0g7mOKsirVSxxI85eqIVWHdT+
zYRrjZP3j/raCOzyotqn9lREUIjacfSerfObjy/vCxbVXmmWW7l2bwDq/8x/bWP+9eAhbp/8WGTi
3lh+WHfJDGa+2Qjeva/p3Eus74cL/2HHelTOCgW5G06zLwg16wbWgZUG1mJr/VgywY6qw+6H7oKi
j2Il3cZWJNum87Dz0VB70ViUiAmcGbwzR7ATLk4VAhx4Qek27zgX0ho7DQEl/jRGLEl8Snbuga8U
Tp+OBzxBbTgv2M9gcTsc1JWEUN7qaGe6XTlrEHsjPbDABP9jYNxW460TVSO2iNdy1kke7PgFTLAf
K342sDJa6rVZmnz2qBGP2C76uVsaf+Nn4u61CKpxd1yn/py5h7VG+HGONAMhTCRYXCF0AKpFu5su
pMEXdgQfvRStp4OU0Cn958lTSgNFzsGiJ3wU3iwEmLNS5Ry1uYsro7e1UE0GOrFEzALfKHhI1yjX
L6qkY1k4p+GlioGl/xuDdtmc5f3XpB+caGwo8VVKInvzZcUCIkNP9FDLWjFDp7mwi+965XU2sAhe
H4eFDkDjjG8Yvk8cMyJ+nnw2foCbjKiTCPUzBWjD/9BXo6JRDgXEasdWB07niqxll+MSSR4Sn05N
pF7djD1OFVOZVSRrup2R+9JAYAfXLmOIujr05LBFm8bpk4G10mnUeEz5b91B44PwggVnSlaBgkEM
vV/1Id89B0oOFXbGUCIKb9on6+R4+UPQ2O10oa1nvSvuvenzR2VV+ne+n896in8Nx5RBeXegKBfb
dcGpvQo9PimhpfUvO0zmZUPtedYxpd0pw6xz08u/qY3R+ixbS+Q4lrbxiGyaNvTAYt6gIhrRxvFk
OndZJQbPQCZDOKj7pTLWZgOCjV8quUf41iNu01zjpgdPLYIwzOIY1OuBYlNUx9m4NoAsHxBwYQC0
ozfwwQ9LxKth4WczlLb4PWiuWtzrd2tGM2CN31hzMEmZUEm6VhJDKLo/igtW0u7BNju+Mts/3CxX
qFSCSUqc8t4Q96w6DqEU/RYKILigMWuKPEn8He/l1OE8n5qTxpOFccVGygEesWRnzUnK1naAjepL
ukzeW2rAAjG5e1AOfVOzSdxxQ/WCOn6HScYsmdTPufaf25cuGf/V+FxJojCXgmX1tF/RkVodyhBt
LiyAx8A/ewkS1KopcjQ/iJD8nZNc+JSMegTtU5j1+f1OF8zYvuOY3wetk8B7dp+5tG59k3ejJ+wF
SsQu6SI7uq/2oBIcUP/qr7Ay1T6ho3yINrW12zpjeyVwIHVcbvupWpXaWrZz/sPgskdJvmOSYeoW
sPlUrUMgByt4IB8JYcA8G+s0mygtNq6opfX+RyQ96wYF5OWwXy+GH7amp79t1zjFZBZG/8vHEU0M
2QuKRuphKDkV5OtHziL3jfiGu/e20OzjUDubuVT15VS/xFivuxEGFdXLwNmkjAqeiemkl6mjvxXq
bttfeTEEl7PkBUk0c+Ky88vYJCtW8JUQQ5b0sy80dPUuoWaiTzymVxkgUYBiL7UNkNwpumBK+Jo1
CAcGYBZaNpJyo1em+fjukXfvQP7u2mIorPBZNlulLRrGo7G99+0Pyp/kXUHdvP/Wy38QVNfqY8Wd
aTUVIElhGR+7nYME7p8Df4+no4cqokNqD+/HTUkBCgvpTS+CF4SgXlf3lvWalwiL5hctGZrinO6A
02eqLrHeZhNMDkt9Ey4PMx2SNVtAVOyJlGOGiMjjz9H05nwUwaLm88yJoJ9TxF5ZoDMWfXtTE6g1
yBSn0oBBF60tp8M1r6enw7GPt8t1l7QRX4vIUTBb4NxK7wV7s+iqcjbr+zxaO/YpDIriKHTNdBED
mVnAVOXxYmK2dntq6HATS60EnkStrWDTb6nWUZJi2RGxOMpfxJp3/O5l4PKH8FhGmVvolYR0m3an
nA/o+9YZCwuc5Vc+Zi0uZ4IqXmwpaPZjVclyPs8Jjr9njgF4qIxhfcMkDiCUnD0jzUNFlrr89WIt
v/YnlVvxgt79q2Iujs1BRA7m+a9SNbojgVK+gPgatWRdzHwk03yXZUUsUc8WZ57F7LUMYPw7E88n
Ewgg1Eu0nHPpTs8N0iBa/df6t1e/GVuZRcJOlwEz4CjDHcb+gAjlr5EMB3ITCCKeNxXTmGFTD9Fm
+chk7mYY9eXicVUOb57O0bU4ohAhD01eCoGRtfGsYgON38UGO9g3UMc+7vPrfkfU3Ugocc4Omsxt
PZqkz/MRuwtc/byJpWh0A2Xi5IPDaAIMPXjAHc1gL/QRm6Cvzn2Epza0ify0c850AdWvuL3+5Iun
PASY9q5ND5qnKVSrtQd8XY9BWbuPet5XHBiwdscLO+Z1toQJhGn8q7zvheU4whij3t85ycMul7Jf
UDyttUIoDtPFdPpsj1IUUOBv9dcjD1pECt8jRQxTYUeZn/BTL7qBu4SYVkUV8+BwPxHk5ZD6MqJK
oYJ5TldI4M2bH1JYeLnu7PD5Bls60He6adRVClEFxwi4bXaPXqYekx1GEpr5UC4kGdJdPeC70X4z
bS2g2/1DPzKeaT/YUFaAD8c5S/qLCmKOJTmtyZbZx/4UbEKbwD7316+4ZpJF7W1fVNhoK4nN2cjp
yZXJlzcDSfGVdAm+x6PRftvudPmKSbkglPNmHpmP6Ovj+fNdeoDrw6vMfZtF5U+q1jbdGh1CiIVQ
D4KaV+0RXrmwVnRzO5Oc0Z/6ZNArdggPSiQAZElUwbingT4QKaeTTbgXUMVmehisSDW4WnqFB10v
OzgiKIjaDerQPMDIELvnzpGpy9VEaC7VvhkbvxP6CvbCgP1Eb24Pn2thqHmBYNTsLHiHTW6X1tRE
vtwnu2k7ohXMH5hohz8r2qj/kjPG5GVL4sNB8n1kNS3OH+KksluDjA96FnsLJybv8D5RyvUo4uiI
Tq+o5xhnQxlyLAFU4uaPv9d/bYAYOSNUxPQsbifB85D8I2742H9xwEw54HVLc+WAiUj4kYRS1H+S
mhh034RmN7+VsrSPaJyvBwKmMdfj5RPJYfTcb2I7FeFWHnbz2tyicOdBIu2lSktucWaQ/kehgZCb
YmueFEuCCsBdQlA9l3liij7rlqYRWcZ02bsDg68o843qZSw3olunSn8bh9xqa3ltLGS/EgtZEMpO
QL64x89KsWAS/iJCu/fICKffE6qEXA9JD2pZZWYzka33dZfnryOMS3VuG5nRJmfE31PEZ3Iv+tYK
BdAJw4nGIulUAM1MuoECgeMliOBfITQ3LOMZatv6/ikCW9bwCsJ15r75EPyhZhFY5LKqJpyx4Z1B
BxxAfcdON+PS6kysPxLaxuY8OHOcc3Qc4mCvDSrNdqs6WroK1XEj3l+N/1sMNK9nLSTPz2Lc4XXY
qkNsdKYxlCiRAO5DzqnPcKRBA6mzPlLJmxH9H/HvKnVYGfIagXEjiZXUoF4kmSjeyncvlDaj1FzP
FH5fO8gU9QXvx9zXSjeze5AOG9dZeCTtmxG/2TkQXwIHoXaC6YR6mWfFDak+pmH6yTF3CIAMPTbD
N4M3BHRKFc1nQa+WhBTqrBuY2R5vLvPmVDDEqfsHeA69bk/EEQQjjQn/fD9gVUVmW/g09rlyPCgU
L3mgV/dYkTFu5hJRAUCC2koI5ApY4jgfu7TO1RGxdVw+os3uY6Aza8nViNZud1ymECLL5vWEK2KH
v0GKPOWz1qlaaqdTTXEyKcVZ0DImO1UdPor7H/VRz53X9HM2VSTxVe8hYg7FDY+0+UfmZxGjSm1f
qqb/hJ3isjPpytZf5O/1LWR6cQt/Yvu8E+DTKagbGfaQxHy84cz9e90X/YoAkkJg8D+2VBUSrCnh
1FFQ7axKdlQdXiJa7VXPQvEjrE8om1EipHx8Z2t5QBdWTtnqUi83MLniqYU96ObrJHLBkOFD0Uom
O2TN45fS+gYrXtgOrghPO1D++RNNBGo/2MlRVlPF39zJHZxJbsNbBE2xMxN356WJSxdTgTWKN25y
/xpH/l91Zuv30PTECLP4xTMFeL45XsJFdk7fidcbu1zN4FGw31vQB1yRT7zOJybm05qCZK1kYeLY
RKVZchUiox5bhCyZV6OcYDDyR2eJtV17PpAhANJRCj1evogzgPkPiQJV70hgclUivmZBQNioHpZz
RA9DpYHAUECaaGrHg2wF6F2XLWpxQY+c7OpOCvDAbU6V4II3ykuLu0S6cgMBBLSRszdunqp40tyH
juOMR66bR9tFK5xm2Engk4BTuWfC1WVKXWFNA+bQP7hxTLc2g/gAY4JjnOdPID3HOCyZByVrbjL/
zBu8RoEcoKmET4uR5jtoNuPPq+gLrcFdpdVRnUD0tG2Duq6iWP13eenflYlqWvcMnZIU0iP0jLke
GJTTTbjD9ahRWkASbGrSYlGMyRMcLGft55E/kBxd5mud30sY4IUG0pdQV8/Dx1JOL0JHooEaCraL
nU8LscKZe+mqg+cmyP1GSZ4F1yf+6BlB0NwKcnKY2gDcJHFFJrZ/C+rHeLOS6wLMhEWVXEXs3yVZ
bEFdH1BTjiEioSjcE0LxhrtO8xheo+pPS9xIugb9E5ygnSSimmYW3BktoXxj6C5speJUG0Xi43Hs
ZnRC3n+yyCGg2LLREtMy5+X9fn0xVwazJdI9mbbYEym85huwiYJ6CMOHtwIQMN9+UYMx736QSR5k
W6w96c9N65vYaSV4mEEWPGbWmGdAZhbkag2A1BEAkqsaDf/zGUjrf2bjGVjo2fg7/EqN0GsIJVPf
AMOkHxT+KIoABsuwLF/c8mzh9kzwui3mH+YPkRzdd8FGtNgULlER3AsrFXZ2VnbAW9LDMEoM7vlR
WluUy0StMZYUbpnvCPnrcJV+WvRNYOmPf1ed7FM1tnYDIBQrw4csM+7hmtFalfjbR0X6XsObcfay
99mSWr5SaSLigVxj7MxzZRutZhAyEHpBBbuKzpyV/2/ZxA7mRsPPvO6g65y1Al7WrUsBBThlNpKc
ePg0OhtxrMqWDs06HZEZpR/Qg2kejCDR5FpwQAPEKajJsGsHnICDGIzfnH64ZO85H3ekc/foUn29
UJeVVx7sIsMk3LysnuTTBJgYDzqic+yArKIvIH1EFhsA1yQJZ966iNCVuGrWYxnV+CaJdlO3yNh8
kRJut0zbN0TePRHxG49KT5Rzf0WdMdYEVXf50dSZJZ0ZiiE8/btUOMI820Gauk4YOEmJtzpgsDAM
K1hnYPFF+sQl6Bk/cjeJ91Yeu/D4JV9IcTS28Q59XKV+D6+7cDUgjbw9D/1yibM9wfL0bU3g0ZEF
r+E6i+JkalXKCydHkZeZiBwFEGO2caJTb5BP9DSboAqOXD7yQuMBL1tqhdUDYUH9S24CsRDkplMJ
vmcUjV9BrIICO+J4FVCslt8UY8Sxl6Ql2/nJ/i4nxUwqbpURAiRkXAESYfu5PsIiPEVOgyjYEFxx
15NBujord0X1iGsyueUsNp0X0QSH2ggmCvd+/O01c/5CJX+Or5mSLEuqGZX9ISHAcTWs3ShPnSVO
Ozb7t4ksxko83qROaBWTQcETdw6tuKZn0I1QT1YKvhUVHSozRGqZ8SGZsTV4BQmfodQPh6khMnrI
3CdE4oxaGdDWfYnEtn1blbLi7zMelGhrRVxLVg81iE8XV0w1QNcm6dXkKOOPSLM8EuXow3wg+nBC
fPk22PETvuYhIszxAQzi1frLylp7VpwkSYjoXk3tdtAIrEoO+gdf8fba5Dwqr7QbspCERDD6sAe3
fbxHOnKyCQMOGUhujiRGz1SoBTxPBJClvp5kAfjWB3l7wB745FUiMfov3R3F2cvzCcf7OHbPEH4Y
Rj/830oPy5w61taEthB2UPBPHrdmvPASZx+z1utuNDnx6iDa5fUBV+ofKFvhrhCGmLBO+M5tXWQN
z6iMqmDSvoXmFOXw46EJw+5jKpcX3VIYNMU+XIkutK+HRheKJ0a4gbcsKVcCa01apumrDlb61ppt
294gbsrdZpId1mHuOD7iP9eN5jKXQEHyjFOu4EM1i8f83gyyPORECTsqKEBzJGsVsuL1xrmWtnx1
eF5JfiAZ2M1vqZWJf1T40hzNrqg2z7FnpMlVnXuaKrH4UZZ2mxzrqKjJu3cxMH+JvsmbNHJ3bOkP
E9Zi0c2mx2W+LGj2kYUnubOIIPWPGzod8ZQ+ZFywy5uZjIbHEZ4bRK7ID6gBa6YIYSEr9N/sk80h
BhhrMiEwt+5AOD08nr/mOIptOMap2idTImYMJGJk9+B2obPN9weKDpMFBjXMh0JQHqN78+GFjDqR
8zGllCMtVjf4Ec1jpS4jRPeQRUtEF2sHyjGpgTlZs0wKHmCkJ/uGhIPraUZ6d7EsWmaY2+v0GkFg
jMRyYU69+m4vtFoDY0j7w3B7SnViiT8rm5zjKAGp0JsO3e/ci9I+ZBC1+bq4DayzXja4LGj+0fmW
r7qUuQW5ouEoFDOlnQ7QyFoOf9Ha5hof9ZMcDKDF7wfXyYCxg+U1/6at17ytTPktU+SyIYO1JGs4
+U5Mq0NafXD4mQIDe+bMuRIvmaGIITpPJEHLkBbP5ZdoCr5DheJodmRWgH+nEOKVmVNWC7fwJUd9
o5anHBaOenj0hGiR3RXrf+yYyHKX9uhnSNDbbGzAHuxyU3IjRfwsDvGS93sv3uaT5NqLRBQslsNu
+hU/2EgJe6lFO0MasTCDqSgdo3d2/qForxPl79j3MG941/Jr96oAQ0aVn/4+fzBxx4qWQZzgx4Wi
3PrR0oOPNiqNdBshY7FwgfgXIclXMS16Xm6QYRacy2FViUQipwo47v7UNOHse6qqiy2UqlP/52uX
HkB2W9yAP8F9/nBV6kUARLFnZjPLzb9KWzN2rD5OzLnbitCNBL7qYb2sNUjS3Pk4orY2RMNJAFkZ
OX9hwZgoUGn2sM/nDxvEQk8XjQ2JR05V6g0cuk5ibP4kR7qqWKTBkKUVA3SCVP7rcW1ICrU0F0qZ
bPehScpE/jMESyCA42TJvk1PjC5vuJ0l2VqcIVB7i7mGkWUMK9mRLj1ozId7wrSdab6pIl0NTbkC
feJgEVQAXtFP5GQOStUpJk6yzLuX/o7Uk8uFOTke1CrA/0DGvnQvPLUlIbof/3B6J3mtsRH7kQTB
W7fqDlhCW3OAEnW2uwWvt+ZZ+uVLkgsvgGuUxtzo+gdf7s6iMHiUL3NY/LxVGrwKRepw2RSB1OYD
GPsn5fsUMMGNvIGkhlaxTuoL5yjbjdXjPhlf72NRSt49bxHryNJgZIGvf877sL6pAFvKl5QCe0Q0
IGzOLz22I1VI83j8FJ3+X9XiXJcMhoQdROIohw4hvklGe2f0+MnYLMPAP3ZUzDRF6s0vlo4zdzl/
iJBOp/pwrKKYhKk+fLLyNP1lOykT9Tri/HMUTlUORmWMO+iSzjZuR+ni4Z50EUnoq9bQk7wqmV2I
UrYv9LoJTtmu5jxcUoLHsoHcD1FWEdFHZcG8bky7XIUzRq1a6F8LyLb1ctijhP1+B9DceR3EGkcz
BGK0HrgulyO4eYqClNUv6IR4mhn+4FYfYWFEDIzgWm8Amv15wU3fooTW23OvtBK2HDCkZY2USeKh
rVXrm5sa0F2dG7KDh87qIZSoqaYsgH7e/jDuv/pug4o58SNJS8uz659mzE+V8g4Lt3tsJM44bq2A
kG19wEf4K7eJ6rM9krtA7g4DDdHjz3ViieQm6xN08k/sRUwE69VMwwzu/zMAz0LwVtRpyUSUt50f
os79ojX1UxPqZ96HFeCcICHq6sSh3ouw917T2hmTdz/2sugCvKFqkvFtFtfgxZ0bGm/qdlXs2HsC
xnpOuWohVmQzzTUcUtYhSZWlmRMBvKROcstoa+TNKVElq4hZi3g6wZ4cZobS319IojCEhTYbfl6w
e4IOV9bGNqOteGskNlUvI88VGUWYDz9d6h0Hbo1lxrnewcxRami4MlbuzYbvdfOlwOsWEApLEUK2
lKBKjGAXBNh3fpduzWdxDd+RRiOeUyzA3JiB9uv1lmF9K0T7nG1hm51hn9nFpn9q2B4B5xKv1sYA
WQHWCmCzP2XE7fV1+ENa4N64unFvzto8lBTNxPckWnTXKH7QF9BCiWiAxixVXY2xrMxVVS+j9R1D
m5sa9l2f9xp1Ane9pHqwaCW5iAG7fp5x+kPXUFBua8KU3wcBwLLd/6DHUccbVLAtKAgIOALMGLmW
2ARwlarggH08abqnngzafv+koBml5QejwQsRbmU+6e/JCCfVfPtFYMC1c+XJMpC9xH+bTSNQs68f
g4b1AgQTCZHhQqcY9AxyppoiJKFqX5gzVX5UuEghMmcO4AL7e5Uvuj8z7ivLxye5qN230Nn0t44V
prBW/qvLMedM5KFN417JlTPoA/tv+fYIb41EV1ao54Jt5Jlv4iuxN7TIym3ZzTUmyeNwC2jGf8/i
NzZhuhK0i8hiismngI6qpHk2ZOtkrCoEWIfWpeNu7PFvkUVNQ+7/2ocLbnJwBDv1JFbquz23SmMt
UsiEfbR+nx2FH5sQRD7HZlucmpwYUJ7DsWlmQR99UKbvWqvr0BBGuS0S3v9Fm+boW2osR5qfAuer
06RHGATe5I0Cjp4HnIjuv9Htcm8o898FzIAFd+7MH73DcDJ8udtrVQcxqDQXyFlymSdUnwBZ8a6V
5EpcdAYXdRhclbV7QAzObBzaktBBPSq40P1tL8RwWxnrc6A4Mkdd3W5+poznqzkVdD/5ciuR4K7b
OQjnQ9JWDlmhFT4qcsQk0NHH1zvHxd/0IacBWQw3h03d7sUrjMD2bgS+ODCEVRD8NapHpuJGa2E6
7735c4ATD4yNk1V/h9WBgDcqya1OtLnigbKuj1bY1JFa085Y/tO8vciZI7Rr994Ax+biP426f1aR
M9jPaDmz2XaJ+aewOsircSPeKlk5KOb9rW3ox19t/19bu8E999jkhJdpzTyq17kse+r88utyuhed
ww5zlpweTDb9NAb0sfI2LTWZH0jwjCGDTiMTigWGbYx848x7sO9LrHjbkFymDiyzXSop9MeoFHoF
5v/nOOTca4e78HdO1uT4X365eJzdnBF2t9+qmTnsENvu/HBlWkSpzY2GvqJvKft+z5NU7rRuf49P
0k2cXJHyYk4JE1aU16qaJrGOF4LXLktxIH7Mu4nZOvrUOkWJpz6x8ExCq8swYHTWeFvtLnvaUX2v
8/PhFa1s9xE/tYSDbdJc9E5bhpLro9HT7IGFJsKKhaEebkLMmY0+OLdU8DmFsFyq0c6MkF6RoocH
vn73ZopYN3di0ygIDyVMZ4Cs+nt25AU9LIr3k9lKkdxHBfkBX5QVibzOGBJRXuAI3LZAy/sjiBX7
ebdVXamlTvvup6I0pG1B2P4WNzBwJz64KlUwt6Za/f3QIcaCdHuwmud8KzV3Ls43CHpmijoICwNQ
uYWh1agadGkJDuKp9SVnviKvHN2A3DcbBBlO9BVegfCD/2YEhYCdRZStVXytVAADGR1HK2dBnKRh
Mzw+sgTOz1xmL0Q+bavB3YT7JxZVQwRUgXcCjQhI24WjHDpNd5yMzaB09QkOjFJ6HLdpToPmguQI
vJXmykhUEDnpk8wvWHB3MbwGUM2gIzQhXlGrxljyClb568cgEhVh3ur0EkXive2h9Z46SzB7LTp1
Ni22V5I3E9C5ZBkDcsXt7YZVudONRZwMa3xX2tyd+gUtPhDwiJCAYjRXh98R3gy7UEO6ThjAZcXg
nrTTmRaBYSc7AaS6Te94X8+KPoBpAzTzKpFTUNj/f1JP2tPsXrXv03vCAKEeYCrtsL6RElRv0RoF
nRR1CrRErJvKXK6CCLXpKxJCFrzepmUmEdBnPkatDAnr0FM7QJ5VhgKkwINOzno9FLMkrFCyjLyA
7wbbOoOtueTtViYWy61faHRiBFFfchQ6ea5LCNavwJn2HjCVkc3pzp65oVXga/naSrWEqM6rZUZk
Eq5cXS6sQOoy7SBznlAcd97orR8ke4/UmwMmb+1Vu9WxgzlVzhGWPc4gFn3bZP1pN7MqoSWp4Uro
QHfNWlao7usKCYi5CTe6uJ0Slc3Kqtwq98ERHNahcX53V1chRMvh4j39tUm5zxPL+uzTCXZkgEh+
kly9BTVm+v+59L4a62M3NYiOsDUgOe+IqZzQB9NaoeGWV29NBOy3daSWgOv95Y+aFqJlV0TtYK8e
lBmSIFsY+UnQU5EBaXvwjV/ECtdkw7EhrHgFF0x13nf/yI/xTjrMYJq+XR2VB/Z/F6FroSH4x2jg
TfIrc3wNAUONtXkat5goewHcQ4dHPBFLFMlU2KpmLBokHPO2ml0NqOFnwB4nSutLSCD0YKhf4//R
E9E7KYs2AcB39d+tbZh2UZV8AdrXsYKy2xIZpQZlOrfANaOpJg/3tOHEFSje6U6L9qjS5nvsMhwC
ARK19LQ60D3z0hPsQZiTm28Ah9+X/fIJOFk0jsrxSA60E8o6pq9qgSOntiKaPbSRvh7OCO9xbJH1
TcXL2P/m7DpxXPjdErOYXYuAUmPEnipUTCwtMUhrKzdG6qaFvqftQJbAqs7BfkhDJsdRxueNNkid
alGzRbPbHnKVhi3TTG8Vc4XPFkHDUqtSzvyV2Dz7HqZwWcbVLTMhUxXlCa7DMqTX1CjKlGPy12mQ
vPLyQ0SKnAGGGidR9PJ9MsPAffEsNkN6Gpph2Wpv9mZlKpKs729sI/UudmtWBhYF4NRlbVwF5JB8
w38Lzd2LGj4crCvBFeNuunl4wtiVNulW0GSwVNLexbSiGZSkBafTOwZMr+69H10udeX31+1D6C6Q
a2PIBvfklINMTsY7svpy5IxARUHEoBh+vEVOl4kOkh1mInzFyZ92K3j5XzTzX27zlDzuJy1ol/Vb
cqFt5rtPt2Xbqguxstr3JrmUjE9NGmcVCV0Yob4g5QRX91TpBFuk1N2ejVh7AmoWI8O7r4JIQ5Ng
+VvbEa/9eqJQdjJSNYn9NDXeez+3N+QWkL+xNIekVdtt1Jl4NZlnuP5nZ1owaltSYx+3bBjwKFhs
YpSk77cioXjqip0TTze1L7e5xlswgFKyLqPV9YksoW0/t5CBZfw/SzYN501u8H+VtmCjGTBS5ToA
gOZaTCjdatRacIFRcK5bR/BhzmgFCCtHaTCuND5zPLvRCmxC8YrCliqHlNsmNIvsLinMuo/KY40w
hkcJ5kwkDReaKDIL5b+dzeDLoTlCmx+EHgvJ44dp0iyIxG5kI4irr6MLGpD5PqvLwLrJZnfIgRef
rQUhA0XgEMOXt2gN1w7XCFnMlwdVAeGsng6wL8ahF6/nGDJDaFwF5IUCeR9dUiWboM2rVB6sVo8X
YOtG414YO5JXcc1bDIFArwHZciwsun9oWOWyMXydSaPtXNin1wTsmLlGJY6YGJkA7jGfa2wFaUfR
NRwXr0ifUZB43hBvHoQVbyEsh0UVGzrecyZsOB+JIyb/CcS8S4zzyzrNxN/qaWTES+h57t43uTb4
MOAg0M//7Qc7EYniM2OR5ieL7rVkBvjOn6ZS48YrS2h5CyulJnTk+6ji/fTu2Sz40GuX/es4Rv2B
xVnY8AmKv6hzu9G9kDpuvhbs/B5xliGlNsv1Yi2ddLRNic5pn4fXFHtMHJ7ML1AgQA5rau8tRL8z
wo7smqEiDe0Zky6qGM6+NiAgUiJVDdr3bn2hOVLWFB4fqCAwHf7zspj4plB3bQBxlYZlPixTO4/1
9MVlJLwys0NxxVxaK32D/NUUOJcIOakaXej4S8JgJmhZBZXIrYBku54r7tetkOUFkwMl316TKAZY
u957rMrwPENCCcXnr+ss0pj+UxB6Oskwd/dojjNiHRPO58u4r+3J2QMihNQqbDQ5xmGpgum7xEyj
HCwaptYMB0Cnq0rkNUtd1WWdkfqVxmmLfG8HrBzW56jj9duQssX+EuTiIuJoxJc5if73tcVagd+G
ABXiweljLhsFOR6AkEHRUpa0jwdsRz4Fu+x5UrajqrVaamaZMwrcqyiHHv+nxUUO8oCoowgN0o4F
8+k79bxxX3juubFvcLtKQMFEMCPmYzh3zQ6D0oWAq2zqBuzIJUn842GX2LFQTkLI8tYm/+NdtKss
DP6qA3Xh390iMQ2dQHdfvCYvbQSv2ww2C030WLFvqUk0upEhmuAcB33/JmI1DpgUCuBEsdRKoN5+
xrmf5U8NQhL8Ac9m1sLKZ1uO56v2AXxYxS7j1rSqQGa5X2o5vTxDhuZkfpInJe4vs+Z5K2DLsypu
Bx2S5J+Pj3D2woX20m1mlNKBdCIhQnaizvK9wk0enEV7SLzz7vFZrRvihCdpoWneoXGAGuHh6TC/
5NAcFD/8ScJ0xWfcT7qPwB9ai8f39XqNpOv7V7FHLbetQ8CCgDIxLUJR6zyC8oqqdL79tT4mV9BE
9YLunRv0uuznwBoDHaerwFcN+w3dnVdWmA6q4ny20wOrQMlnHQa64dNkxVu2v4JIyh4Y3v2uRIqU
krlE3D0DDze9zpT9dkHjQJCDd+ci5rX/hcNNO8OLrOj48MWDNFRjQ8tt6TT3Vp+PAyGpb6kzLQQA
4Mdq2bcN2xKlq4z0cdhAn+Y6Egs5x+dS0OZybqqydc+PP0H0S5o952NC4q7LPJL9eY4WaYVFaaSn
HCQ+x5DRr1dmzhmu1C4ncAXGJvX7zzxhbGFWj0UxCDIF9ixha7rohJKN0kxIqIff4mJEnMDYhhmP
VfvluWtPtytHFfFlL1TQdU9PdpjvGWJcfVaADVJt5RNkdbTzzLEdDaiIL0gu2D3f9Rx+0DfWlzcA
hq9Ril1IoufPYeI7kEPPoNBGbdBoYGyjqqnlqO/GGu1ym72Lqf223JH6a+5YiEkF4TWrURASpSt1
SmNGsFQpw93/VQdbmyyiJXr/yf5pXDx4Ln7pIp3pg6gnxhWAeMJCBB30Usvejfx2btwaM4Mim+qn
S1VqoqXghW3/UmurwlZFgZjJ3ZWAEorm+HiTC7jEacsfIuJ3dymEQO3M42YcoYHYgEfP9s26N8n7
Wl2AXJzpWit6R6kcQCsxa6qvM3+XMV7EIXxk/4N7a8l7Q2eyQ19CkRcThphF1oHZbafkf1p7MoFS
4TDWaOmXh2VKugS+Qx00HeuUqPSOyayEHR99co7n3nI3A0//jdxQTDvs+eTvwbwtY7kGjM4sxGgu
UxHNfp0q96urUSJf87Sj8/SjV1AfXe0xQQ6DpIbk1yeOjyj0Hll787EcQlexrbLL7li5bkyryaCb
9RBsZEVWbE+W6goprBlzywRUQIrAbinOjP5lFMpAublVqy0D3kDOaaSE6mD3WVxnhmMLKgduj7kj
QfokRswK80GXgge9Icw98odUsaj58ncUdBmTndROSQD7qEaADfyGw9HT/1osEa+cFRIKTK263mTu
Q5E0VgAXuJ+NZzFgGh2U5E/bUTeWtH2pqMoqn+qHbq8pvoZw6COxWdzEByJD7MlzsDY8EmUTSMC1
tbKi1dvpLOe6V0V9QjhAaFo0gN4d1/WmC95qTLqfL5B+jipULraZp7EeLoXr8anE1wORdkuZpoci
DNAongpdoqOxRQyLxHS+Fpp/DrCImC5Edmdv9PdNWgWcGlYrD/7ry2rfAQqpUaZVcD9c4HruMhsI
7wWxES1TaB9zIu3bXwh94bepOhySpkQ3HPyKqpyz3YHC8hSqq8hYyLOHqAPAIIo5FiPpb6Szy/fk
hyDcIEoJ5jqFVaMea1ULoLBHUAEmjRyPEG8NVgnrBp7FPC0pItsKyRWZiSLlV6vLasutmJ5VvQPo
DAl/tw30N3k4opVOKZQgkg06YlOkViE/uqIY3MZzivGHV8IJ3fQz1gxgFPkTyPwkRiXGJYO2SEdc
c7yq1Tf+SxuZETMaaGUupAwMlDBqziS2vZWNesnVpJt44MWViF3m6cPMJNBDyeKf8oJMWbNHjVWw
1seMfa6d62sNr5w5ipYNXcTTvJar/JWPrHizZfDqS9bYBEvXFNUIu0u6Dh9ddYmvf0OatnVxrzmc
oUF1Sj1FVJdxfRCSHw21ikmP0OUfxntSdQsC0jeA48jQpq/dW2y8MaJad/2XN294BCnd1FLE9za4
SuBSg/nzy1QesGovNBwNbNK3saafRTUlWfBb4PCwMiorzLodgKqw3lFEvepFl9f4upr1la16rNYn
HjzZg7ZOUMQBPFEGuZK94ZN5ba2gnBLRwQQifr69S/+OtFSRT3SPG6sYTaxoXdNoUTkSWCIrQ0Vt
yLoaFeWutaUY0ptdYoUbgj/hcHHYrrWIL4ZO/OnKbZ5Q+DUFDSxdXzApvHYZqflKp94ET/ui9xmz
roOQRzPTTRuEhm5VzmeanLgbtoMPtvyNp3KKQBttn5k33jH93DKB9giMzFIFvNBVSoCnCePi0IQZ
HtSEz+42U1vueKp7aHGayJ1aTeqs2Qk3m6q+LeN9F5J3OTQBG7V8qFPYsJuk+mWSdz7i3AuxLHQm
g4cDjct1uyuHhYVK4AXLwv7lLOXCdpWW0R1MBJJLnIJtMm0icUh+3BUgxB6dlVeBV3PivD40A0/j
JY71BuV/RzEpVI3qPzmuH6/Zwgv+73lGJkjkT95YBLcwN98HtV7pMVRbBcnOOgx6LS4oeL/rDC6L
L5WxnYXQM0yRzz6wsfCbt5B6J0AiKHdK/e8m3McFXCsYZlu7zHD5Ge7LtkUKp8NYC783hMDQ1qqX
PrEEEDka938rkD1MHHF+Bf4VWL+z06VkRk8sq0BYrX/DykkUDmmz/1LWOqqpTZGQhcMUfz7/15+J
6/gmPtSgvoSsEnDl+O+Em4QPFfHzDueTuT8T2dYQs4EH+6vHvnfylCDxKqmjjXAUAX2ksI3cp3hH
Dnqa4crDxsDcFzBr5POHaIS9AQVAmuqAzsVG8mKv9wll2r+oaGqqRFextj3qHPaxekhqEiNRcqUT
bsEHnRiOiaTuzN0EtxTbKqUqk70fM/RageU6NzR1Lr5wEUHqInS8Wx93En1KjFqcBkzegs2OQKrI
yO7xrsQuHEVPwGIQ83RSKmoWGBuVB4afnGSeb5cQYBtxtEADtOoJxVCRwxV8EWWLDJXG5wnFFAlj
zM29kj9gGjne85g05xyoiur0yXDnl2SDS9hf5EBunjlbpW5HxXSPULze304GXgwcO+CgLQmF9ChQ
7t3wa12x35BA7TSgp4XuHXfzREG3Qi4R2jS6Zc5KaXDM+8hD0Y208ERfsqHhbBBunGMgqO6hwM78
OGPRv+nbRzBZtKzf3gwh2v/AvZIDthK9IPG6riF8POXCK3BdovmS+tjO4y9IBpDeYPdeRpEU4y1G
/b+Kc6Rni2lpfZ39SlRSvzIYSjzZ2hb06szc+Z5fhyGlO4S76fWzcRoByNq52sbUE/+h+7zZy0YM
WnvDe42Av8/MnVdB37aWBRuHbC7dn3/pq6JAPCKzbzjpp+sPbyFZOD4XsTdFVyz4MGlOi5VMHGDG
LymDYTF0UjG8ziCYTFq7vjTFVv+zvOZZBOwvRzRmJ4DAVF9tB6Ur5zj7IoZHhCaKrXe+tzAb/Opn
OKUNnRgGRmIRUAcPZehpJmnWtb2uJHSAncm9iXBgOQM1a4aCUe7TwqXVL2q8abgDSLSfvzE1K7ko
LeqgM7XweZVc5o76ohmBtS879Wzu+j7L34RwSQEcKbYXx20TBdJ2SAcqC2HvZsLmAcxCFvpIzdXt
GXk2NiV0BbWu59hVr+IbqQPr6noIZlNsRvsU+XPnWAuPq3LqVzPgUUQnPPX195XSzksNvmqDmyZS
Et7H6Sp7m+4kAEukyLQ10hal3QVjKFGRFBVxZmS8DcRgfBpNQYSfPufN8hsieyC/J42PS6TWywKx
ug1YwR8ldHPoDR5PlxTold6IjdamsO4A5vVmcY44uM+Iyo5C2prwRh0LeXhjzSTb7aHa/5LumvKM
U5jGeqapGgDB33nbJCGlU+/rFd83ulCo/9LLlg6FHeJixovTygSbUUMKstf2VOiezM5HLvOlO+p9
5GNIYIcNUM6eCrk+o5AdxFywb/ISo3YG+hnMtosDdmmfwph8b+fy73lBjmn8fvd+YqRmwwJOUOWZ
ZQ5wUOjqZYXxfp3/U64ehCx6UE024SaV96ZqHQzUL92vBYB9AqTrNPnn7Y3IOaHQRv7zsZIeDPuq
nRInKmPdGL2O+WyNrl1JEy7k4H2lhZQzGhdTqCmDj9LHk5DRE+P4PywOXetnkvL3bSiMlRM3RiOb
qIPw4Ga3FSAu3Aq4j7I9x7FV42iQQRdcCVebEIlQvv3YLLNQi4BDTIxD+7kZPUPXUSNDrLdUAY4v
/4pii9tD80oB7paDJMhdsL7m32lYNGnCKLtngbh9JJMz8/QsQdyfAgYmktWDZpLpc74lrCDRXeZr
k7A2guuFDis0ujNSmgL1LnCQrFCT5952qT2pFdDmNW2m82SgowyiQnnOeiiRBqDvHCA2/+ciRiLw
vq/2xh8xICZ/jYNDLSSyLTGGOer+3IQ6FPHq5HKyzf5FOgAo3C1MgyZ8vvaUfMRMxA69u826nk9k
gfQOfc4BLNgp9zTobjAMPECkSLSwg/RA7z7XcLM4ywX1TbYD51x3h2XaPHN7EiOt6ufZ1YZhPxdq
C6lRvxwja/BLmwWzk6uQMCqbj1AUOXq05po7to5uB81ltdpIWsnIZyEf4smsC9icwb69DxBFnhTI
tyekscdf6UO8jiGTPqdj6zjNade8ccS6jbYSZt4DloB4f0B32qjidBQjd1/AhqWZOmrA1mOp7xYC
oYeuieAHW98Dkoy4c+aeh5TqhdXJdo/vhI/dUAvLF6bfhGJKcRnhOfjsF1wE2rMxRngiGjSegLAo
gNBinxeHqnsBGYulV1WHE/I0D+pJTkDTNNa7LEycOhzowQtq5PWCl3GDzjQIWuU4KD94WwUdxAS5
RDJC2XRiFG9nDoV2N7KOuA7d0YIm02M7CZq7/0Z4M0ex3FYMjaA8WKRrK73C1dobBVQcZUu9xLtM
q8SdWjKKJ7oeISN29RG09NSMF7yhSsnZ5vA6f1kx2eLhKe5xJwDjDZRd0HdujfPXVzz+4f9o4W0L
a8FjIkqj9N2lCiaCJGsK4voeOyCTrnzqLmCZeqp7tOwYEOGoU+WlT8tKGA/1MnTWnFShadrz/uwC
K++6d8YEKdbVuJULHjn6d6dKlxb1ORuhVgz3jWV8t5x1AX1VC0H9uCtJw6nSd52id3MPbuZpgy9x
6ZUNsJW0HBBfhcVM4bk/VfSUIE1OgT0wAgLnZ7WUTpikFRIViFszMkPeqAwrZxM5BhX+WMgRECbK
FY0de7Xl1GSQUifoJKnipg48A1Gko+nqqtqfM9S/qH/tkgLlfMg+OO+Q+9u0zpXanqH9QLhf97+X
wGEsWTmlQc+n0rCib70HhtcuSVPm1x+GfuokjY6JefR8AruQQImTGh/MzvBa5zASoBmEDcfzItJ0
AmqRcPbPntyZ9tB0VJkm1USEVZkqRyRr4a0HMMDWqioragiWiElI3I1FU0+9rYPqHD8+PUPWhWTy
Nsc1CQ5Ur1i+fN46n0WgLto0S0fnJieFN+WV63pKsmMDByqKtK4w5cux50IKRoRxSEs5syU5DcWB
zD+CYHC5JU2UI+Ns9rl5yeaKZuoVVXeFyqB4X52CJAEf1TBMvW0HaRjIz0JozFxYy2W6kLJBDmA8
CeTDQO6mLsbv8RzWXMA3Oj7PoZmQdVVFDtLEoTvO4NOLBm+sJ1rf8Mun8KXz6EkAW8YHeDZ5mLPw
IUymfmb8PM1v2xXR7PBXHuj8lqvNf2PWXqXPTRTclTiPr98uvr+qsgU3YTxRVGbwe4P6NUhAD6/I
yRKkRfdBTs/1WV0F4mCFUxnKMV7PJJAbrT0yvjXlWYFx3kmA7n3MewEKPyqw+zJQYbP/AKKBYfz8
Luxx+rhDLrmgML/EfgE1wqWRt0IZz51jk3nEc1GLXf5r9QtBgw0+zT/iTo/QVvWl2p4XVc9hRbFv
jrLADZzTi6MlXvch1vihQzVEQixf+x0A2hWLmpl5Wfur87IqcoylFVIyMyi2uY5EuGUX8N/GweYj
Gk6uKNLauVIr7yaSIjXOgkoUCFK2+0cEGNpS1zLFFAINyi/G4UmZqgSbAtuKZJ3Cy+6dcNFkNQsT
RiOCD1UHG3tOC+60ZP4WdIlY3wOqjVxX6Y1PFdyboNA6scuzpf18Ql1JvWQt9d4Sgx1vHDCki/D2
tjALukORLfLBPeD2hGt5pDoq0OcnWQRr9GShkVXRBZy9gtB9X872jNPrDKOszeQAyMW429cN5kcU
cqSxCSSxFNakwW31orlLKPh8yUMJTLGd80z2IvH1VAFvSlVYhs2oLoD8m4n6XCWUrItySjXbk3Np
iTcrm9jDOX1deSb7ipC0Otus1MB4ZmrEWRDpH7KdD6weQ+W9LikoC3jl5lxUhILFXAh6QZHwK+3z
m8uAv3DXwyEr6eLDyDjvrklXgNq5zau4DFYJ1S0tVSIv2X8Pu98luarS5Oxzsw2TLW4dGEvPdLoz
TR9KoxhUIamgLfxtWt5G+cFW3TzKz4bjvzy/9dsMVarDaRTLWKPbYX/JuPRIU3I7E5oZKDffuYBw
tipYHp6Mf3prnNTKaqjSPQcQnZLpEaEu0ujpaOJO2M4T/K1OJ4WovemmUsD6h5EMybFcCYeua+fo
xYNWXFvmg1IJIOb32BV64gs3tEoLkjusgZBjs6ECMBUkVUSsGH4r6on2utHiOP1ctzTMwh3LWgwI
sm3XLMPDFbPMdv6Zag5sHXNG3TwGOEuNaJVDTr7aDMyzeKZGo/a7n9DFMAZuoaMGO1+3j4qv31i4
qJbA7Jg8Pqk35QctxhTwTWGOhVQz1092YLFOlTgVnQ51/LhAXd1yOJJERQhJT+F/U9aaM08pXnH6
IDaO2En+OLpjK88QeT4DYTwnZkPAtIuBZhdGxCEIzVWX3ol34x+pPlTJMfRd5MMtQ9FLXaouLpri
B6L0d6F7OvUoZDQiHSoBRihximPjeYQkzbO+j/cewYT6TsbVtLFtJIP86s5f/gRfjjbAcAkoWMNU
wGpwzyq7m1vuqN4NU85I7ED7k0/H5EQ8ZkkUEK2y4spKXuwfGqpPB8pvUq8E9Gsq3q4uDpXLFV7U
LQ9h/F55urdjHlRXoTDxkQyWv9OMZlGW/JZyTMlZYMDLsviL5ZqCdysUdzUq9iBVOzy9aClDP2C/
bOkQy4HofF8hkr1OKE+5tRA89LfljVKkJHMkjqe+doQGwT/Nx2VY+LUzTq5kWYZUSsqacqC4zgck
QhHDWd8Rv87X3hEYekHqWIjRxDDp460XjiDc88mYdCvvXroCwzynOJYf+MGZbgx833CbSFZ60WC3
o0QpsqYp8KNyLjNuyp0O5pfWif6e/MsI0h3HRuBFBy58/DiKoUz2C3Xcv821ONQZT1WFBm1e5KxM
RsDvFsEVQ0J9xXwMkemvko3KziNUKgUXqJfdxPicl4H2MADtNrfFSNeFMBMsA0caIFIp1FJZSI3U
mzO7Yi9cYtGhQcq5bdZhMEXaqIQS6Exv+oq/dcchbGP4gSfnIILajeARYUPihQRy1sTHPmWz/1Js
eobEqI6VaAssVd1FFXxB8e2FbEfCyBFnM9WWiQpkW0U7hdbbWGhigLs+zfBjVLO8htPnBR/w+PFQ
jQTs2eaAsLiRa3tVtGh9vdsoPHCak8hXCP/YS5jfSrElnrkZvR03XgAs+ctvCD4JKNN/DX5aHAjL
DBqOcWG88zVa+vkRZARJ+lNym7a4rdPds+ASvP1mEwDaHzCv6/EDZ+uZGnlr3zjbGB75vc7mSHJI
x1Bwst0Qq36adz0OGYe9Fmx6WfuE9UTJvJ0SaWxBGLryyEz54iYTyAt/ox8OSM9x5XFyfrDZmEHY
6LoNdJJs1g0gdFGAjKZP+j9/Q/q65JmWzBqdCZydRXUTqR2DnYZKJsvkKPw5jYpvikDVZseJg3qY
mvlu0sJfGOwyfDmjTT8PCjqE2nkDqe+QtPmzV9SuGXsR/SEPOxpP0U1dvFy7XWeRPCEoBKXm7GRF
ppnZl/9Xv9LVnKIDxZCbcGzH26f13DIyG1W/oAlx/Tvk4XN3B+2TQVHaHxYmzi57RJNJsoqHK1Gw
uCanwAwFtlErYYzAA8/x30/8ejDsDypknJwAjWGF8iybO/LEwa0qzmNP7k4z5pVhA6rwJT1O9RVq
tytVPBnTIPMNssjTfq6qkFHdvRHddW0VNDIdgOybRqRNCjJafMfv81uBvP04usYaIfiSztXa/d/U
uPHmpE+SW5EoOY56OcD4InYLV4/xJ5Gz4WcqlTSkxbuWVtvdNBSScH9DmHXcbNK+UlTnES0cVSRm
+a+ldrRcP2/AtzLH7T252iuzj1S12nYcxhiMI+LYNppRBoNrFe7DJUy9bc3xFRPW86my7OomMwir
Cf0HkMbPadzx4X/D5GhhSWaPbeVNYcQ1RmJjhjANpX9K4G597U5J6Xq9vyvN91P84pXMyfXwbJEY
p/KIzJ1FQ5+3gzIv+A/Ct1WBC6DRlhmb6jnKPByoQHWHaQ2FDhze8vr4AmJB6uQOspkRRI4odVXf
NOmg4pPJSfow4FtGH8+0TI88JmEMOVkLaWeCTycoGGK/QG7iM2f77LKOA3Icu5+748zk4Ksq+esM
TuWQwU7XT0GZJTTRpLOvqugPrzgvfN5OZE4B1wXwjWmEnrqLiACyLEb6AsZ0rmcHukk0guNQtXqa
bKJPHpm8f2ikVJssdulTp/IY1NqxVmwqlqzU9A3o9DrhUKorVENQbzyV0EBX/gKK1bk8n0Spe8YR
OhTb3V+DFSs3OMznvrB9F6wMfXWbysNM3j3qWVEchfqbzl40gtV2FniUcCCgSv7sZM7uKAbYlA07
AhMX0m/gyDPnXUHXTsuIjXHeVrwEvnK2M6DvQoYtsTOrQqGuL6GgHefeKAw0NcQy/3BPLPVOSXT9
qVkDOZAJlfadjOESxc1JaDFlFA4eoQPQ3WzGeRoozX0Tg7HmcXf8cKnX5zgka2/mE/6qCzC+MnWF
IiThpt/hhn9OUghZjhu2uf/LuMw9XcjyQBm5IZ/49RMZQfJyHDkesfXwxGVK1NZr67viGsWXcDUO
1LyKmA1R8LUM17I2cka9x3UZLCKxSmDtnXgw3vGI5992f2aNCsfXRuxCV7KZ+E5LtQkXatzQIkrP
2T0quScG/vsGgVz3PjyakJ8rFFclbV9p8xRuCZLf5yl7MmsjtFHn8TBp+CV0BWJG8sPUYvYSvW9Z
wTs8njznXiqXqeBNcVVgI9fL8K1K/n3oMr0HSD2LRlSncK7hLzTGytNoX2xk/7Xy5l0heFcllcaN
99ycjBEhMa3QCYBKN71n+OGgmWGJHT32Fw0VArI1zkPIzxVfbGzM4b7F0MmWUo9Wv+Ed1UciI01O
SVIRF9AMaytV4ef6G0u0jVdCR5TBQ8BC7wAuGeF6npE1vA+9FpzphZ8qMWFSHkCUKnZNYUtwjWXI
Og98CtqcyRh8YiZJoGo+8UrWYw1KdI+VAaSTQTbkjncCwg+ck7y1jfTsA13IrORlDbYLjFaZMGa9
P0mvRFlvMLxW8dCN8Fwhq8fJDuUlp29BpossKOfedLrEGcPiQbK6KML3iiee9v2goDpRal6B61xF
F/9/8+R4RdRo5BmY+uprUcaYrmD+Oc0BfI88+clZJBtB7HaQ60eA+qtwfQBjzxUASWCoCGrSWZzJ
h9TH9AZngORsZVoMYlFRlqNtSs5tfT0ZQjX3c9CFpPJW7v0Oy/7ivqL/3fzfhcRsXrZtbkjxA4VY
HsN9L4vOKcf5k7c/FHBRVu5RGn5R7oSUmAkzwESZKkiNGmyZnT6ozrXNzqCX5lRCrJs7ga6mjFBY
SEeXoarhm4oEdSnjYsf/oOGkTn1eZalUM/+gGl6PpshylSOk3r5nrl5WsSqWKXB6OcgTufLEu3KW
cg3zOkPX2wtdrX/Es+pIu/4Xn8Jbc/LqGo1P3nUZ4j5Aoyar7QQcmfOcK44yCgF7nFK9nzIhFFrV
JIPr1Rxm8zR/5MOMHuNLiGUD65nfpewtNXM1CbH8NPCYLS3Gze9KGhpw9Iee7yzXkct5/n/4a8f+
dsKMmNsoAIJjEJgizRNQguvvNBsfmXEqv65C9iOVYbZMDk91KEc6mODOCry7pMeNoJiH8Rs/a5jY
813W+oiwO4Iw72cNDNgMfmc3NTFFNu1q0nfY+1gVxPMWNsNyEj8ctkOkcWNyAQZOjomcOg9Manec
vazk6+5TgutOcC4DCnLX8eDIUijX8HUc0GHAkBII5N0tURsU+U/QvaNXRT8NrONPE3NNAZiWZBnA
lnBRWy5d6KVZpbEpHLO9yJNivW/SenJDR//GiKvt1mcH/UYhF97vOTsygj0Dq4CPzhVm/Oaqa6+H
pFfebiHX99yWyByqlBgcyYIZsyFl03xaUA5i86oI1KpWOcL1EW0KP74frf05skHHjle8sORp93mf
c/PTnuHHCqz0lRP0BCYs6YYxbzJUMFD+uXIDPi1XJeqSMGXWUhXVu7NOVYKBCn2Yk5AUjGjCE9uT
0m1G+4V/YwLPD/CcmdXR271QyAKcHdj2Oe85mD6XHM0ZPzhoV2S0Ipp1vPm92KKh2VJZSiFZ/6bA
vplQp0Lx+iRsrBIv87BqFIPWgmMku5MwjrUk/u5LX82IN1ENQu65w2imldhN8nl3ooibvrAIoGGk
deEc+S87vJZW3uygxERHpnJvorgE0YBPp2HmZlxMBt5w7emHH58BvYGtHnjtHGaELwUJGmprsAt4
nRZ88GwPptQ8Mb6iSnWxlAsabJlLdlFGNqDaoYpLkPesokylIAdDF4IH6cgeiD5nC48WSNO9vCie
kJqoWNWwhj0Q4EkZ6BNgzj6L0H26to+AQVWUjR5mKB1rdot/mYqzlEqKyLVY9KHTdbrnsZG74YgM
qLqey5utFZr9wI7euyXLOe97vI7nogBghQQqRXaM4AmddDN7Kgbi4bY2nxDgXODSWSYn3kb+xDJ7
nuMz1motOn346zeQzIcUe7xLApRqj/mjbLUYPKzjTnc3Dr095DF7EKaA/6kFizVPm7Spspo/JzJw
NI0Ua8ApyLguauzVP28a8CmLVqMuKsNh/LEqvncCv/tF9VJFiLGCiOhuwfe9rFMz/taSrZEdik68
KbFTo1fr3OLkW14y5i4roiEtFqRcdGXRIzpQPXh9p0FpghZ+qQ4MypcdCFawRkF2JUlUBqyq60jx
soAJclbuBYJXmGByKhLOyZ5dl6qXBKsW8LqTtE1Upf0+2EB5ICzwhk/4mtVUnb36JXmuYDvkXXg5
GwFN+FENcBuJhgr8TpfI+98pwdQcN1QEEdalWMNl3IgINhp7tG9BRt7GEZgjbKReDayCiZClTGgv
vbQrwopfoOcWOuYR80TmpRx2btUP39bcPlM/FOkeA1SqTgfpR6N+jepzW3zIHywkgZZ/8PMxM5aU
NZwRHRCZaVdZnE626S1ZrWMhNm6WiISpi5+/3biN+3yqhnDFY4hGNMRhkIAspW9uAjU3xV6KUwC0
NfERYw3B5HgL4/0/+ofl/xANyFv7utWjslkbtSZi6DFUqR9YXJB1NF7b9+H2NyuKcBGzmIE3P3jo
Hnbtp0PqDtclNhz6rtJP0tv4OGNsWZ+ZBvGLAvnDZ8M5wCAbCZ0uxRMbaO+yk/+Fpu2PrnpWBVDX
xJfD0NHcFF0Cc6J+t9x8jsNIcyYwW9sjbDcWmMAzQv9H+gXyVASMu6GF1B3TcEWPFk03CLQ0rvDP
8HS0UOZV7Q4+3yNY5m2PDnGevBF1OCrkqhBnJY1YACO3mTEdTrnfS1LvJip3nllALZFfH8QmAhpz
4oT8x6mHW4dnHrLs2Sr+OuVt78l/8Y3PaqFBTOZif/+KXLcTKE5HvF7wzKBkM1wnQhSnrqmOldv3
MzbjooPsQ47Jb3UPlchQPtb0qOeuvoCcEow0rvk50a9lBmDD9u4zMnbu7USqyV5TbTLjD7Ye++sq
OZXRmKbIstjRy2c+QCFsnJvCycmO+UHhnlC2QDXVQnDniKouUac/B73vRqhM01GAlZhfASIJwwVB
YpymqUyAooz3IYDeaJOwoMQx+r41i6FqjNAsDzUSUJqojqrtgBmS5HGMpjB6o7C4QHcrwB7Od29I
9YlDkUQitWT2mk0KAMDTPvyFRsRnhs/hB4OFW2/xzrJZtg4UqAAgbtRBCb4Fsp/dsefyTv1pGA2j
/dwXYqTDWmVqKnoT7s59yX3TchuM0GkGheZvQg1IJY9n8Zdjth7htHfxeiuFSq1CuX51l+g0u0DC
0Y1m56gNN3iygAVjX8TJy9ZbHbOPPkLW5wnWAtCkPlFY0hVlRdMRLF2B2G3PJ3rSvovXIWt1oDSV
+OHoaoQJlyE5QMRKAEPQdT8jXLbwqj2JeaeMwCKxr9AEbr0N5PRooPhI8vsl3SVoY+MsNSFJMOYc
Fw38rLldsSw9yKBlgYir2/Wz4jCC0cL0UlbtN8rnyAEMi0lVUYPSMf5Z3gbKhAU4L5+BsELbmoz8
19bd9S6EdX/pYoG0IPP7hme260CB97HBhLGU0McYwtHvAi3iBsIOkdgTkoNOZ5anHrG1cWQd1kaN
m5XAx1DVMa3bblFaU8ak/jNML+35/tEQTZiXQHLiIaDNFONe0a7NfrKq6PahzmE76Yv9HmLMycHy
VPzz+4TQnpLWGK432lUJ1wpKBq38H+Qo43qVqCMqtua1cj1XuzU+r0uBKl7hX/Q8B8BSF1as/fXq
VBeaxXyA5XGSxUi0Cp6dYUDVPktDOZWY5Mb9AagcWvooEvFhw0Fhu8YQugAX2UvQ5Saz3WAd1qXn
40yu/Gb/o4Fz7DvqZRnvNBRlm7XS7Gxrt6QgI4APTu4mC5LajyRKUS9dcYs0QkRgR+sbnjw+ZYCv
U3dFdXr3NoMhSAezNBjmIhmjerGDIE3v7UzSdrmr+0O+uJzAbdTbvZ/BtvObXABxGs7kofRQShW2
zRX6hCHBPbWpme6Niby1baJmM+auMuM8Y7lxaOVTrQJUenUAR9CXFayfM/evAf4E3+m6eJSsqOQR
oHHhhE3lLArXmV6vFxlMdrsx0MS8RI3W3uv+BYG2hsaWJzqyL8vJjMPUbqHAJCHu4h61KCzFFEL1
ocZAwCSaJCXal5kFyGW9gjF/9W8s/Y0rUgGWeX8XCczHuz8ugyZHZ3VWBQeY6tj85rIcpV4DIyQe
McbM8tKYUqAe+sVSuGAmQFPXzaWEPR5JDlXXJIq+IJpTei61t9ZVgXWhDuWjPWFgYZ4D0m71gXQP
CeGGT538x8QyXE759laipHFnh0vBMq7MAa5rZek/JnuL5aWzVujhOsY8XWbr0ifD/jC78G8y+LTu
5xljIuJ3Qk02KTiNDUXiR8mfmGOYKiD8alNU0IeHOf/7NGo/nqGvk4klfVS0G2AjW1HqUWtXQ3SJ
6muqMMzKHu98qL+qSVhnOYIAODNQnecTar1Wxb3JQErDlh0wH40LPbEV8XXGuoB0ouRvWqMbpPJq
R0wmusYzF+kVA53pJfhBiPOIzdL3ZOfRwHGkDpc2zA5ZeYSChgGz8KyhQasFk1vWpyW0K3hGCt3v
JPaioPwWvGkBp5vvp3V3e9nJmMRx0lTyCEQ4mQD8O2DYUFzwS83ReGEhzSx86s+k1IMrwn0cKNoI
PfSsoBOWxNRZ7QccaS5iux5xo1k4LEbqcWJG9Hgwnqfo/1+GfiE4lL/Pd5vJ53OWCF20Izq9KQVH
rlJBCp1Z1P6BigpeyiU6MmUndrtje9jAD7lLeO0QPkIji3RvrGC5QzAqu0dbAE4JeBMPa2k4HfvS
n1GUfoF19Hz+14neCKAIPOxUJ1RwmNNPxJ8nlOq+txLw+6njnYihnYtZRDhvrjvOo/x4U/o8gNmv
zFYoaTVA9C7go90XeM4CzuMQCRABq80HIqTP89hEQrxCnzQTFrvIg++cEgB+hqjcUCfsIaB1BSBE
MK+o/VStY/+Hx+EsTLtcY23mXQ+mUuxNEfZ1Kkr9qA+46xYlin82p9MRiXcwLxG6IfRVl1SIHElG
zMGlDPLHQtcqnOjyMjeX1gCDOJYRurhjDFK5MLGx11MJQ/ErdFvtf3Ab+uvD4L34lFzwRmp5tLXC
WpvijfL5MeUWLCUkBis4wD9Ys9g0TcKFa+F0nDb44dIDz6EQI9lM2wovsNyJdqOCoTU3uKn9HXRV
6CuldfDKiJxeSlCDavnLeu1D1QFhWsakt2nYGeTnz4fWjNCEV0YTc+CMM0DK5LQ7hBb830UBHQR0
eCC5rbHQ14CYVVBw5qCqP4WLiM7HbZYlFo2juv7jzl8dQktxfJvZCbpH7h2CS50Gm8LPqP38O/Pg
dso/RIW5ZXzM6KL1IsT4WoFUq20I1MHhgm87Egpt4FQCURt9eMDLEMwinBIjI8KCdnhXT1K9s8rb
1Ic394+1PLb0tc7zoydLz7R5WVqqeQRpVERDI34nKfMKPHHQSzuyBlnofbm2OY27h7IOoe2/j3xP
6iWCkLqbgSrAm2IQ17nQ62vbyayuNBQmZOsA/Q24v/EsdGpKYzHGKay25NSif6EpLeS6b53kZwQX
eeFRlgdwvNqlXGQBZ4HESkyds4KKgZio7kcPrLrxoesBnDBps0mQRiSIVDf6m6hAZvUdM8CuAehn
tLA1OpTx0kPOXRTdkpIJkaD+K2v8ja701VVNEgq1EwjvfGf8xdw/EDF1UkJ75/XyZPjh5tyUH1an
554qhxkyN6zsak7UJx9U/Rq4T18vMQQVY7x4x+PCOJD3b86x4HaTONsjQRtWLIqP75R11CQ+BaNT
EKm7d1OcN/1XsDyltsfRUyE6Hw538l22HERURDQkTX3Kno9QEz8htIu2xYNmopcESDnBcPIGZd3d
lLbe0rVEB3kWtbBhZKpyKlnBBGhsjblqYSAf4DyfyyvED+B1uQidb6dMUqsxiBKk9ksxTKgaALZp
GhjU8mIdmh27D29e+yrKgT6f10RGUbvgGjGrZN+YMEI2U8JK6WacHqS+tYxI5ThIVwsfFH5Tp4DQ
SXTXM6XK6keUGQBmNYV/K4E6/H8Fi5kDvnnL8TvgBoYYKuOBkTNkICZVBuEWxJXsm0EvtmnhhO7p
QW+pfxlTwdrvm40Ro/vsISm93aKzvDCjykzM/MuGQ5xXCWH8VhtDsz4oyYc+Vpmbn2YWUao8AVVT
DM3mqJyAToleKofVydsclHjeaNAVR3GL6syMgJl0wwF7PShZ+cm42WhDkabfIVKQGvUOhUx8s/P4
xZxHRkn6B+TP1WWatELa88jSQy/+3F9mP/zk75cKB/Wy7qunGWIlwWSCvQhRM6Pt1cv1sz8fSwI2
tWCz4Kq5WXCPPN9fhuQshdh4pLMMSQdWWRD95u/4FiTmmq+yhaOOQRqBt9omKTuacFJbjwuXRTvZ
VnQY17/ejIL+xfzyCoq74gcDiznqtJeliAvgcn+w6oKp08kipqEx8ns2NH3Y1xRznTmeiyKaRyac
8DVjArH8fdTW7/e4I5W85I7pTdIiMjsguEmgu+EZ0DhFL7zap9uG4g3h7w8ejtuZCZH12jfI5R+t
lVpS4SIRHDEjzYX15b8NeUu0NyVbBo1zu1m8yVHL2LpSAdd6xxYKOnMIdVXW5q3Pw+vxg7bnqduB
ppVhwC+GdgiiWS45Lx6d7Hi2ZE5iL8gUJZTJLWks/zLzd/XqXTiIIekc4+VWrlvp+SzqNMjx9zgV
ii0vWYglj9F/sb8PQUyU3tvOG9RpTX/4ac6MnL2eNGUVHvmy/+ABmcKucwGjTvy4eStgSGmxC6g8
sl93Rfmpa9v0zng4VQBqTFVR+in8MgqPmDO+iY9z5Z/dOeWCMDKr2sD0Wa6OjCNkR2pHZufrDeqk
q+HPPWlGAfAVnC9jTSyi98egBGdCuEJUm9aIDt6UuERsuQaIZPmyIYcCeXkJo1WNE5EfOZPvXVLQ
qZDR7OKeEwW9czq9LB+XXbseB7cwLmsyV6GZJHY3Ufs/6BJkszHVCx72zUAfZclxqUQSNqbtTnNP
pl4HyOs6zyd6i7OE2Vdns1S/CYw9QqRwHf/+XJR+7/Q5vZhABL85r4toymQ1SRIkxql2qm5HyB5H
Sdns4H4SVJGv4h9ew5W12XNp2PJj5bhuxlCRH33ic7EgJ61fIClf+sKYizLCRYp5qnrG/UwhZBF0
RL/w9UPkFG1d0mGpYZaFGJBCisqYHQZDJZqZ92SI6WPnWZeNutXqjqK6RTT5AB6k9df3QBKUNWSX
YCGXk+leFxynNBGrejK+YouFJetadp8SrO3xFmpyYu4RLRkM+cNOvvynSTGqF5PYiT1oe2igTvgP
vpMKeTTkB40BzNd5EZCbVJ+nsS0GPQxW7V6mvZnK2VUWEb0SGDkN7VrtL2iMHv8bjJRuAGwTs71A
1YOhq6Yowru7oFVxBlVQP9JsTVKD4az41XjLZlZfI8TnaIR5GgwZCKmTgdwjO/LN4EZIpEDHSi96
MSbwlXlmYQ1R+9wy4aa1DqTnz8kQyq+JuvTm4z175tmABFV/lzJ6WNmLl9AVAk+EDqrTvr7dQJ6y
CfRGx4Tr1OhykdRyWtYqjPPktLh0gr0yR6EZn5/R6lhpyZ/BfmwwgKkVPIe2KtFdGh2pvPk/XS22
Sz0SGnahXDQNNtEbiNghkkHobwC3lWKMvLQB1lnctdRQtLDpAvA1gsWm5IxYnXkS+we2LWJaNYhW
DPHqZ1a1+Y4+B+uzKkvv2C55O8NjaahC7HLw44KPvbWROqBRSwmx906uSjDwiIdMidgiYv+k9GTM
ecx9PR6jv0FxIQntV5Ld/hWAKdydPaPmr5gZtn6ICOTvllpfVXLvVfqfqznTEwqBCxtYgCwlPwah
jTepZm4DtRMywKklO9Hsd9cISbv/7IKCNnHWrXS22SJZuDfyn1WKghwQwMyKXUIKQ+0mLA2JGOVB
NDTy6Yxn5jAq+ThGoBOQ0rsRUUvcTN32ZuNzdq6+nTpawgBYSBA+FSfeOmnBlAN/Fe81QweSswVl
lB5EEv+2XznQE6XFdwiquP96MD0Z6s8iv8tgJBL4bXNisy+Ir6CSjjaX/344RW1TzAQk47WloaSf
Y1cC6XtN4KXydOtU/7iB0tLiW8a1R2urpZa/0csok6NIC0keJ0XtPGHwi9ZW1NkDljQ/RSUFAKKJ
hAqAty+JmJWk6ykVMmdowfyQPJ9eCsJxniPODYYZquxH7uEsT8b5s0qsqed3Lh2X0LA67LJxGpWF
U6LiwFiYHbqAltY2hmXsDBN18rKwOAlHUVPeV1HJ7S/scW4kK9Kt+NrmoMWc5P2bOdO/YFtI7R84
tCsE0CAi6n80mVwfx65UFuCjd/cs1NTVNdbDZfyPXa2SgtDHNcDPfbwrGTeeXwwADTLvfoj7JgtN
mBzHTWSaSfvbvKR1WnbJrfk++PD/LPlyMFtep07i5kjwgh0Qrzx6Oz80MCIR1CvDiju7eyH0h9Mq
70T8pLR7srbOHV1TcTvcvr4kn8Y4t6+3F403HC+HlAovcYHqgfvyHg7K1BF/fKMSTgKrL+37xlnO
cowQwLan24zV1wAt9/2GzkCYqBzEofG6glKMsNqUIlOiH8v2ehrL7PSYlsfhBeglA90F53bGiCst
tdVbENHXe0u8zefn6BJZix0+6anokg2gqByXdcympnL8IHWn3UeK3Fc6Q1SiV7Z2C3SzocNFhyw4
3cz2tJgAI2yT0KQkehx215qUG+lVHkbi6w4wlYnknnne9A/iH7dM08jb4hxwqqqvcD/JHad+TJAT
tnGzO/PnuNVvYLVQJ18RZcwW98e2AIVgjy4zMSGYhneSvvwpTUaorZN3hi0+umI4kHZDulFLPNo6
oN0I0ei5tLqoBCslYzxilIcf5ZhFlOJ0Wrrgd5Ro+k/NkByHHn4FM0CDm/qH4dYDFD5AVxRM0eIJ
tUSnTk0zfVtHSSIQaHwk7Ea/ukGvkrlbtAUsaeJpfiOHULvVvB1TV1/EvKlTi+sDSLGvqNx0THZ3
NuaEhTZf1kTv1QVlzIOf/adoqiVg9/uAczzzJc6v+x5msUGFe0eoGgDho90OnwTRgoQXOfOzPsvN
8E6CkN9Ac4UW14GANdJKIl8T7U2IkC9BS4bqnr078IWzZrfazFrC9EtvR+G/ENIaxcjrxDQAg2bH
7IrFSmy8VM9IB7Istsl5UwaFZi2ZlnH9ri5lTquP+kO8Hm+QAUgRmeryU74wDw+dviFMTlsib1q9
HC/6y9Md0EmyJtyakhAtQZD6DdLn40Ob3bRFOA/uQST4Iqk1ctPgdLJhS4islXdVZsskrCvJ7GTb
97LH1FDBT7ZWgFsN/UWlfoKkGhKY/zfJph1RGnwyLnqjynytUbHmY7sSFnoJirJonFtexpWHdsUb
pifavwofNxlRq2Tl7V40MSIP803IhZuK91aK5ERDFboa3XETbYrDp9V5GGUtBi//2Cyg76ErK3de
rpqKt07qOfrTA+bmESegHI4ACgf9rk8rkC5Pz4BeQOYwTa6NXrppmzjz7sOBPChWp+fZNfQPpcY5
2U03fd3Mxn+IMXZmhfff5f5nfjRWfldNKE2BfidoH77j9XinQlsDcex9Zo5x1orN7jKD8dBNJ+Dz
kdtopvIhtuO/3yxu+2kKEyCxbUSwJsqkVVX1M+/T6x+6yWBA0jdWVXzGWMbkWrTghA4GlSbm4XUA
B6ibLB1jwwBhiBGrx1ixEcfpBBRhT83nIqiT/7nNkXSKxlQQUwJFx+f3Cpgqbwq0G7NRm5HGH+jI
GcKCy13k/gsXMatbICEPT9oQYNYgm4e4+RmeAnm+sKPucMs+cHYJDJXon3EZ038hTzwzdFV5bkrt
2ZLezhLTbqjqV3n8HoqyQmPbrMI281/fvOozKRYU990qkYkLGDvkmQCIMF+Y9N2grl3pt2WJXA/e
wZ/ZHO6DZi0hb0cSwSeaQNl1gRIhOdGWcq0/T62uoXV+V+VVcNwS7Z8JVJOmarBI59vwMJ34FEg7
4uGY6Uu2Ug7mlnEe+m/WEw4SLumhfi2kUjZDmmBnR3DZtaJukxuw5ccHRu2CUw1NTGN0Nl6gPdLG
xaNXi0YDdtvJdPlzo30SgUJxXJhpL5JDXMPShBGAILyF7p2EHa38j7zGjUczjIywrTweTTt590Ml
+vU/iHHy8Ef4BN4v/0D04ckq1vf9GdYdTvYST6XPbx27EoTw9LnmN5aj2dbSpVfs//23ZOOUQJNF
URZ9sybZZ7tPo8Pkt75FL2yEX01jYb5XCFrOIovidaDFx+S+X2D8ZSk26okdnfLUfJflcDLnl9zY
hF3LwtmBP2NBX5ffeK7/XrwWQX8f56pk+4k5BvYOzY2ZaUOZIr6IhXyDtTim+e7FiAFezzMRptCn
Vp3PjsJBDu0lgsqXwdb57DcV0knOQ14JkNBUVqKSTGEjCJukbiEaVsjfyK9o30IO/h5CLEH9JfWe
sSHvTjCXsDrHZzOVanpDUt86TLFkY54EBHIE+R14NR2vvDIHtkrcrpEJUBONjxzyT8kPcXGapp/Z
+setpU8PtL/48lg6gRw6iCU6Eu+ht2D5w0kDr1DcnjbWPMIOWTImQIQVhk53RUe2xiyt08XtZXqk
eBBEeWzK8+SL22VRg7pmyV8Ia4Q6mKbpfsjfbL9eVo8w6+hbeivLLYEd8t5pxIefq5ArxzY2T/mk
Sb47ZNtgmeqzIyc8PRAuwPEpRGIE2RGaz0xn6Ps4d1xL1Cd23qIoxTEJ0UPiGefOI4trb6W65np/
cGVlFJ7P2FnCtYLtDj9XzTVqtEeBgBeFq4/lPtD9NbltydEhYVqZWMQU3m7bvbQTfmOe+EQWIP8O
sDjq55gCnKKwXIqOMZpiZDdcaI/ul/SE1XdlKhPspPEcUb09IDVOWWkHM8UkKANQuOTUBOUq0onL
cA/kAd8y7Yhr/RmDxVcq3/zZH4Wnp6jq1+kecEbUAaBGqVsT3SqTU9XXYQ/pzZAwIQbBuL/NDitc
WWkejr7tK5TvPJNHYWzwZm4E7Lr4Ieao1WQ7HxAdprTz0+btqi5ct1rZSJgU1rjbrG7X3VxeDtyL
cTBkbZUszt95py+gI9+n1ODyk1qib+oRE868DpRwm9qoDbwdXAAXGzXmPvyyETebUx2rLjyA5iEU
FK4f6Yx2fF+XpurI4dmYbCZdK2JSM57nwmB89GBc4RDQL/exCar2DrFerkEcG1k0yskLCVh6DAab
d3q4ajo+vLk79Ku63zy5+o3Y3iDiiX1enUWjneJOm2YZWhOcKp0OLyZ6T8CSuxoXJYMuQ8JV2tzY
KgvGDy3u7yHuDyI1Q/JZuDJ4aaB1EARDVaRpIPIrvjhZ1elFm7niOac1RgMDSsOXkEBOuE0nBFHd
xyir/DtdDkwvg/mhqp4qn/daOWDmTtfR4ZLbF2m/cP68ryVeAFPqtHKiGVmJFMCbHilOkT5FpqgG
PpRMBSrTJNQrflhrFH1l2jiCwiE2MzYlvdosLb3YfTjpAhubvmCms8iSvY9VcwtFWMoUPof87Eh5
6i0hxzJIe7GjIdoSOmkFS2WkPRG7kJbKaTMXSTRMAT5vLv1BwKIY2o51wdgIBWBhOn+DnukWlrtl
3R9r2yd3DMU5Hr+ct9k1juADhyuc/EN36fDPEApOc3jQ0f1GJAN7STVBAqurwrfYPg8dK2pXVOvk
QP3UFYg/gPHtX3hXsTrFSto30kUAYtOY/scdPoJl6vLzaO0kor2fykJIdHlbIpuni97ZxSyAnbqe
qMYFlK1gHgr+AIcWNQcZqvDRug4ik/JAWJMRStqv2lZ+GWD5yTccVzQEAQZDDkoSSE7pYlIUQF2Z
rXtIEr2loOqgDcJt1IrI5RrWFn5fZrghjmAszAW9Adi2mTlkHH+Z9ZFOWy/Lt9tn0qeM8Wjrlzsb
PJlUnWZfxxHE2e7tnfaEEpUCE3HzvDxfKAVgtQPxJkNi7LpoXXWMNSiefQoJIoOhgoizzm+IPhhN
Im0jcZEhIyMBRIfdT5i+TbgPtJvDeg7lILRo4kygefiwoAZIdxOVp/rQQxxseIDQIAZiTG6P0oOz
i791PaMRgEEjmOeJWvKz+sxWca+yCr8OxawKx2yuSVvcF2jH0eojauTwHfMuQfaeIeg2H/LueXS3
mENnSRuoOqXbMSAoo4pj1/qYkm0aL0/qLPJikrb02hiAxC2OGO9QL8vNH9SMBT9fDdj8y9WXWPXp
kNPWgbu5hmvjs4XE3qIK2TDXIXHe3ffrHnfVuWUvDkkRAuyTUJikh7BWOwcgBkyFdKYrMdMDov9w
TfdX8dEDiOVPywxI3ZKqpgUk8NO3Q+kLIRk0+aRYxOAJ9LyrLbWYfk7345WvK1RxXwblSL8vpkYA
e/u0EBj7esxbIemgJ1Mnp6VEDjGDrOmLVOqgRWjzNp/KFR8dzWKrO7SpizGJPMdOLAkdWmvRBZXB
8IQy4laprvVWuvP9Sua7CltwaXgRx8UHpV1CjvZxba8tGuY8JW7pBFYRHGmbMcW8L6f/sHNQY988
O9eEeqLd5fhp8Njp96fgFqokSHP4TUrzl9CK7Rvj0hSdUl4JFa8XEcoqYBdmDDsqlRA0PVN6UYpi
WSUeJ1C45sm7bWiaOFRnWvcMT3bDDEkjqEYv+1TSTIO2cqi8oqFKn1z2d3PbNCI/S2bMgVOxh906
Hygh0wKMlQPIxxi9R/fJ86ZkAO4Oz2DcJU7daEQ3Il1566RgYugN9IxO37C8PIDDxHQZw/ZxFd3F
0mAWfX0pMKTyI9cwdMaQcN8f1tlf5WsQlA2ZYPC3JKDE46LA45a9iW3hdYxVFhyG2C2xuDLv1ws6
NzJIb6boBpWih4cLJVt48YZbSEck/Jzyo1ZFxsiSnKr6pjdBvCHW1OrCWt77SxNYl1BPvHePA2nX
gHgVzRbd8FCt96FhdkkJlHiFgPiBPsfk5ZmjPIN+jg+2UahYQoJD/f6adQOh+GpU3C9Ez7eCWEmy
TvJ4IxWNdu31gKD7uE9hJvkl+fv7Gz7T2wTGMfacU2D9PuTqCoIoE+MtJtcvh1TdRbqp/TL1Utji
v6FtpHa0KKvMpUwa4C/fJzh8GD0ggQv3hQGD5a5yTs6ewZjwc/OfGsqcU5vJQfGU8Iiv0WU2pd8D
maR1XmQaFLChXvu+Z6iN095mqlPAHnfGJNbDVpmR9YNUvimPxOTUuEFEpExxWIQ/t+5wjTN+WlB/
93Z4Aptdtj7H2cIsB2FDSlcyPxw6gi0hURg0pwl2xieEKS3ntEwRpOm0gyu5NhA8kBydVSYIU88v
ULmRvfBTSRxHvJ1wBlVGFJefLmGrbTxGV8UGLmsatXqYSkdSL2/4hm506Jleub398gO7JHp29Rt5
r38StGwqwcm6vyjqf9JZ29SxX0sE3U/NVsoD4xUqujKiDW0PRU8d4lXZtBEoIzCtdF+y6qE7zMiy
kvDFSnyt0+6DOYBELbSqO2JVqjFW1kYX12+aNmfxEFsX3L/47bi91u573ya9dFynCHXxdGequ0qb
/0RV1dng4LCyAhlYkF4118q9z9PKDXDyf/BlGxkJEaA7Xjll82gMOMqeVNiIsrngMscLuafSsguE
GlLULwmeL1xB1TaiG/wIeAPaMuiScnn6zBssMTsW3H1zysVQS/pcWEbK0UcgFbPAqaBAK699m6WR
NZl1IBWE9l8p1qSrO5GSqvHbXPPnhr6DM519cutC2PGQ55IszF9KiAELZZpWibVWoqbP7ww0Om+h
alSdXSUhGEHraBSTp2bUxC6H+nvZXC9TRNbEJr1sqfrUanfwP2dEFPULxbbxxNBhGi+otqiegiO9
9f3gfQCzBuVlJ+lx6lS/f6njfYbAZP5x9oUeqHem/LNB3PoGJtmv8Q6s90iTQZWysSlFZPjxasZo
nfEiv0HKJm9m7pRsd7likVnTpAp82J2EF9CyKsFA59qbQZblr+0Uvy0iUvXD8DBzyWWOtNwVYVr3
BLm19jHDnUH8VihRKRIDhMhLC4qsJPovgHyE9f6X7/euzXqnV0dZ+AiEbjhYnCGljJRPtxKQmF+o
58RWYaexAqCJfPx0xC7HsEcqgXFA2/30+7j4GhU9ddvbJIMbG95Kn1HDTvyV86rBuId2GUyhsbqv
QtETmcYsI70tHmXy8VLN+DZFB8CWZ50sgE3r+FwN/hFFr5y1n+rCHtnRF2NDbGa57E4/yTIP4PCP
VgOi6P4AD15CR3K0bU1TMaycO/zmqu0pwfNfTpMz3qIlQzLHTvJ3EZHMGfbaVxY0Keku3sVhex7F
OtZiaKNY6/6FnLxdbm4y95rcTSgR0VENH7D1SOAjR3ufkl/zksajvY+eNp3INzSv3j0XrnES8Wuy
FOzbeDfpdjqpsNNmqYIXMylfMAO7B1OQLzZffVCTi72fJItw97UMvGQMke/csZInd2xvcl+5Inyn
j4IKwYgQKoECU+Vu9DD19gSe+WJ+MOZ1jIF2j2JAxktXy8ZccFsuWG4+CTp/ilL61lIdRuB+DNBI
ookGIbZ8hGoUhQwbTGDUFJaDj9Vswkp89x2KHko0VAyHkk1mI3WRjS75/HGg6b38w+zxzwwd1ggV
mt8bFKCn2YcU3UKzYbanT23gER2Tz0Q8vtDZ1A/WLAsqJ6LJJupd5zr2Z0nd7mZ4cy/SaAv67Bgj
QW7BcbQR8nLK3W1i3ggM/FGQMlmstOYa/L0Ta3AebaUJKPMYfN2WqlOIALJ58fsCXaIEHeXdRT7j
akQ1+DMUvJ23OuooxSjDWlWWFU6JJcg0f8lnYdNzXZjdXK+topuWJCCGxo9s7wemDxZo2iI8KPXO
c/XtIyrXTjW9O2CJJ3cuXpMAO+yEThbtHwtP9EGFsyrigkXuZYUnLzcyayMBEzHcAKV2+BHOpNwX
X72WygSGSN+gLRaSMTr8j1JxNKzHDphy4f7HGb9ukT5xWIwCKpS7kVhnw+fduzZa9kUPzkbWRtma
eAGybFAoBTzLvOJN47lld/TjIBwUMH7kpLTEBUqK/u4AjK3Q3sxJsnF5qgfECki95CBFsAVc88Mp
xYPXjw0IvFALjbYHhIALEkV4jz085/+FwhMMCfOQGSeZsvxXXRG7IzNWtnnzJker+37b02b++I7O
97LDaUwXG778uXoV6vPMGRc9gU6Fg62luds6Ma1DezbPOwPrIQUfBRrGWcXzWWm56bD/en+ThD8K
p47oih5gdqxDvk1L0kvDEdUEnNwdUSAUhp3KFxt/JTpb8QkFmL6Yt/ZMIIJIAfC4jvecMdMT15Rn
iZkbgnnyb+cibuMNQ9gdYCFt+9k5NERD5psgxYeDwg9JNtW/9bbOzi2c0Z/gUcOZst4kjfG0/dmT
K9BNgXn3Txvc15HiWALdvogTTTwcFyJXCpQ3MZQXzeY1s4X+4XNJ+W0ofVBZg1eN5WIu3qD93/Z9
4nV9XgEk/2FaOlM0Aff45GdL+8Ro/dk9IJsYgum54wfkn8ualWMPTHO0FpS5KjN8XKL7g+Hr63my
rJoFLrScbuSbLFxYemoz06V2HKaxg2Bh0flR1GCVm/CbT2OiD4g0txrS5zYuKcYwdfHx620tLLQN
874TyUregrKAi60NuPad2Yfq30DE7csoj8zI+FEvnCmk1W6G44XbNJoSVBwPSWbxZfFA6kUzbFwN
6HNfGXWaZl2aDQex+E7OyBnbw4GIzzkL4e5+ByCYGx43gnH38IrsGuwjHyk0a9dIlcsAZjXWWStQ
QMwO3AFJpU1SH/JBxh2+dScHSraMymMh6OiVELT7L7HTlsWxm/a6CtbDHcOGpgvhBE9XH7jzr18D
st4CYpzDgFmOIlYonIU/z9m/M/xfGAJRtHFYIy+g9BJHfOzOwb2WTTTNWdelpo4NPM1xDNIa39m0
Cj+v2JVizufPQVS9LDr2tWINN0Yb4pUnnsMQ9lvrnEAdcfICPjpiLPmZrDbGLvLLgoSlLcvL54e6
t+E5Qa5XYim9tn3sFQt6Bf4RKWK0VAvFCaRoQcfsaXX4kQcHmD6Z460x+B57nK7VOMrucgbNSZEe
h/8iDlV3LtjDOlcgfWdJaZJnad1IaImsMxcioLc1EevzKdd0pUWIEAR7tQ7zalxqSy/Lx5qbFV3z
tO/DrUBaedvI5JMR8AWnXRmSeSnx7wydPAKWWg1DqEL047sTNpa8A877dNlIBmb2MM6HkT4OWZiO
zUTVpWaTPKWF4jU7ypJjF38LCYH/JJWDnmXVR9lhv/vFnQIFQtUUm/4IgUPspfWI1P1ydYrax3ic
pyOLwcARV3QempYF+JRIyxlQn2ievBhgNzLXh/8c05VMzB89imsm6Ibx7NMdzyVzDoGP1XtvWeuK
ye7d6ccHufAb5dXHFk/2BgM+tChnm6aKA0TudCAGhNx/oBZqGvkLWq1CetWy96mA52C35MOu0NR/
i9ZCU+7CbcnEjNtG56yG88lqvr12kSKQvHUtPgWVD5E+cIkzN1VdE5T56YstRdjZp2QgDR8I2BPp
L8bWX6KXb0+fYwOv41ZuhxMVQmE8j/l5D537hDUt20AIFDws3IJjrEZGtehgeWomYZAMfOUvkq9c
IKcBxW1/yNrRkGjNn5tpZ4SXUBpOHCgFcW04+B9DaoXYdhRR64XpdbSEfA7GqUFzaK9Z9xc2n2ye
6+AE57IqWY4jznWWKh0fO12npl66hWqfvnE4jbghsskdWOhfZEqPs/du53wA0L66yBhl2d87KgQH
QjVqkYP/EEv24UZCW4y4XPfROKWAsTeFNx6CjOKvFo0udxRCZBZfm5ZEAleGeMI4D8cAooLU/qkF
G4ANIBmiUQ3BeEqBT3RQdJ5FDYPy/lGgfz8jaH2fLt95qu6ZNKwajbsvYH3HJ0GVwJ5EbzK60blB
07dMD0pzxv7aovI8Fx+toZC2gmCIciJfJVr3BoCkxaSnZNSu/wtfx8lJ9oLQf/yFGMpIkK++MDPS
g5ZKxEOY0f9+ozXbD62k4rnIWDpFqLUSsB1mmMZic304g4Ydy+LoLoWeHMtejATSjexwmWUJdrBQ
ADw+k5KpJQ3L8ooyyGIKEFMBiprd1WT09P6l9hnxaCtYEabb2v5qzdY44O02AtFyswOC9+phAScM
RwzpEUeFhcXJY9FHQQ8/ocjlZPDrNAuR3Flpt7pmerMa2dZr6mR4GBaKy/DBucn5Ime9P/e8ZSHD
HfNu73iKJReWVb+MVjn+LYFbL+HGE4YAVpXWYBzryDOKX8EPYHs9PQ1CzAVPcNVo1B6B94gaGyLo
K0cwKv4FVc5QiXr8zo8ZH/y6kpEkv5FIXYLDr09fnN3dP2Rbkb1/Ys6+k0YWcB7Ns6tGrgelDVHr
pgKec4u491Ph+6EY4rXmyCSVZFMLcRrC0HNYbERZMhikSgkNLeevghb0Bb1HOroRbESb+czt5oWk
o8DprfL4GN70bInNtS05fHtt1FcCqWXD+AWtLu2I7kZyeevy7DUG7U/fDOv71SMgwqVMpnivtohV
QWsM437I8+rmwS8+Yy08IFSLQRzzvsxc4WzO8jnKeNBHHr69LJc17qWwqLfoMv2Db5NrvmdaWf8D
/OqFzhZ61SxLpCXx1A4paaBfixXuoO0SnTC+NviDIb3uIiPgQb4ye/rxwWrYpTy/MQxoZW8Etce0
OLEINP2OjUwr0JE0jeRFoBe6dqPGsdn7OUVPJErlgI06getw59MMsh08wz1Sfy0/4N3lPbkBqHg/
QQmmbHyDCP+AecA0uM7cdhxh4KTW3pT7TSFNC4XT9LV7DgdcpbU1vqa/LHc9fmyCseVq5ZlOwdhz
2wooV5krnqdVAELPhDx5PwoIpXoszpUtkwJWvngjq+3YP7rsVdkvhAcyw+B0hdtNlZGQlELxnEQu
BLLPs5kYG/ptoKRL4qTLZQVYd0ws7b0cz2u3z5ttUmpLHDAPmLGl6qUGAoGUhe5j5g8Pae2WaL8z
cbWneW6by5VwVQwUXtwkQdYk4/5Q0jSPYJk/mDajMFN3T5fJz6MwAKjyI17TLni/TvNskrIpRPlz
NUS9lMh8qVr6ImXttoKtv/X9S1HvGegOkc0Kdu65CxnmRSAktVaPnBcX2xifzRft0BNDPxAlr60I
l4Vg0ct7IBGSZtSN1NLJ+SkC1FS3wsuzmGiIG2FdQoxvRebrzklC4qeE4q5d0lmPl6xpni2b3oQL
ShMgPGj7fuXcHkgX2yW6Gn+TurZtlEGOMTUiCbVqa/ijYNAzcBIHrT49rSsWXznj0FTple5cK6dA
lPcSWHpvhNmajgGM93+eDvGGzqjivAdfUx+LpNKi9t0SYoUiP0igeITcsh45FYg4b5MrkCfIwCrz
SIuWeXJD+Neg9NCPjEYm7Ig3OumNOdcdx3L1zkm5HoFBN8lM7GcsAzNWuRh2y6tX+oEbqMWAnhXD
pkq6yCvp6MOFWR/kGm3Bu1P/xPKZQdq/NXufmbKE6CBM6i+MVzIqfOfG1nGLMPLoRY+ihFpQVCaD
YAywy61+uCxRMDkx+zhJWHsnZ8a+Io4xq6pvbzubpzov1waipgwzG94yGKd6ht09hsk71P6/BDn5
wMEq07ADwwTEDWSXe81AprtU2HRrrjpjHxq1pUDpu1abRFL6RHYGoghz1oSrTUpaUY83/Ju4zUmx
6aMnC0qObRZJbxHPtFcb6T9I/dx9NSgwthfZANh0sxpFacn+aeffwuz1vznON4nkHOzg0yRKhm0p
2twFcB3tZV4IiG+moJwsns+HXwNDbPgyZdTA/rkirDxz/Ajsov0AUHsn83MMY2bB+UQ9l0pDfmn9
RXR0uW7owj36+Rd4U4t8hyXaR/+I7jd8tMuzqVqixfELEJHGfBgo4tCpPayxKSseNHOXuAj/nbMV
UpFFW56XNRgOLlnvlBTFjlSV+wC+kcHFOeFiriGvoS3dzRZ9kDkXRRMyHdj++FPnYvPEJAUn7B6v
Fuc4YwOqS6RckRfwk1n5+rlorq0asdEBqvzBv9qMPi+JFbE06y0iBPbwWq6Zlgr5D1YMZ8VUy03Q
i8hr+1GSA7FxlLSiVYY10cdO9KY4RatgVL5m9g+BojKS/CSlZtqhlET1mCIhIAsjKCDw7MDT7/1D
qE1I260pF0XeVgC4XKaIpJSzszCL4whQGI/iHLTVDuKOciZSyDW6DHsL7Qe9KrMaUjG5uvgMdqwR
Lth4Qd05IPaiVJE5pV/hmoiQ2lkYevchCINmNbiHz6D76g9kuwTsah7C8Wy91P6PXVRZb6/12Gj7
7FTGYX9C21SKaFrZvAcYJjxTIBMZ9ZRtgwLZwnObQWbEhEQRjDt2qfNPJuXO2bOvXmvHjZWmNBs+
B8SyH7WNgB+XcIudGs0R+pY5EqnVXtedghUNKKd/D0oV+rdGS4u9bpooAqUzqlWHC36l7IqGFdN5
S2PTA4nkxHl7OMSOFr/RWVxsS1DSbrNoo4xQuJH4K9o0qLTNybAJk3ooJtKoe7QuRAv9R9gBMYD0
x2oVxLuHFWHerC7QBqod9Db8oWUVEnh//nOa1dMHYBK3lbinz9XzZSplxDuPW4kEAsaSwQp++aFo
ceDdra25lIeQiNliTICc5Wz+p3XdGs+x4gBZpZnX8X1Kok56zLySy57Twbvush/eWPXZAaBs+kr3
g8K2T9+7xM9s+9DXLcpkoLcs60yBiBLJ2JvYzAYJXLYZqSguPZqTtnu5vVhAM1ocwxTpq+2TyA3m
Bn3Zgzj7SHjPSjg9LCe5pgZkOJojtklfUn+Bqhyk7jRE7xeqeR5sochLS8TUFW9ws/IF4Io4wDJG
xIzFp74a8WJQOOk8XiTv7ehGWB+AsmjkiFrmz/f5XPfFH13Jqrv2WQAESnKErV4b0F+HGXLRqA5Y
BHqK+mYhYPaGAAHYCBsdfnjouzKA+0T5LgQAMIN5Zw2F1eHrIdUkv+WKDCNOJvg7Rmg/xbkTK40M
496kCpmAYV/Sjrup0fZacxzdt9sk3Nm2AG72AWYGEF3DLSs/NCvBITdsWskdTo0SvBgVCcFALgWU
cawLw0FFGZ4rp+ntoAFZOHI+RychgUUouzOd3TmVA8pkNWqmL39fLTw5N8L6prTM6T3nrKxxk+d/
TMUK589aRQPR3KAoeF7WfAOeQtXIYNacVkNWiVZ2+kRfxIhUYzfb3Hri6obkRUnowAV/2WZLqe/R
POUNuhuSBs+8YdpY8QIT2zRRLAnr0E30VScifbXV9fg2kl7wygrBp1fgq5He90AmY+LRo7uOJ/Bm
YYhDeSWm8I042MUwG0LwacOIErqLemSBRl02b0kA2Yk8fHhXRRrs6DJg+MsE9Wx59dl8VfV3j8Gi
JKOpwcR/mruReTaRO++dMHF/WRa8nlxrj5+ftCX7LGWRekN0BxK7nZDHmmFpH2aqiTtxukmQQ2un
vcNLw2Bs4Hd0w7oWC3JRwhEsqb1qWUop2j20UaTzr93P8nnMGiNmi0lZcijQXm31Qq5YVz6BzZlk
eUfr1Gkahs4T3y4CxNjXKICJycKjwHWiLFuWRJyyNtUty1uYGVPfgwKx7c3tCOa7Vu6reYG8RWrU
UDuICgul6wa2vtAriClbS9z53fg6ETF0uoml78Py41O4ug8ix71NtT3c5WYCMu+cdUVnSrXMBHdK
6J92jf2VnCc0x1lr7uI6KizlLffhRxbq1LQJQrcxP5gd2GE9/+HV3kT8dSY7mkJL4W8U5A9NnHYM
2boTVdwxQGc8hdHK2qsYdLavJi/kL+WCu2UWl3+HiRw0zfNMr4ZOUPYOpZUZJ8Or/Uv3dx3v/vFw
ety+yFL/AUSofxEXEcmxsUKi3lgbAe+cLTOpPB+M+eQTkxYQ36x8z9cOBE+1oYS+Nja40qYoY/l4
PQWJ6rzrX7Mskxnf1UytBgdqXhRMpE9Nxt1ejLLGPWA7ZHMktwFKKDfwDsU3akAy9a/6sf9cyt3l
hXSSKlPMwApx5kyalFNjujL+AdfAAJ4IvT8azDzqfGjiYGb9i6v0NUOLPlTQwEv99IVkUJulxv/W
aOTLP3OPfTr64fjjxRhZOSbY9TxA+lnBC6MyGNf9qgk9Y61hu4znhyKHdIx/Jr6OEpYup9icAo3l
cybSsOHPaenUQgqg7bB4F+e8um1qxsnyT+seyOnVS3+Zkv3kmGdqv6+kYEnvFhuX6xmIRCoGSSPp
Z8rN8OU7UkJ0qfxau4Bo2V6XORZJvP+8rXtdeqQd4tBpgD8NexJtdevi923rAxi08HNZ/yGO3kRC
NnaySQZI2XnrQwQN0c+Jxc2CVCIPDnMZnQT0ek1o5m6X4hkFCAfGsNWLivL8qwoU3gbXCtOqfDOj
bba+uG3sb6ip8u7WGI2mClIVcJxTRu3L/wEX2gsxtdi3d810nMxuR0R+LAry3GK4JBMH+ywuVGdb
vRhH/vUZ4cCNaY2HLyWq8volF2bi+clr+/fxHWECa7x7tm2RCAa2k9jCW3cyu+v0srS9eO6Zc3vj
bLMqR3bzXiT22F/qvfWbfZyI8pwV3qaX2AxGUb+NLzd/FAqrL+dEb+MGGkz7vYVHC77Ca7/K9U5z
ObraNPE/hQ87Mkbq7eVF30cKVu7lm6QS/6GHZ3QRNhB/LtSb+R+QTzK9kdQ2tqRItV/w+PV9zQXL
OhtxKhtLKUjIa4X3Ldkotaq12EA7EgRikloDhWhgWedbX8S63FkuuZLmVE5vd/ZdnCBPG4UnpQre
XzrCSE/ygYSK0Ly1ZzX4XCneJUz3L/YydDimdvbAnsLcMj0MC9Ge8xIP9sV/CVxjEdSOj/WWBD5I
Zzy6CZvknfO8AQnrxUtfMKcbMQ865sC/6MJbcf0sIedxxr6iglbAS6jMNK9M9WczFWQbaeGaqGDb
K6ssca0LSOsf90CxHqsI1s6CKwyka8sn0CV2X+OHVFazFqI25kRyx+ttwWTZgfb1BmWDVk8KGH0d
ZIEO5DSCNRc+958Phl9jgfW5fI5wBM+sG1DK5Rn8rjiPjdE0EtUsjjk9M2hKDyoQqt8+UfGXb5VV
pVdZ2ZZdGQ5UMSjq4g9VOyNTQnLSXHCtRW4OIhLnhGPjwQqJsSNKgHEMXMVT5SCB86CtJIKgTmmr
/CEDvPAB9hFSRe4oEz3q9FHAS0crOnbk2RcoWqeRAGIgWpsZSmSoWLMQbwPBE7TX9ZjRsuvFGY0S
xz9jsH+8gemNN2FGSt31Cy8gl/0ZWMB3T6JDIdW0TWX2LN6YwDUETH+hTPrdFpwYxoftOx2kc0w4
4EhG1rxNTgHkshYrLabFemY8N1vlcvPBDCZXDvfdko8Drg+HTqnIuNJO+TLHZfs9FFH08kP0ABPV
A/dBiHfHas2CTc8Ae1bDV/sbEsEwoRd+1n96//73Uyfkw7RkVtLE/uDY2rIgkt9c1SREiuzQcCFk
9lWgRdR00cHqudTeC2aEmVjK15H5ImfY77g25DBGFBrfCJMsE+CcBo4w02+UPwISwgE3EexF4ns/
f1z0vlvPCoqvL9VM1ChIRYgSV92LLel8mQ0m7wM1lL6x8H+GovU8HtL3PdijP4OAQfJtZx+4EgcE
hHLSpV09zQACxnKjxynTzpHX/rjlvGtZpSMKhXNVoabiakUK5Cq/uMs42ir3a8rVlWD+zhI6pQay
WOA9AnU9b4b7rR4jUmqFnM9NNzfEZNEkn29idBesStIJ4C3TfH31lq9qmonJlBKM6lkfQ7Ld9qPD
a7rkKjKsZltNrnRLAtdQsoMV8ZwY11+GTt89WmDBh6VinVQ8Kh3CYZYq3RHURxwhRAGFuvM9n0XZ
7EIs2mcWrtc636w9LJoEy4s6ip48GKVu6s0x3Odu/kacI17AmdwH92fSKgBW9udFKwoyPeuP+BAp
W/9+I7we8GgiA+4XgrQ6Kxl1T8JNPNc0NXL0fXNuIJBbgsMsIu+nUN6dJ+E3Mid2H1zB9x9i4j/U
IR8d36DRFwvq3NLh0vamlxsK5rDAMxAjyN4fSGI3/dxPmPJ4+RkadNlrJKHyzHupsyfeboUvpbq3
6xyvPyiY8sMRIDEiEjvHqV6KupwSSC3Nbj+NvopIx22/iD3KGAPRDpRnLep+hFTHMcx+pvgofVP8
hipkhBHbgaASypiP8w0fuV4UAF8P7uU4jNT13vQj7TlqDP/8T2Dyiu0n3ajH2/LEFG5d6ADkPQXp
/Wb8q7+I7d7p24nm82rwMa3yjPn89TNP4l4RGYSCV8laVphvSEQByMFFZFr+xtBvXs2y7otUh1J/
+P7Xux5A5HaGzGdZM3IPnsbQLMvap3/lxg1FD2FkmMA2uVJ4E9jz78tlqASKSGebzKG1YLMG4Eut
ZUcu86z1Z18YXj9ELar8qYtGUwYwHCsgi4NlIXvwWd/qkOmNXGPE4QwsPzzUmkJ6lhPhc1QQG7Qw
WCqGyD0Z6wuSa1kYlcX2gvWQ0U4E8cLJkKJxkbTjRC1NQZa58K/94f1D8tMs+G86Z/4vwySQhhqp
N3ZcFOKGphOHSqwwTFD79BR+06wK++kJSLSieibdLELHtbnFWwMe7knrOG8ia/z3oPhNplrFgdZp
Fdee/QYjUyEzPFvO+MjcyK/DVGmgF2YAo54L2zombq9pQERjfl3DkG1j0LUzmtfINTBJkx5IRh55
/eHmV2jXUojsE0MhCqHFMASXSSSs1INljwLzxITJ0SwgIgCHOe+Z75g+3AGtLxW+12Fyy3T/6ZVR
UkFY4YdixBPLhiB6C1Vct7NsfyhrQqJX1xttzrIS2wgIEFmmJaD9d6qgq3by7xBwhltKNeJd07zM
0gm7g2EPijZ2TqLootSihB7cJWTC9UmxjxdaUTszw85ur/ml4n+9ClsPlaIlGuux9tQaw9LgkfSP
0L2IJBzKuVtMi9fFFSLyEVSxmGz3x1ifUtJv5dN4bScDpA+F1RA6pcWtejHLDZUXE5Cl3fwOyRlk
tTZOefwVNn7bLHXhxxIXtGYrYuBDn1RtiGnXF6lD/dfWSIJNySxb/hd+mkUZi2Jy/a1sbz+0k6dX
f2gSeUL/EJc2pjTqAstX1VyCYyR0zZJVbBAZ/S9Vvw9yJnlYHLz876No9CwkwTIHVwgxHPzuoj3X
164wde7Hx4nBlbaPaLr9j6lmbAquGyTbc6IimBYFb8oXmEQ2iqsJTYjHVl+kE7v/kO3c2kvKlxJj
HHh8W8jDcVjNuUNN1i1z7XdmdvnMCVJWLshoumKII8bK8FYykE2/r4lT2yuzsILCD3M8/9kdPFaP
U3D0S8+ZtwlKQqrP31lwLSAJXzSqO2SzfvBjWqHAtwTYrXkQlox/Fj6j23GMfEl0zK1zxfiDnhs0
qP1z1gn4AmOqWpxFP86VT5+0A0zVhsipnbgvZ06Rpcd6KgICOgNAkmbAXR4VD1SxpXU/pZc48/le
+XOkhfJszpJekrndxgn1yTmi9mc3NtGjTNe6PxUqoTVYKatfwNoy5fe98GZF5srBLpxF2VKQi+Q9
iQsPRxYO8ke29kW9LdBb+lbkxGpd2aHwZnmkq8lKJ+LzEuLIRfvp7QdUaSklh2odwRJWrHfhx5Rn
NIkwyWS09B4wi015KSBchUy2dqVy+kH2DUdrJPwNzm/PRb6dSH2TlJsEOVjMMQq0S13oIYAtPz/T
1RXX53Udgzodwo7A62OXwULNIhAHV+R6vUmzOWFlECUExuE0qlRKDpxFuRIvn2UBhpKzwsuxV9mQ
aYpqtOxP758iraxKdbJgcWMsTjJHhxhwOlJXlhj+ABT+z6C1iVS9CUFwEE9RENDZf9KdfD5t0kvW
Hz3PEdvq14h6zmCI9eh6OZJisnP/X6CphBHNX2DCHQfvs7T6Ywfr9yMZDFt/qyX3OUwbYlR8iGxm
TbPwmkhLjMV+39fU11jIlQ+5ZgPOwr884/u22nkmHQXZ/4Tqlt48ZCSN4RlGvV+4Zd78aBOFo3xA
gWns8MOlI2tuuPGnrYoQKlA8Ecj1PxCNTBYUhkrKCWA0DoUlMHi2BhUXkifph5VDE++AaYX4A7np
np1LRftjb1HTDrzT3nyDEwzuHkLIkGmxkxrlfwfm7o0w8y3u7sfiP8mrycNrXVgoDIjcsOrp1OAc
LWsYhw9JH/maWP5dacmX2MO+nYv9hXv2vVU9fZHtkW+j9PzNA30p12b2QLqDM82KjOest+z5lGEH
5GfSx7yXTnVhpO0UWyzS2SDsPB7Kd6533/mrCtZc0RyK8HajU/AFb1bXX7+tyZrZtFUMPx/ugmit
ii6d9mYbevixuIcBdoHxf9/VduhwuxpIn5KTemF3eVuMy/bjTa/YcvMQ/F0dRUUq6ffTmHzwZusE
P8vdtCJdc83PBmIehMFyrB+quOY8GFfB++zvkj2DuH/cOarZ2FBIQixEAh/nip3R8re/sy85g01K
XBnUOXb8vL4yKGxXFpDY8V/bZu0iGA7teE0J1shto7cyZFT29oDEnsnHAXyANh54f5e1qSR8WhJB
lZH54oA+A4lov7MA60V/HNMe7in74QOoOGgEACX/o2OK/0ORU/WxyQuHbjw+XOCFphKw1QTvKgwX
gAKGBaOSVggl7bJWPUb2l43SOWfBtVoRslypK7EWy67nMvU61HLCCEZLAlfkNVkuquqD5Zuq0i8z
7pvtdM6yoZ7B6upurrG2xlt8hHENsx53CfhfUqHTcc3D8tFk8IDhNA+ICaV29jJcVer1AYi5sHuk
dCh2l5xSXRKkw7fRxIz48szwthLRmnsN2AvDauohg5j1w6zhSdUxSH36lujG95C/NF/OvxtgKvcD
0OYnJyA9m6CoA6p6MgE42tIRpUyYIR/3OQY+6zNs8kn46DCnU+Bvg58YoKzO7aRGkIr3Aj65pSzg
Wm1a1kW4+RTg5V5VO39EdO1f5v1Cb4BlAo4O7O5F6KS3IteSxQTUvdvxidyLpANZzh+y6/ywbGak
Ym82JUt4sJc7o6Z5iGAvfC0OqRnByTiWtkCfnT90RBawmknNnIWa6RDfHIYP6ZyqmSICuZjXUVi8
kCMGWkdo9SMma4aTPmtnSnaNgFDEQMTERhcixrrbJoP/egB9AaRSTLB/Z70UEfIg2IdeANe/vcbc
IUR5SnvAq+tuvHlSZV6AQ2j/b6+es+2znFcRcSvdhT7CUlK5xbOpbEzmOb4UWVDp9z1y7rSQHnYq
NyNHcmM/mgELJ4ZPYdLJxHBaUpXAMpQBYGIxYGV3UbHPCKmcmA1fYJ4sOBF/5D4FjmGtVJI9V8Gg
TeHCRiJt4Hbs4YEXRlE5WiLyEYK16a4TglEmgkk68ROs4aUxsdSak0KCipBaOsnXixJLMnCxEKso
gdKDlbdXLN2DnQaDbIyDQAY2A/FqywyU4yM/5bx9i7wlYqFsu542J1vV9wWb0GWZzWsWaUTZG0c6
3NFdum0EDkCnu0ll2mfVvIFBzTkq4Ob+tCn2i9uUMK1LQk2P/Gb44DFK2k8m4qGyHBEn+Zk0dqh0
1vcSyY18fN9j5/nf9dWcs9NWbkJAvz7UZK3Iw74JZcjG3ppCjfUO/9s9yf3B987zUYdCDQq6KjCz
shzky4q4ko6x3mM55OvY6OOrjw1qbWrPhMRjKnOKTCh+VWK56UU9VzpV5W6w1W358nwXx7dKz4MO
mCwWvwn+OOAKWdmq8OmAy9kuvJSjQTmgXZI05LzvB+TR3Vo5u+UJ2TFeF6cZjjymS/X1L4CHqpFu
9sBDebrRKI9OQvRyD/2biwMDSCyA7kwtVwp1vwTzWfFVM+LvPrzV1WaMX31t5MLqqa87mMTtHtkJ
zQiKxi8DrwV1JaqYZHyiKb+IKl03G/3cEXi/ZYH+Z8lSTfNaPLExdlPMt9X3iGy20HXroiZtU6cE
tyqo7P8zbV3N5vU5AxcEoUivWwI3UgTWlAcXpyJ8z4iJL8/nNj1rvhXL4miojY9/SrBd2xoSh8y7
0Nijn6Pjbz9HW+bAfZSD2dUiDfU9nkJRcaQf2xphpeDF2246Asj39iUYDqQX5bG+YoFHAlZ41oh4
cBjyyI/E39BRieBAMBNlasH93Hc5SQw2gV7FNq+/V6rRxcD80GXamIrOU+OjDosqZk0NENx8j0uS
Sy7tQinEU4XYujd3QLHEy/pzGCjLsCQu1o9hibKqpMiBlhObmfKqUKsibbYwdwpXK1f61+W4oJkV
1TjCuHvW6ZkAOa6d7CCw67/Mu+bCG4a5AdbQFqbvPjFox3BmtO6zFlYzQlCuzCNhkj7rWHUtxkkY
DC3LkC/YtH4xVcYOXHmxJv42Z5OjSGgCvKwYFFwTgU/SeQY88agdJnixRcQ/UubilB9I2XlCUmKO
+j7AOB/XyC9FnqJFLWAxE+i1fVJIAxVB6S+2g2VKmDyf9CsaAU1Hy0hRxLKgEnCzHeJ5TS9Iutme
DAspUp7NJg5WJQZfxqavDxfqYb8T3p6Ak4hL9dVhkybr7lWK+U8k1oM+O2hrzeOBz3DFE1OMoUOC
NwgLUwsO0fHu6ang1AdjpbjZfdLnGRHrkd3+JvQTvS+vOaKW6z5Rgok7OZoC+1nTgOPioGcRuPxI
eEAGvRO5sJ5NLCf4RYSqqTCkn9L0Csyh1r9VaPEirlNBzy3y0D/1V4ivzkw95RU8odOfLK0OladA
FOwDKTD3Ht0qwyK94NfP1RJf1u4lioWQYtIXV+W9yJ6Ofwm0mRl8usEp4s5e3ZJPGDpDo/EDA2ut
L7COHPziuOjUbeMK6JIvdjLTVYGjP8rgp/W9E8Dg5eNU2zr6I8nh1fmnNn4rGTNC/5sA5RtV+9Gu
v3HeaNnsdlk7AM5lyxcVmD86oFI9iFU0oVMzwIfkJyIhHJBxp/nR9RBxPppdnYlhiRTR/0EboBAG
lsgkZuPtAN3x61jcpeC7CLdwVj/1hDoNjcoSD6hWEf0YXSWswz3didCdvQ5ObpKumf4eWn8FEqFT
YNSWeedX6EEIpUGmuYotaL623dhbbLV5/GPbxc9iO0w8NUw9kfb5LRWunPDr4s4etTQd+5ayCV4L
jpqVAPLGCagDP517Wpb7H/zMjlvdVCDXfkPk5KOQJqbP2/MzzMygY0mQN1i7C4HISBqtAgv6r6eh
zqvzlpmj/QLeTJ8JGx2a0l/dPYsdN0b3ZDcFJ2jbjfbC4tXeIwvR2aggJ8n7JUJmKhFUbDwC5s7X
OZbscMiA8DfbJ2fbz0Ka5s1vCh92B8GpNRUIGfQnqdO9qLCo/zFxzxoyrV7hVgB8aTOV3VtumShw
R9BUHppdJ7stdJtRGaYioe4L0wVa/uP63SN9FBU2sQtIzV1wF4o9fylGlhP8C80Qip4GeV29h61a
XXZB1j78vwazaPEJn2fLGua72y/QQREHn8W0tmlr8zruoAXtD3dbwpXmLthllzibZeordX1RGI1/
9sc0/mhnN1hmvd+LPqKLUMdpJRImq+VxIQglIhJw7f8KF7o8EayEBTdnqkywVLx57KiAiFhqFF5N
vdB0Bfg4CY9d9uDcBwYZaPoS8R0CLLa9SFLXwIYZaOAa+wI8C/ZzkpY+TeSUiISTZOpYfoAsDQzx
IEUHF5+qN7hWLPd0m0AIdxv4UHujE6+/nDJ8N3BheMu54D3U6ElvnywB2tbsoPHbo4TWL4SoBt7Q
VVFz7SN1NX0Kylvyz4sgTHUUrwVaEKoBCv55+xh8Bhk+XwG1UOx89bsgJJuvQtWdAEmOBE66f7TI
fENytLkO28jWxzbauBzrgBDUBhLaZk5Ah1XEGpt78kaAZwE24iB/5ak4DmVhUVcBdMLSf0cEJygy
0fxsCxYsg93sk5k7/5FGkJsouHx4wFFC7zFYrfyOrQ+ooLXve228OJ4rVR94Y3hgHRTU6FrFHcuo
s5LR+9x24CsifT0pQ/LmXbxo3DI0CNRls+J9r598EnzZxQD91KS65L7Wy8K4YR1+KCKsZu7FDOdi
oFjq/6qNSfiNKsZBmPUMlfKJAvXEG05XccVroiIOC9GjgemkePzLoV8cR4SUGSIPFZbSE6Cmb1Hv
LbBTaeiVOy+zvEnw0P47fs4pKF7Le0MKfe34gSnCtSwRQj/mFCOcnPJyONm5OQrjRiuZzPZH4wya
RaMs0VZRDXBsfoF4bOIzWwhQPALUldXPxxFevtYWBAeNbfxAbDABE/U/Nl8WinTl9AGjBo2MARW8
m263KVjCRKViIeX8Ms6MEqufaeENe4moJctwc24poqbFjaMSesDHawnAn0rVZt2Gx3MXGW/FGOyj
1slnnggISbO6rjSNFKLv1lnl50vPuVEM6hLFtw2oeQzsiC+m9gQcs4mJnLYUA5AUb8eH81LQSV7t
bPk3z6WRCkMCRiBGYD2bYrHp4n1PtGDaaWKpzoWFW48xN2OfoKHp7UHaWm0yPPbzigHoPwAxpM/S
UxaDqk/qjDxhRTYsz3mSpgsYIkxIj61nbSPFaVbe94LMThF7mLyNHmjKQEZjHQNSV56A7jvKEqRW
ZYebED03TXn7SK2DxW9S1NE9hVHsOjg9ZzMYiIh5hYoSYDI3jqMzhtybS58RdIplB2QmQoBLXOdP
NlGeppXtITt026TiQUOA1RZIZu+IgBm/Vfhlp2Z7QjYWrUU9gAjnaMG7buNo7V9Y3RwiCViGE1Md
WHdbqEpcush3Pke+2K7qs8YPKtCq9btoOpa0QxtbeCDt8nVAC5NCVXOr5Scbx7UzQsReVTIeqgF+
jia4oj+8qyTN/7pga+P4B9rEkK349fbKTIDYt4uavpElfMA0WerQvdCHhDHCOMd8jvLdPRXUWHXe
bO1rSwqoSX0l3HPwdoN076iim7AB6XALUaERihXZyvkeCEXJyUJEAmY0xTFTv6yPKWZDrARuzW/E
2Bcpsn3rlCrCSwtGlXWmYf3Ynuevjt179Cbkhd+3v4d3E8k/XPWkwbnWnQ0owVebN6PTIJQm3CY4
Zj8kvO+o9rjL0VKmqF/2gUwv1RuGt4qe5Lklbs0r0j1o7GVtlQFs7PlBTF6MmQaO3MrBxT85SuzN
uoxjU1hrpfejVWjhxgLTLTpwBwR4A/vYf40ntDPKC+jOq4hi2M/Pt6aaRJQbpw8Cvee20gmfCBpe
7jlxObbgQVoHyi97haVKRX8XbJpbmq23qVFMmJc1WAWvmABTeOA0BDyI5Sx27QFym/Gr/9Bqjzcp
2bSaqHzL5IlTgOIrP3+cBQhZ34sP5/CRGFYmHvZ2BwVo8YB9yHd3U73Of+sWr9s7/yoCfHms6Mob
ii1RdN/0E0dlYYjToFKSShL829dx0U2SbNKfMnmM9148vH7e0lfDtrajqr0csE77oDme41X3eOJv
TG6XuivH1jPdHU+ddtpt8CStRmXcrybV5WJKQOpD5+C5J4FGb3BBRUvpnPN3X20KROqz4jhT8Wbd
WomRrVOSs/aAS2uZnhxGH6N30CbBkIwAIDOvtHA8ElQ6GL/r+hFsb1YLiMeQZuuH+lqETqST7uIY
UZcX0WneShQYQZFs/8XDDYkVyiA/wN8HY55lSI7ihlT1k+IAp/V3zuqSI8kThG6YPE4iQbga22CI
0TJuv9XidVZtSSUxmquzRkSQXWKoDokZokEwOxFOVQ22uwWLYXCLO1LR5BzjCgYu2IoQEEf8OhMm
WVHRbL9sIDTH+mkmKlr+65KNA3rSrKg3dBYhdgoF5oud10frL8XHhDF5T9PcqxYaDvCav8eg+HZn
BiHRJ4TOCo7iS2PDXq276sn3WeX7XqMyImOUncfBKtYhV3i6lBOO/EkHUWnVQuk+gSgs/56enIHr
8VFjGsgZSsdWzF+s2M8c2o5CrpEhYNFdUfMXdgUOdBEXssEFX3XQnFT+gHvnIW4VNvkm7ELvOvgY
ttqQ23RIDmn6iFzZm3p9hq/kF/OuqPiuSm//6U+4VOrWv6AvFb+nBKzWexHGvFNsFQN5nlbkZO1y
MgKaRl0d20ZcNR8ualJ6lX8ws/GjrcovPZm7uS5rkc1YXRy+g6+6H6Vc+U5wrbYyL2uDRhMrF4k5
TAqNWxxkxSlplAyalZN3kbTta/GdDEFs6JkEUsalpWZSMDwrT5V1JI0n82rNNBE9Qh/5sOE7gkye
8fT49aq0/PKA0wJxZInjRP8fUxSEIFlSAs+IjUuvVau5vRkY2xqcF6AW/8vYc8otpIEZLZapQ+Rq
ew1sA1GyllOqL1qV0nQCPs+gpQZMpz1oEcx9u/E8qnaMRVxMcmMdPmR8W1fc+pNQlZ7tgKfpaTS7
JKn/gQkh6qgOhShL44G0w9wvP5QQNzlTWeJB7J3ER9yXncj1Ye3K53ItA22dN3bdI1fe1cRzJGue
BSctM4M9AZ5SiJyrXHNyuoKWYDXDNvz9FvApOYVmhDVGd1/IbFZyb3EtNlZaoaofSHIgTmZ8b1Wb
4ZDNhKXVtLzqC6QunzzSNUbcYwxphWwM4qHadI5ImPTVoWmFWX62ocWHHR14D5QRKoPC6cvcAswy
ALn2lAEQYGh/flTIkINPe++9EBWr3N0esHXA2UyLZeUJDTV9WPTNCR0tBVJVBqthc4vHvecERJ1o
JSnYfd5f84p1o1tvCmE9kE3dbnGbuEj8UTJufgCBvC9JAiwczsmsupusuUfsDtdJYbZ71PtTNvcS
HWER/o7P9jYREUWe7HMQprDWl6rMpV1b4kL8JIxSuGehdNVDw1ydl9C1LvvweVjvQfNBFFTneVuo
ERbCVPGmujlQ5dWMnwHaI3vEPNWvZp6+6s8AVZRTDFoGQzeGTwjWKd3KJxLyErdsT2UwcfwBjbPJ
AMB03JL1BLwh31bitFccQds4fBfAy6UxCJU+F1AJ4zr1rrZi5/2LQhQpQhb86/fd4YGQmFH3P+pE
9UQW5iALg5tK2v2iKV/xO9F2DgsXLGXprFH9W+X2BqIYv+2hBEWg8u29YZtd9Nzs6pmfquRnwpNF
934VSOqp5gslDPcTUpsjtUWb/wzvz2ubWDIPN6g8hvyOh5fNLEGbCzxj19J3b1s7/6qEp7u9XxJg
/y68muwNsHYYCiFjWd6qAt1MUWQiFdE60AgwFC8Lh5riAcI+fBEKV8LCbdkyKai5Pn5H6q0N3Sdd
i+ww+gf0NVhwW+svv9/LTJLdCzqoqfhsWpscgwlb4T5zwUpdLf0NYL1yPWP+gNU9OuIbWkaLVy2X
xB1vHj22uGQNF2kPQrdp1Yrs4kmdWMy3Q+QiS5H2Lgc9zkBooVdKGRErQW0DZVH2IvasplhY5Oo4
vx5brs+CxL5yVAztahujkBrWHank2Luow/kd8+GYGcncEYL8GGf8FmQbLwVrh+asAdJZSf2vhsI6
8AJSFDQzEmtF2wI/vQeFwNbK0I0IJmjx/TnNiI3kWI/YfyoL3GbggFX35sjoOYr9rj77Sa0IGD9W
HJPjYJtCuehf9eB7cRN14lMqdYsE1Ewh+3uuysvJb3TSOUNpaN0cEQFMNQPfQQHAgLdUdXxQsYO6
gYGusYhy/Xt/lmeOszE89Al3IUO81d4X+JBOH24FcQF6nVZLn3FhWJJUrYO5hTSdffwK6nLHtyLE
N6i5FjaV4GUGtq1/QnsbkN/wGL583o0QgmDylXfC69cF6e4LVFixU8Z8ciI9cVhoYDyH4qHPQ/wn
lGgoD39Rzzlx05VzJSnhCBX8ISVGgarg4O6cjPMNYAFNPDEXongTmEeAGw17f9lqkO5ZaGEzuEEu
YRubQYHHpxyUEUfKO9YBjHLQC60rMR+ICSjAHG+JdAHg6jGZHdzR+OZmgySbctzk/jfwSwo3mqjX
2ylK8wgnJL1Gj9KzdC5iwUNVZIEBV4MrJm/nvtWP94bJvnLWWRKzKuYptxsRKn5uqq/+bdPMMndk
CmBeP1cT739qp0FdJnAImYMeLII6ow+VdgIAtdEVV+f2c45P9jyMuKjBh6103IWFWl0ieFzB265w
6u1jrXbNSlYCUO597nuCDtcOVzN91l0HQ9I0Bm3TerXqSQ+1CG2EXrGOa/+26cS+xDeMELaPOpD5
EU/IDZTEnl7g7RbpCylHulICyK0AmE7r9jU13dj/TI7VwNjTMwr07xmAV55iMDlfzTVHVSlrQXW7
dHAuC0Ef/G6SnFfk3ddm4YvPN+1+ruyqHH6FIuNHwK1Slaeh5VlrXYisbZ+GXliaNbgpHUP8wO+c
MCzmOy6+GlPVyWTrcAVcvxXqCwYgCbL/XSA9QPWKUD8dNfJhvu94hEra1qG8gKnJQszAYXQXMv0+
BRp8IBnj4yjaAL9YQ3dc3PrRs0CKxKVbVdfwJ3FqFGMiquEd5ZnxnKctBocx7rdtVsndvo/krr57
cBY/wCrjuzRID8Zhe7xQWNAIoDeJu70ta8dWU/SLyKTCZU/OKoLCXGHkKNF3LHCAZjDw4YrUsDM4
WYKqTQCHGlWuvlEZxoabPRqRY/8FlZl+HuLD7eNcEa5clcdqv93M585vnFaFJnudmtoIX5FT6gpE
lPj/LKY+dKyRhbjwZ1iGraJFYhvd86xXhL6ONZITvYXLGiHS5DNYPw8z2SNfSMI9/kIEvV96eBYt
nahgGL5V4v2jEvfit91aQUqum9BIRzEO/zYef/i9v5NZFdmrs2E+1oSL/FeJmx1LW1KZuqtxfciQ
pzlGEJcfIWS+3RT3epE4mcwdVlGt0Z9zrK1TLXuaL8pir2Y8v4Y8mj4AvMO4qu3MwmiH5A/DKME7
w+NNeQTSabaIDgJ4CDeTMY8f7WAQjU3N44EUnJRz6QiY1WQs83/SqZnD2bwy0DXvTYzCUDtdJVra
81AAmW7o6Bp1lLXfgT8yHyNvlJuM9qIPfeieRr9veyx2xCpgSgNz5X98I6NeDm8obaetymi3QX6R
NWaMXBymwBp5oCL072fwmBBGyLIfL2XrA9PLvFdJbxfgFJtJqtG8J+j3Oad+O2XAYkbfBDLBPwzU
7c8uaobFwN+OsiSjcM7mQrgb3TbQeL+GoPUsYKEo8V7KvcE/FVrVFIA+nmjL3awfa7cOSGDaNkmL
jif1QnQl/YD1bgtQ97bks1F0xPTUomcTZQYhVTaeqcu9rhfWWFxAqoYYeTScZIPLCPAShSTnsJ7k
kfyFqZOH3iV2s8RoUZEucaJq03c73+mijMdlMWULqp/Hd5zTUDyDimZVomU2liuzbNaOn0KS+62f
C4NszJMV9Fe59EkXoHIn/zv83lpc+pgvVMAae+yN1D2xJzFWmdFlDm/4xa1YeDT/qjYswaBpGq4K
WdaPsV8nJ96kunufGdS81DeQld0nmio670L6V8911UkwOZ8k9xq2ibxQ4Ls71sI/FiicU9esG6/s
YkK2/6ldIQZJj7LG2V0ErqWMs8UD/17ai4dxK6aPiKgLJ2L3b8czlUEk3VTbLEfopSgcbQ8o0Gsz
fDbn+e+syBoN7OhBbeE2zmZYKTaBL3g6VvzaK62lrCzWx8ZReQtEEKkLWWCQ26KPcHoKVYAAvo4j
qr+Fk/uvb/ilH3tcfj6OLAE6DRrWYb+QzlZO3czuATtZtKL2hII6ke733DkJ80B0xo6CUzmw4zGh
ouJack5q+EXPKIApVknvkdVqMwhP60mH/BqinQySnZ3y/xSW9mereNfAm5gKQkN6C8pmgK1VplZR
3t0AkTIERpzdkf8Etn/AqHajqP+3WU+oXmjEjfqe4QYiojq8RK0iHjjrhhZCcTVil5CTbjrYQ14b
VADdqtQX53czy20a4cNvxhoEeaGyYjjDgW5dyJXmTFE7GpGGGgKU0JllivzYXff+tnv8wsaxmN8F
jLKuY0IXfTj65LcK0jAs0T/h88ZmOx1AQlKxt6oteUNtXdDHwX/wokT9we+cHlV0tDbCyoa1Nh5d
TEj3rxRxyF6H9j5Gl/+69wap9m/cSCVVjl33RUmlk1+UyaLfm9xQO5AhOXYo+IPHMsq/KKEiREme
u0x1IZWGYtp614SrtGxjAxgwBDYH0GcYN2oNBGwRVDk4BIqrlqmE4D081jHcmc+WChNeb/b8XsZ0
QJbexsXMHnaez+8hVpEN+yaBEDNgBw2w4KQ+e8lSpf4IfRABvB9oqALcir10t8MlR+cMKvs2aQoO
d2/m/xohM0LMCNg119czVtXDFQbWsi4pbsEK856GXgQbk9hnBr2Sq53ScFlMEA250PzJzpwW8kUf
K1exLXDVqtSRns2Q152P7jNbYjZF+BY96R2j3ZTBrxmfIGv0HwTE5oJZQxHo2Hh1YfbgrINVuiYO
87O1ZdOgxjkJOgMQFxSKEcyYvyLb3CUrZBIAxc2nVbkbtr8///JId6VGKBZamYz6sg+RbgYoJbKj
wEB+3ioAU2SvgtCxTTfGwTNLWrYXtpmFPBD4TDpRxUyQ5Dn9ldunZLFK8rROkka6ilNeQlyBcV4M
bWelujptwqKiPhYQaWDYc6x7m2B/ZE+cXBDbzUVDZm5VjocnS/CldFwQPCF3/Bw1L62XIdgwWBoA
dzZcqpJXydA2DUFdXybkwsMlv6Q4C/6qd7hDroF0qr1uf4WgMpkia/Wk1h/83FVGyWaZdjw7fVyJ
reu5pAFGr7GlgGh0a6wt71KYVSlH5zwt5pxMvrrQnPBX9bfep349xlPeRUv+3QzKaIpqG1C367U4
WCRja0l5WDttSGyzUTqc+jwadnDH7sfsatCi7sLPX1Q8X55RBctmz3VkhL5RgngjsYM4yeo/xAU/
Dn6/2vPWVCxQYNTXw+RNeeoXQpkNIjjfC1TB1lLwUXPOeYDrPRortCkdke44/2r2rgTLSxgzo9nT
e5wamWdz7ZdJKCtOmbppimoeLtzWOQ5acvnZn7WUKuBcLb8/5qXqWuJMqEJDM2SqnIfjXCBtL9ly
QmrLFB9+YgA740NJGNXUGt8tz9rOr2Y0LXjqv/QKXFa9TM5gmx7lm7KNnDrZmU6UDfYplXK2wsi8
dXkLRzp5HL/bpvkxduNgOl+vNBp4Q8IgcM5voIz2xUgbyvqPmnju6hnAx/91EmY5/UiWEJhT9u8g
1y6gblXnyjMiXGBAz8zzUeFcjvwmQO/FP+9qNRIcgkxwZX7q3Gt/S+UexTsBunPllKfzF/0I8vvU
vwWNGd8BECZBNFMtD1Dj+X1Po8ymyAWFaIpolTT9PZKx6o1/QVU+Z7CuXjs0IJi8yHvPhjsxhMCS
+oOk581pHykniF6k1H8OvuGTds/0wvXMlggtAiEHeCF867n88B1tZM9tIxEBCGEdDfnEv+Ydqmdp
Mt132rmlEqrnqLwvbHhnRn20AK4Xa9J4VjxHsVdIiZCUcNfRlPQuqbgJ+4yRPLHq/q9a1LqiNxZm
vPVWlXEdS1/HDKgX188cA2XFuLKOEKF52sBth4FjqIWmo26jtTW+9Jf3xqnDOPupWencR4GJsVOl
1QF4rXG55HDj7B1AIHjAHdoQjtQZZJFliq4EOBu6vlBZilksPZqdv10vnYKKDgSVdOTITsx1szjc
zoZT5hjsF3LHBXHO7GHjKIC8ezBd45n/vHDlxKYdISqWsqA5Rb3GK1lygMb8SxaYeTXMMtyfp8YA
A2spY9I91QyEvy2lRUx5/qKdIJFXjZXKx/8U7s4EvNnX7gCDaxW8NJINh3XDNOrJxu5rZykcw5ve
TMi6b5uTVHBp89e36+zIG/FHhlUfqd7wDI8LQDbBeB2pa9Hrp8kCXrvZ0d/d/WnLMsxqKIAwJkr0
ump6Pgm8QCvT4v3ECtnV2z5uJU+SPKA4ePEO2LBG4V0vcFMJtCX5gJ/cKBbs75+7fz1llrk5by7Y
6R5cvPCf0J5Df7kJgfx4/BBmJ0bGl7OZn/OJHJoDkK2bJqUyHJin8eY8CZE6TVrF8Zufs1dbCN9q
QmVf2wo80hvVYlzxeEnLm97/0wVo4p0aO2j2kJOwYfYx8q/+GQdO0pZi3rPaPGyv6q4FFrkGS6o/
Zu08ps4KpqInGnxc42lXKJ3xmPMno2v3HnkZQ4gr2Zk678XaeX4D17R5CKkjGQ9yUh6K4HZKUocQ
nqfjQZG8huTlA3IhsDapCZiTU6kaIutEA4ozgPhBDZx1X73DzYr4zAlClQg7kGrE6Wr5+fbKXuyO
wRthsMouHLZqGW+zDGtoAqQaGWqepRCGqJcB1le0u8O9+CGbY3ZqjVuwlp6ioUHC2TKoHFgcCUyr
H/eBHQpXYQ9Zynzg1lWG6TCtVl9gkznUkUqVwzzvuIO5amWJ9+0VJS0VvpzxM5p259ns7lEKHfXE
9UlzRVA0H8RGMJyBsUt1Gfidx4LkkzOKCP0m0CITq/KqnAHqBADObFMe6cZc2CJxDq7V3C5RcHQ5
wWUpMBwpkWp0pgN+X31jh7n83IPBam/Dvykb0Fi25M0kf6I5E8E3sobBprZpkWfQl39C58JX3YZH
dLTqsD/6iwycvff0fO1/oNm7nHXoN+xb8HjyOAxnpDNnzyvvSCndaMCttOHuRcHFKJnCeAQQufLm
CGQREGGUScvy/WmP0bX4Z4pfCjm9sD5ttaylZLKN8HV6ohEcD0decmAmU6iW3PfOxQbJbN0YDUKt
oh2PefD0A0wiaQf9lJqjFinpVJ3AnMaiHyb3FQba0NbsAwG816g8QTKn3Y+Z1JTe9QIkMP5y7BMp
nL6fhdIwl2Sv/qB32J9eAafeL2SHdcExvr9F4hTDJA3TbdGm2Mmm4WvZEycaIGiQkpAsRYN1kT1u
pfgd/lXDf3uj6fkRNIGwgxGA8ovQpqiUyMWtasUMrr75eJ+IyaLTQ4NqIW7thyq6J4Ve6Z8dpGL8
2MDQ9ZrY7YGoC/tnK5heVdgiU2e3Hx7rv+KhoG7AafAYPhTVzDKXUIpJNCl0xkf2jYssYQmWqAyF
897aOoAv78XW2yj/BaPube146FUbQk7MaMcy8g2DooAyBHA2mgxhtPIk8eEsjLxDoN2QLvpitKip
00L2G/KLJ3iBiXw+5+4AvlPh/oZBxoT5OljCbIAaQegyAk/8nhd2naSMfOlzNweFAQNocMDWIFB6
hpz0qyc44cZlsZdNUUvdPUCXaUSibU6ncX1bysld2N7LeoaM+KdNa0FnzCS56LyMFEecRefhtCwg
HDpxnecs4mUhA5phCMpP4sskxJoQLudl/8DtqMtJFyTuOuCxgCaiCkBcd/oDe/UXl+2DA7sNjCLB
PrSPirUFPlZHkWs732OLQU8PzGLG5tObjq2sqMJ3mTeKd60hTgSYGhIX/b2GlETNXeS1caxbyhml
X00zf0JKEAftqjSPnWAoDj7MKg3uPqdRwcEWTSe3BuqMTHZ8m/xG5xRP4g1O1qcjFaWVNj+iyAyE
t+u/XyVOnE3HOuPDyX5xP4/sne1Qp36XC6tSfiEFZ6bLO1ko1mQGBlZ+9soZbnTvs7XBgOoNLb68
E6BEwAZ/FY7Hi65L1H0KhOMokwPhxJG5sve6a5m/yDNsBFbgHF/Act+PjoiOnHZ4bNIBwRnQSJm/
Cqvs3ahiSvuxsJFoAYQDpuRv50TRyPw6zCbxdNanwL/xNgiLvaXQhm7f8XLnr8m/ttqBeb/mtqtx
3xSNAGYGluLc984enJysqHkIkkWjIAdkbJCHO2iYs3xzXPjo6bWmw7L875auNv2fJ6dR10GoU1BT
x3eVAYYizNMBCOyxXzM6EQ8dEk2yyCsocB8+GxX+/8xHIxs4pGcqIBJhT0Rq5s3XjmETTQKrgjeC
LLFHYyhvM3y9AoGS7Jinl2NBhK6M4UNFDqgrBWmuvEgkwZnB8vD4g9Wk0nF7iitJd3BVN/IqAF8c
znRLt551DcVZtWTzujS2sZm3W6VJcFvFdiU0YiI0i9e01J8E46gf/jQBnd4YoM2yV8soPqcWv+tb
vljTslnVysnfNwu9rbV+Hw3Zz/X+prT2kuQiKCdYDSlAnx98Na9Xr5MniYz0wOHBp/MzUftdxU5d
A8l0CYGcrPXFI/QxrEFw0KDB2rPar51YH6e8kONDTlNYYGbs6gksbxCrVEk6+sukvIlKMqKB2l/z
3UchMyp3H1S7B4R5OE2i2zifS0pDLiYh7sD/dLmfgHfclcADmPDRinf0QvZpSD8ZGECZadABr4q9
f4wGwpM63hGwXduJqreJ4CiupP1XfMta7wC3fBbQFhA5qmKyWBHQOHkR08uAvX2Tv4Nv6QDwweLC
ifTqk9wYfs9QRbWJ/2FbmanVX8GXbwrtVztGdOfdU/CApySPu3oQHztX8kSsxq62F2WdBMiF18Kf
ofhzLbWRDHQnhDwFDL0NrkONEs4AE6kEQDn02LKByocKXmjlpiQjP/ZqjWnPR3PX2cfT52AL2lgZ
5SrW4CfTJlHGupB7h6QCd18fGeeiUB5qxFqxaDdYxwnqSm9fcaObOsoCYLR8tn1ZwJ+tWJ6/ra5P
ziOHPx9tHq2Uy1ihJLWxwH/0bFfePzjj9382RIcLmhYH5DBP0jXo4ELPMppruF1t0PXapE9wcQyk
oduqj6+X2lVzkt2gU3CCmR62orSfmRniruIARRqbrplOwCt3A3OXDts86ia9wEFegpT7iFn836Oh
nevBp5K5W7qqw17NtnE091NiOFioVaajCMRW7D9dQm7AJGKq5P/kwcSk6niRjSU34n1PFFueGFne
BI007XrKe7GP9zaSGp1iu0BAmLtOGT8wNMdK08LF7Txe/QTvK1JmtTRkZRMmM9sgLfi3EytCdi0+
OOmcRWBbTje/DjJoRj0l5nPcyyQMtH6IyIEmkHHqFaQt3D2B5uQ8ZO7necNYlsz8yuDc1kIxN8S6
Uul7yGjyQjD73F0e3+KoSBGYI03QvD5O7S4E5zb6Emi76ByAg//TKtNnV+pCw+6VhB6fXugi9y1m
uptF1ya0/mEf5NDP1gk/0kDpHNMC3GidG/x0y1ttpZD3US/7qQZF2ymU+c94BQ+BUmEp4SUtxQJa
ZX2y1bE2z4fJmcWsSAr0BYEq4En+dbZCcxUpGda3nozMYVE0BpgoJWNEf48eLrpUFSRAA8s8UewN
Qz96SEVfx54RMN1beabV0bB7HS9t+bDUwjBJKrcVt9ptvnwbRJBhe6xK++dTuRD4DEuTdQFaB/4y
cwG8yhOrr47flobGe/kulDDLjI+fcTipYxfg7iHGgFUKM+I0Q+73dyHee+4Zd/k5Xd5fje7U7LwT
+dh9dntMGzV7tijI7nqrhDTKyD/LI1waHZyR+nSl+ZPo4NF9hRRV+RYQpHtx7C0wOs1jz6R8DYqH
medl68x5phxdhd/EJ4Bb6SNCI3lXatvo+piuetm19O9A2D3vkQuUurhC4qVaSe9xz2+yhjr7U8J+
7ou5olalE1VdAiwGg1b/E4KPO97bCl6OpKuDHqwxdymqhMGOuLXshQUGRxSF98k7KZ37pRipRq5/
KFEGoqJQrqeU8KFrGy1cq5cadJJ5Nz8MDHwlN/guvW4gjK9KKzSi/Is0mABXgTFkcvfzMQtnwOGD
MXtNOlNHku2uMZfAyEliw0y/k76NRHNinK+aSCjPo4hpxlwdUspS8SqcAkDF6qzhp4CKABTmIWbQ
K1e1b3h5oJEzD6dC5LhOJ0ExUGrSr1HvlDApS8jfRcu+H8bCaq42CYUxlslSC3LTdsyDyk/2bZpW
0MGuXcAnTwO56OEFEc58EzpCoCVQXj/SEWXimV4BRcdVGyguZZfd8lqMvLg/U6RLbK/LP1XzRC/9
SABTDe9yhiOwMsAwi/fdM+neGTzj0La435TzqGuoLE0t8KvD9vdSaoXFgsGulmt5LhU2MVll6+Mi
B3E2qELMcOWMQVhcybicnp4C/fL51tETX2W0Ji3cfiI7d42F3nixdR7bl0FjMdoGEw6LiEI0sO4A
dp7mUhILNIMrxmmDD+a+y88+zv4ZgQ+WyrA9yi3bEowVUbF1Mpf68acjDAbFiMzeaSGScmQ09COX
4AgE2gKq9iRMyUfLoU24YYN78jH1XLoomrDyQVDK81uYh6L7B9vDD8ck2ZQWBGm650OrMK7VmYiY
qTgxQn9HzILyB09tCJBP7YASYkdC6cAfMNHCI+pxVNhLzK8fUHp9YolCNJgornE3OYKTlgp457pZ
qTBoaDlNJcD/ke4DhVob9kjTOicW6O9+a+M/vFcd0oh1AEoVO1Feiyncd1ppiDWqyqP8ioVWZrcq
dlHB7K1e6ppF6FaiZv16KHwnZwZDqSxf8Wes0A6wdT9w00WelGYu3r+hiJSA6v8KUExSgmRfs6nv
ANJIRpWdaZvefAoUChIekM0V19ynnfqUYgiPfuTpl+U5ovbsGD7WfsZJs4NPVs9mFDX8VhrmKXkV
3K4qoFClwqkIxt6I99yUsWSYg95m53+mZpJLxNkyy9ER8GWw2LhzBvcUjTN+NUJ2Y2L5eZ0MDNi+
1Uu7yAXZ/+kxGkT33CIs1Km3h22JfyBjPNzMznn4QW0yDkA62wwvgDbPOG/M/CL+RuDTAAjqZKa6
0ORo6iSpsRkE1si7QfkRPP8EtMfEqg6qF/ZNPFDLFhN1Oup0VVWXrVo2qY9uLESYm+EJ6XvssoW9
Z/sY0/yZFri5ewBn2P0Ndvs1FYQUaNNSTRsqIp0G/xhOUkbebtwqIJcrLxryX5YeIKPybBpft86V
yqlpMswDjATQvu/8Lt6VTe7TQWUIOL1YQnMvDJa0oMRc3nIUjrbHCiGh6NoRwKHY46y54sU390Nh
0iZiAzvB59OBGZnVs2nuT1Oxm3ruf7oz3PWksbAycGKw29DgeevSE5EMZ6N1LU09XwHLAzOa7lqJ
ejHaUwaYq/ETd079G+aepjErtdM9OT4Um+uy9BrkcGZOSVrlrRhzQ41IGOs26yQQW2NaENX8I2nO
yfBWCm8SRs6r6OdHxepit9UVEFTkMnKRoyQ5oKJgBrPBWRtruOPfQjXb0LFg8G0QyKHcOt84ZdMU
bDdQHXOHQbS0F7GPucdmNlDzGzXPx/CemKANsoBt8EuwUorfjzIPjyRJW+Fq/2KcSDn64yIriAmJ
V0lOvs5aHkp067pF3D70YQWHNPLdt/sMwirRAA2I9UxKTg+QgfqkiwFfJ+X/ZB9tQDciwWzREhuC
rrtCiadYh52vgl0OOcr6sqkIvM68ToCkqR+5b+GkfkOlHoI0GUXYPcMZ9wXJadDzboPC2umEhoWc
hJlFDZFRTVlafHEuULfdS0I8TChxok8Iuc6PSzF5m/hgjnEsclavdRKnNUUJqOFzxAUD8dJwRpfy
meOl8DITPue6+87AQxFs/ofcJw1xl8p8U7Lr+B/jN4G59fVLvKfQC8cf5s1ng4pymofFPaFlg6aj
g9Y+aX8ty7ak20DnngwWMED/srJNJV3XKN7oeh8mVy106u5WIOTMzE2v0dMLmlGr4VtpxHp1N2oP
FhyTUam30qVmvvP0OVPhp03875Wd1FZEYi+w9AZPeWSVUjENCCnSlQ/iIXQsPBPOtJ9fmiNjGmyW
gS1JSWl3Pk+m+X7XsUwGQuHgFnIjvI1BIGwNkVzyTwyq4cpcW8n03ssQhW5LLrd9va+Oy9HWQcGC
+v+C11sqc5dIousuBiRGK/q7V/aCJeAWjeajsUQvgplmTa/9I33NpihjtSH+y+50TckOy75EqZ1P
7h59YPFYbdtN/d8hdm3tuE+Jat/cUkWSetH/4rkrQmvY9rlJPmzx0eYmIC40JBrTS54ZICDQUqhg
9HCoaM6Vq/Bb3yTz2MAzxEGyFdbsukRyxETgddaZ8/DCuxWIp07JAJgJkU7I3gBz8JJvN0sa9NK+
M5KLnYluwPiv6xgnP6iMV42HO0Dk9CdKS518irpRtsB2wz6X28D7BHJxQ8Y+lT8X+xWFN9j/gbxp
A8azqrLICVPYXFZPuTua7Hw20pK5/LEq9kjPmcLg0l8nBqTFOV2Cd7OpLRqlW2hLfb5gYhVHE61p
rWwXUi9a7JfqjROoYTq8DmhLfplpiGww06Rkmmze1r3IIKfCR1GXGjMRv/bRmhp9XR1sVHbF8V3B
4FBmTfRmrrr+4TJ4gtZ+mT4QZFh6teV7pUhbi+OSTkt1I0sEPhtIcQlwQ8e22m3G/mByGxBcU+3f
UAbPjd9+35VGTBtTKK/5w5zoMeRZ4SeDOkprG4M2ciCPtWuMy3SL2xolH4H4tiRGk2+Tu63Ho5f8
FvIoKLVFZQ7jg+t/nJ+MYJBUIxbURkucBKJFNPoVTQouz4f/m5VV2ieO/F3MABu5OfKPph8Z3WZq
H520i5t+mOiJP4U67uuqSpWxBc2d65NNzHn8SDkk757AtGoW1aTbuE0G7YRFF1aq8r9XaagUgmEY
oc9Oy7SMUR6XnqxMq9qJw9xvpdp256N1ngMHYjsCN1NNGVJ35sgJs0wL0jRJw7hdyD7E+js/P403
eMauqQCWPR+/5Xvibh2ieZNqsGtZuutKWkxip9poVHCWdKzvgZppIwcL5EGO7wAmd7uetIYgfqR5
FJLUtPs6KwpwMlApSEZUU4CdVezWB+5TJdzNiaAo5IOHKqhAbMba53zLl3rwtbstAnmltCC6wC+w
7wMTIuu55BeEi0it8r6q3loQ3tx4sNt6HC+4wcJHduEJO+a5pALWzWyNsfhgdbY+KfmR8TZWiuHq
Wl34G2xE1Q79FTCTU5DMfCMXpkLMKkfTpXStvnZhRdtFfpWyP+wJkiwKxLI6+sDp8vD2hQn2NPi4
JiC1+aXwB8wiEV69WTG2fIpoZYQ+POMYI9N9sCtnA4+74IFJ1TixgBEXA1mpVGFQ/V3JnLN7iN8w
9hevBqYw6WuZZczyR2rpqFL0f2sVP0CS3XjTB6/i1vZHvDVt9VESKX9rRCxrB+3dgaiYLh9YGh9t
KYG9u2c8mnlev1sVQPcwJiq3I54XMXmxjcsK5SY47t/VVC1p8FkmyqDZUbf1CyegfytQ6v0CNrTP
n1ut3rQTpoQS3YCtJERZ06qpRXdwQUmHt/5gmXQ2+HQdeP6+W9VndHzTJF9pPJOFrT+qXLd1tHdI
5WV4i2Mx/1KtPkybaCwyNgeqnf7iUBLSevOAuHBTY0/PmBGOyA/CUN54BPaHLXoN//AqPz1/UlUG
m9Ukt67oOqBXP+GJP5XS9+9RkJGaOPZzO1i22etyE7dihsZGlYMNzb83O5v66MADknnLNxd6XRRe
4B6mOD1w+HJzod0L/ayNJg3K860MHMl3avpWL8PIOGp8foFua5egHpNiJjKDTzlUiLgBngNbI4rO
zcQC8fnNg59y7lgO15ZBl+2A9jpgZrA7dSCyFCpMjQVp+6Z2sYMSvPCscsr0FE2pFcZPewFvZWHl
Z/jsUHcANwnY1UDtEKE66Us0P52UMkAcd4IQEdrJVFjThSeqj9HVyDv1o96Vclg6qGougRqc9w1J
nbFV0h9vRq3EBvXW3ELmcCIb8S9HxYN0r/JJf6vpPirOsqUsOhAF4lg3UXgvf8v2DYKrlabzZq89
ETpOjzd+CF9t3NvqnUPR4X1QGeIr/uzLGj5SqnyOXX3ZBZKjSTdeHTT3vgcgjzXY9bwgNHkveaBh
urNE/W+rswG9DvoyUwTqN2bPRsmZIhTWB2T+Zn2lcdf67fZlScUUadqs2V37lFhHtJKPljbJYeaz
6gtojqpxf99ApkJk8CWonBDTl1rQRust1vr3HnowfO0z0VMKoV3SzkcGIln74pJeEXI12eNWm7Fa
A9rzOoaLHXtMbekkfaacE3pf1fgPo/sWvZnVM1Xr46HCMRHBVJL9+lPNbmMDn7BmjZJswZg++k8s
rdSEsTkh13aNgOAk00aW3apu74fUOAVADJzSf8rgGtUb60gkajCcmQ52bYFDCfR1e/L3iZTnQbx0
qSM0GdGwLkwV6UIT2SiE/vYZ8Qg+jT9qckXEqQoDV/GOAckVsQebtFJcO2rYHXJ1k3htFobiMl47
JRAM42fQ72V3KrpNVLjT/bcOhEW4D6zm1x0YN5AzxcfBJgD/xJ/O+6U7y7nGxb23HYTYvInlm9XO
+9glU8VPd+Ap2YV6De2bHz45DOTPDRJhYAS4bdbMFxKR7IavQw5n/6rrQS74d0PXROTV/UUrXxs4
Z2tnefjiYjc7e+CF+lugPdF6w75qNstunZsWE+9n9BWzqkGeJKKoqIWPEY8Y4Y+zadbAUcYfxdJs
PH/QkiG7rNre6oyZWyAMDtzlrK76DnWjN3NOTFDymv1spXB25IBjahZpq6ROaMK7QPaLdiv6ScZo
/bGWn0WLtUvSGm5FYHMmkR1X9sN9/7hluYq88XrKlTRZu6PdTC+LAkXAaSkMvgE+8QcNjMT2+lXe
g7Pu4t4DfMXUurssOJGQiSU3NjeL0cylavHr3iSzw8IY/W7O/xasnO5JwflPrScoIgrWL6rMWzyt
r0wm8LHv7nXYB5XErKLSaestxUtXw/ID/0K5Vm+iQSdp4yU7iLcCNEWCo1fDuNHnYCeV5bEolMUL
i810lI3DcfwDhOyXAQPyl3h5/E008xPGERDi9uJgAtQkxAYtJnzoq3wukIxjX5G+aaNhh5mljVuz
jXw4E2DYXPGs7z3bQyJWyKV1y10e1QEkzl99tghYFtx7YOgwAyx4CR+20FzRTSRDxdAaDluyFQw4
2hfNgtoa0jXD9+4WLB61NP+wGEs9ou+KXj3h+JP02WEdkwJNFHOnc6bt09Pk9fYysa0sBxYwjZVa
wWNx1vmPcDWbMnH78+gyqKoGxoUH7EUOKJ/uaoZ8Lf+VuxvkrcfGpR6gbTYYMip8FFzOCNfDmMnm
D+yqw9ByGj4y+tr5CPwS+Ut/n3p6oFTbSsXWPye4xZ1X/Y09MoTMrZx1wmBPoZ0s8HimIhxTa/Rr
lI+0ATULTqe7JQcf/w5G3cYkoAH9YiJ1Yhpeb+R7mZcHE6WVLT7CMyM7uXzXP1eYGiCxTZYTp/gE
StqvQTwRE3HQ/tthpgWn8brNfVoeuWqOo7w7fg+9V1Q6yClkoGphmkb/vKh7YlQGd1LsGGf3BKMQ
XLokEtYMnJIj4kKX6FMUzbxHwuJDwlrXeZ+TsAKj0W8w/+xVvDgJFGFxn1Ck98CeZBgw8QCjd2e2
kEs5HBmizmczpMruWs2A8SnUpFXGqTJZkHaAsUVmzucTkWMGnBx87X729Flrk1E2mDV11DEXbmd8
8ayP4ry0ZqdkAaYbhhp0NnUIXnaSd4yp+GK/dUNLzGe7Ha0VXaoOHCKGhWLjcYK7kCBF5uh5Dury
oTwmd+Z4Jl6jl+9acW616MBBiXaMYqSEZP9grEGWLmB257Lts1zyQbXZzVUWupl77EgsgVNariH5
713/FDVWIW6Sgddb6Cb49WDyXeQ0PKk3pBHKzfrgUH/YVUGx8yJCkkx/u6dz/TG9A209vajHJFO0
FH50gq1Q6BSduvuylu/Zr0Kzs5YNBXJrmQZUrU0MOYEljzbdtBOk/lJGZCW6DnPCFY5MhAUUCse0
dPs1CmCFXISBQMiz9TVOI9ketiMo8eolghaumRPl+NDMxHPXMq86sFjH3weAVGVeUGBbnNxOKhps
ICQzElU6TSu0h+MNaduoj27cLdJGLHQGYT1DPZ5vD0usvBfSFzsDq7bRymR6Z/YiEF9nJ7TkvgyZ
VLUcEdI3snAQ6urnLyo7QzB9EOJqVwaZTqXUx76mD1PyKAh5Mat7KV3OhWa27+8md7BO+utP6DuX
0QxK4RdLujyzRLLj6sZhHi53dgX8KI4CLAJYt53eGZvJ2Y4N4/E852KTQ8/gWUuilzot1UtAkC/3
AqnGkObiRPNy9I+X+PWZmCCAK7uXjvASXTKYlamtuL55+ftDyeJiu0yYFCVS9wIua/ajp9uK3wmh
27TQWmZdlyISRNDRZm93oH2rrhjcJeOuLJnrw6ILeqrWean34rSEZVjAMlbRZuDHbqTbXg9OLn3r
RZ7/yWHe33GQ55KXFF9rcBBj28ZqV84M7t9I1SHVpvSMti41JbHPKmJ7KLS271OFNYnuaO0rT9sN
yi0N20zsGrCbaoGaoiSiS0S950lWf0gbl5cbLANTivPwLF2t+c4BDMGXd13Y1273xtfCfUtJRZCl
U+h1R4LSm73IaFlralyIk7/xn6oYxqG3F9MFyKcwexrBueScqBcnXDxQu+qifwxv4FOfL7Go+s5H
idL1b7b3KIKrb5ZWi7QbYox+8K8No50jF5FTHtcbrrxWPxEMva8lQd+8GV9Q2gPot8TxbEh780it
q1rKHWWsf90B2J+XgCu3MNudSwzl7qOEVhRdb9PMFymSaX3JIKXBHMAp9QklSbLvzbp34LH7TKlJ
xLK9ytbVysdnhx+KHY0ZFpXzCwpG2A9ZQmSOhnHwMoCx1N+ANrV/2FTMvWHGb7R43aLS65MWFB5C
aMkr18S5tnnF/2m7fmF/Wuyb/wdBtHFA+9VZDkIX7o4FZ8An2A2DgjdxrKQQzZPOHIa2DUS2ZwXw
2r5Wvyq9RLyJl+y0PBK6cy4nJJR65w096CGHllced+OJ7ZSK1PY7Q/6Kxb+bHv/YYVMg84Pw02+Q
JqT6/N1YrOVx/M8yVDHQHRlrP7Zw4W48LrricT2iior0pUB3fThlsWB7E4EPPlbxpSjo/al90D/P
tAag+Pd85YXEjwZkJYZN7niBVpP9//wd8C34nKdXOfplm7m8Z8YGeX8ASW0W+PPiaAZKATv2ovoP
JLFhSb3QVsmCsXd5ForNpT0/Bx6oFrASwGN/227sJPOMJI0EGv+W6SCEke52/XF1YRvWAVUIwniG
Q4Y+acqzBoV1TwnXeR6J8R/yge/i8e1tuZlfgzGVNrTkJL59/v7Gkx6cqN13rkM+f4HoMMYD+4Ql
yNxurlbdFKB+F9M+VPpXPurAvWuDEd6Vu9MvMA1HJmZioU9Pz74zIHD3Td3ofZ+hZWJSjQCu21i2
5nkPj9E0gcdKl372H2Y21/Af49nKZ48DFqZ3zzZ2CACZ0GYq9IKoSqh4g5wc3y219BX0MbYJnAlu
d1ztIissc0Zxce84XsqsonTdO97DXkYsMvKq/ceA/qwPw6jr+WJceOrt4PdAo4SNaLYcYLwch1Gm
n1gO4MRWEaSHFvafAzOjDkKiTL7+EIdlfSk74Y4GByZkPAlkyppQ+CoMVXM/aoRhh9jh+4Gw8fA6
Z9KTpGdbTHr36cxLVQmItr0MIgldzWKkfZF33yG4q08/kG3APubHD3VD0U3Xs0+cKIwFPn/iHdYB
8aPVpKsbxvbstlv6IrxoDjERG2rBh7UJoq+3HLjE0ZW80i/gGVafGw2HbrTMK0dy0FSeIVZdC7Ln
O+50/zQVQhYTuBUfnjgA92NjJmZwCaDmZXW1b37xdgX940SwPP0e/DJj+bmonIETC6nnzUhySD3q
FxhnoxPjIlkieUVt5eeVMmuYVChpTC6vikJ1IFq4xZCfeQmmIZL+a5bP+r/LpVszKrId3RZ7DnvH
2jp1QbpHqldbR1zIs0Q0TrtgklUBtJsUoxNLgTt/1SFemzM9gUAunTqhIZlwFGq9eYRWq2YcOs7k
iSsdBT52akEVlbTCmfFWLvNH8gmZI6aZvChI9vCmtT8B4pZKpO/8bWdSDibeqt75dPNQrrFPfYL2
z3LbKqj3GK/6L+njRscsilCmdroTlOuRLlL4TrVaT0CmbO3Jm2hB9YuYj9FJoPZEaNesm5FsbWzs
6N+o0T6AMNsakguAZZCx/J4g704IuF4z1cdRj1N0jNS99YFwwcrad3kie41CVQq6pRRsxdQM4dNL
+f4P7DLF5SsjPtlzMqShr0cGM9dsa9cezxGu5EUL3Sz+rNnzIupT/k2VC/QmqwPFE/pNIvSNGXtn
G1jiKt3UZEZ2q2+fv0074HgHdBVW2Iz487WPTkl6YTGMIAVL1Nf4FHP8S/n5pVG6BwIF5JLfq2S8
0BK0DHAffhzBED8xSCtWvxOxs1tR1HIHMKC8RGWHsf3ayVkrlvI3/1b9BZnZDG5CTzolKBfXh4FP
egZxqGDRkRIhIxf/s3tGaLfMpzeEcr3ZrldOWzh5f5VlPUVIwtbjnbA7Q13W6GtE8NmbEMpT/mmb
xjJ4RCSJ+hWbfGhdUVLBEo8S4Ob7nFuTqmFSMoGsRMxd4XHXt+4r2CJmK+QwLzjQbJ4S6iiPpzl0
bM3wtBFTdZitiL6Ce6eatDkS2ynoZpKIpxZSxSTrhyT5Q63b6zRR/nOAhzVHmP2HJR4bd/xeuuCd
sK7PlzR2Ntjc0DYseM94D+dyL4OW56qreuRxz+65WvyzDe8awEWP9ehUtzuqMGqJCOwDRlcAb8IC
3J6YWctMxNwE9Q28BUEjNGFxCXP1Xe9ZRmgbmwrsTIctuifvuoxcDSHEaCS39Yr+mbLK38U8F7kY
tilmzYYIQL76y8eJRKLRIo6VqmalEQJK7AX/1afhwOjRcMYl6+HichEfd578qmgPI5F70M5GEYGY
UHMl6Rn9tRwufej9MNRbt7d/X12kGh378oy+kbMk5hWMNkiYx6dd9VMTpojZx8KeMp20P+qccM90
W4WSDtCeFctgIT3Kb4eFviiXZ0I9/YUFNp5cvo37fzAqdwgRtyJi6jUFjEReVxwFZIIuHVnetnCj
GRf+QCXImtFE1t8BuOdoukM/bN69b9HuEkzs6gsNjQfhxu12v53iXJOT+QFcKlFvD+Da99u644Pa
vpXfzRZf40YOjj6UcqVI6r2phqsCxL2PqvjQjsYjCfTfSkWEXnf49yFLBQuKmZ3fNE/Y5cjZm+uR
KFwUSQyGe0z9ik5hCkftajPwBYoB1KB7vD2hJi/5I/0/NZUrgdGMdvTGMVjknAF3RqgtiJvnOaUk
rDbf/RIBI0NYRKdr+aOas+EB6Km1Q3FJZXfeM8QaP8amE7kiKSccNLPIvF/TbHWwMPuhwF6stfsK
gBdFSHC6cJTnKNLJfI+oyaPwOq3Dn8joWLjsMP8ITNoTPsCEbWucT+63HMfKwBuZHYIQ2XV5OzOR
Nayy1ep+/a0v4zFpooaVkzjoamA5JbBn6VqWm+4smkuuOp0cdFC76imMx188ejAona9FfqKLkZK1
+wk+a0G9jWzGdrHEGHN3hwy9Ks3hBVa0nk0ad+F5FayCRtNYjwWhJIhs2PgyMag9cdVdZaxbAFnm
9J6Elzlkd0fZgn3g2sTz1Cjg7qRyW1T43XtMdzHUidFNkVqwPZrMLg7/MAJRaBvBRE1dxB6QBbJ5
6UiqbDvZdsAVTyZJb80wEjaw9HDFxmQ/qrHni589CvPYFhqpTaU1V0RrmoNoqAlGv3NyJ3RufX53
o9/28KHVH93lSXXJ03hVgsR5kBTOfFEFu5276jJGQxpYyhTfvf5FnvfD1HKpitXsNQeDVQmoB7O/
QpV7rg5zoqZWv1AP5l6nVu2w6FyAaYTOr6AQpgD9F6Aa85N57PnXS6eG191N2pnWtgNys+04ysJQ
cREqVcWwYBEv/2n7m5GEWMeqoTiqPYOxNk9UyULiACMljn6xqTMVnyvKATAufZ9hkMe64d4iCKfx
wvkqydWObgspRZJhxPD/gq+x1ERJAyM9brL/jqjlJQ+EbURn/iBucJi/NYjVXYGY0iWErm/OsTAe
JxQlQnwKV0f6zwzrzooMQOuQbg3vKtz1Hl6bFS7VikxNpa93HWt3Md4D9x/A1EzaGQ20dGsSDODk
/Cl6RZbDFOA/xp9UCcvNoAMduy22/AXY2AJWDnlYPL+scY76JbIJ0JzdGbdwAjpxeTTnba6j4IeJ
yKIqPbnQtd8/DUAOMNS4PEIyNJDe4D/dH/RBNGyZgSEmwQT3hvbeCJf+UTuSdRlKcNxr8zqoM3L5
vMCcq99MYH62m6jQRA2iU/iiwoLUvCEdZWJJCd7HjYsXNRdoyUHSQGOyDJpNvQHdpbbd30MxPAia
DxMay2BGbeHPGU/3SPu3oS1YfZ5c8xLtR3238dL3VR1a/iuw3IezVwS4k3NWtu0SKoyo0yOMYbRD
Gt33y2LFDChNgpIz46N79XtqT272uyXJw9HOjuQtY6DoyrH5FJyA5JqpPtiXamqyfSQ+oLcF1NLY
K0sav7fnIJBNuc1ypvMmxMJ5seqiJTrqKw8TciSo6j9aUbwnYs8p9dyp1hHSExPNbtPjXMji85QM
OZqGKdIhW1BZ1cDYgMNHGZZRSxIFHZ5WELRJMWBW+GpDJErjmCfetxJG2AwaodKRGcdsDLkJoce/
LN3j16DIyHfWPFcb7t3WEyRxvpocht60vopbe0WjcfLb05iuu+41nlkgfbW6kwVqp1k9JnJXY4Ns
NcPzdNSxhjEVZzE71GiAQhfAXIYg91VFKEoemt/ErZ7dYWpH5DuwFzqET3H4Tbuf89guCfQjm2t3
QpJ6R7ZYFii6Li2+9o1vQj7ZVWJzjwtqbdl/2oVDMT2pcAQDqsWw/VD1vLnpuOwHKnoDV4xqFnaU
Wn0VdznR2UupAFf3SWyBHlmdUUh4FfhGXSEdfSpNAyR3W4YQiYGtpz3PAnwrNdCn2pxzJG1w4p3z
kVTnFIXw9LI94XU5oW0+b73aTIn4Mo9CGF6geRdc6eJTL6moW4cIEYgNEKIqWzQbf3sy/C66U1Ne
s5ArGVcymrRX2/dkDv66Qmr0HMu1raELID/zI5ZpHIAzaRZI2af9PBcj2qF65zKc97FbBpGZ2yYx
RSK0f9saRGmI1h6BjEuHh2d1ic92er8P0VSPdnIBPNNCb9SlzWhbvJ6Kjh99APpslvYrDQflfTyo
duyva/PWE9FMjpy3GlCRxUexEHCQQZ4Fx8FFWld348TMiz6KmmelP3i65cww4DMW5ld2N2+U3r8W
s0pr2dEH41uO/GKErqSVTyES5Cfw80hVM5xbW85KwOymjNsQAAH3B2B+No/Tce776xGM9oWMJJ97
horkcZXNnWynMt7Wm6OXoCVoEwmLe/KvnEWXOEY+0c+vR+DXcwoY1yxfEpnQ1FFYyyvFVx1LPngz
I8zJVfPyDxoxxPQRsaEfnSRao2RMsJZgPPU1BV3aj8f43EaVWpjBuIe5YbFezW3YguNmQWBbRWhA
B/7wT05bY6UhJraz6IgxoOevDq8nIAlEx3O2Ka0D6OqqesEyjgjhO5HfX0H1g3VgdWtyN/H+Eqwl
Vn0oN4boCKtm8Jpe++V/dihhoV0/QoEBciwoWMi5K03BN0deYhpO9NEqWy00BphY/YkSSGBczvIM
7cdmRdfSLA+VaoIiSE4ZLLEg9Cr1eTbyi79spnWmdqZSSK/LO7K10QubFrXxJzKMLy+/LrhRRCEn
nvuNheUuUEKvCSt/Lqy3IfupWOo3bGrG3/vZXOJc7NhfC7tG09bIUVxVAFfMwEhE/B4PrUeqlexb
HqvadPp3zjBJQoAP2PUzAuVd+0jUNBSd+k/O4WEL0lGbt/3kBDPm+HRsnI2UedXM9VZUmLjUOZju
4HjZ84T+7+4cHuXbqH/FXbozINORFeoaLaBtDePR5DUdPeZG8boVVcmYCaUBmhEhT7HzrE2CImbh
n8syNjYlikId7klOxgnWECrzVP6/RE60JPbb4XzCsXbk8prYWhXHezH47bNC2+hZnZ8qiPCfvgvV
D+KpDnreO9jp5w9Nw55kow3Sz0Kkzvjoi7yCrW5YSeiWbOuA9eR8zsTVQ6l816aYt0X+dfzSFYAD
XZ+iVczLXoajZgaX+IPmA4WuHISpErMEM/PKMIUVQVixQkY7Zx7xSxvY7UuUr8i4tCfhVhTtyhlD
h8bkv4MzEn64whC6wuKrYivzoW4Mmv5cJewPATgZOJMDx4dSEvrgFXN1aINtH8PqAIhiPlF0ErHi
23jRZe7RH6HaTaPdorCNAQlO60UlYIFl0POQeUKXVsKqkt3auXudY5x85pm7WgXol2MZV86DZPk0
pJf9Dbg1lLL4Aj6ijen6GgBKid0D8n4yFYvkX0+z9zx0uYCegdg+zuMjF1s+yOhj492e8mYpcWLx
VUNqkxo+47SctuFOCO921tPZqgjZZasUJFxDOMuNFv9pjCpNLQEvf1DJaixs08d5mzN5I0cIzHiZ
7jSyQzMV1h9SEoNR2f4WxZwStvamppzgmNm3XvvgFC2qMAQu4TU/O8FmHhL34ssM/X8sfI/dBEY+
+TEGydJAAaRPSGK5JfCiyjufYX7aiPhF3RzBL5Jguz8YLB0/jLUrNwswWn8HUaABPc9GPs/k1HhY
7pYRjlz3Pxp8C8QUisQf8QN+oWaAoyUEF7JjZNu4eIqB5NqBxhO0mqpOvnNEEAgMwQ+0fdDTOe2p
i1K79bduXK1nsGfJKjUpw325qD0m0dAl7b7jkYj1ZCDBj8o500YfFPURmc1E3oDPJ5CGsSNpZxDq
bX4+NgrdM/7xGBlBGCzqd6IzSP/OZJeJHufHIO3aGCSHx2q3Q0hJwMo++e7Ml1u6KnB02ayaOaGc
PvKssKTTIBIZUTOe9abhUKHquC/zukRtQaKWRfvXcoaQqqGjboMH3EmKVqd2gXyDvyKSbZQAwtC4
zPQg+biDERye80h/+EA6RoNBrBZlnX17BAYxiwfAZCsDD4BJV57etpcohGiI0PdQX5DmAgH76Rrm
agJRiBDHCIpjQ4UkQJuwca2SpgDo/M08gJdtEolaJ9w+7qz5f1lchj7G4cV5CfPzvLchcCnMZx/p
4YPsz0z5e6uzYTAYFFnHUWu0Yp/fD8f1ixzNVZBrACoPRsXq6OWZco+Sr4dJHF2cXNwHIKmsvxdV
5nzLDlqALy7uw1NbOlF8PW2oFd/+4u2HiunJigJaIg+t/uYQz2R0Xxe/Kj+Do2OSKcCGxU0AytuT
pRv4TkJgpiKF9hwdHaaimCGufup0e9IA5q5ncbwrXsQOA01eMPrSihNS4Q5r0dHMn+/6k0TIpwb+
DFdg/Gu29x29rfekXUvMyNJ7ATTFoky3bWibdq1PV/491xI9ZbgWCXg6JJDH6Hy55ryJ3WDUv+4y
Xg/MjyxtQ/fWTXTkcwrPbvRhCRvMoZ5yHrR6cJ8llyM44T4FU7g9NzesMhQPP9u3XoaqhOYhdzQl
mrvoXh0Gz7VtLlil309rWNWTlaN8DTx04wFtjvd62dYRKk7dcBz6F+4ISkzVopeMWLFYI8qaDsE1
iZJdHnj2Jm6g0Vc0lyZIW6k72mGtbJToDgXeh9Tx2ihu7gVIprU5hSowuOriUYTQz4YrK4BcJikZ
50kaTdBc31uBfy60tXbLgwkJIewZtZqUAUx8dsQxNvQ4wrIsHwoHdqSiVMnGBNnsOq5V/eyYQDSR
LVi54zGpU4/vBCXzVCR4jqgeYARITAe+w2MgmLNX8bhdTzyphRWD/VQEVbD7DvFLNUOhGvPBTEO2
wLACjdJLY8BOd5wwLN0wwyS2PefAWzsoxRfc8V+k2rFas6Y3omRy0Z826Is/frmAfCp6lWj4I8mH
DINswb1S1fhHtnb7HSMEh52y3OfJgoIE7qXiD4+ZoM7w4tmLrwkgKS/TI4tuAxfhkla3R0vJrmFA
8FybGe0cAKQNSlZp//wu+5cC1QxSX9Vyl6cIv5uF3/UlBD6ERPCJQxGmCoHtJgPCJrYxI/LRqRWO
QsYaL1sAXGA8VwaOcWHDNXK1wy6ADTK4IUS5Vm1rdylu1zh1f6RiB+ZFPBtF2rNauz2bhjUV+nMC
CnXN3Wr3wO65GmYep8QDzn8ICtIYI1OCfy81o9ZTuu01/aH9ModU10zjhaBpXk09WYkyNE8Ks1yn
EGDiUcaXwxNKHu+9dh2JZ0Eprb8K3FhplPtOdvfWH5nWGiWKhfL3yZO0Tp6A6lgIhni65d+6+CX2
G/1T3aMipJOluDV85ZRg8LCDXtlm6tLurn5hwhUDCOeNdQ0ILJpS7J4k+1GgJwe8IdfJlReCMxIo
cUEZcdQeqCLKOOM/mykwWCY43q0+vyrwfFnxkj3g6z4CjJE6xMZKkCvPHUP4X7PBGhDT9j8Lsqk/
zX2Ygbrxszvf6RLmbt5JIgJt0TDLZ0AGUMgBVu8Vlr0gasY1kuGFlmC16DcCPQ2SfIFnEAcah8FB
Km9XO5oT1qhTHnhW63gmEIN23WhQlxwPcelvqMl6s5jP4HNSW26RM6vzN85sQSBMf2wG3XVzL9NB
D6Hat2L+J6ejyMauCO4IyJIaHtTSygtfbcETWiOShexTqsS8ffs/YIaaLhKlcihBU8tfswkSMu3m
f9BWvIjCxEEQveVRw34+7MQNVxNHi9goEv326HcEsbPo6eyUFhJxo3XI7ib2hFcTBtY450bpE6pw
VAX8ZsxOKrIta/f6qaAhqsFt/PfXhNIrQxzng+tCzyTAdrLxEaO6znZ+9fiVniEXLwai2w6/r3k/
hGorkqS7wsVf+CC0I7zD4Eu7rawWiBdcvu8QHEuhwEChxcw34eVrpBrLx2sO0YpjmnHT/RGFiGFc
agyXLZSEADM9kBB4BW289idM1kYDpAsK4kqp72X0yxjAwVaBFVXnwXfN6OlTMpfxanTILKl7Q2Ll
WrsEO6Tz6FTBgDGpxYZxL0pCej9Sl6gfiUpAKhtoIB5mjG1maySoPq6x8sqKQzUU6WUyjr99Ohc0
JFm3z3+qafwP1b1vJLnAXRC1LJoJciCT4SoQZ4vu+YoUDWS5mUW4kZfAGVEHBHxB+VHarGfqZDNU
azG8y1i2d4SFiL7w2/aY1mZZm+4jFCzY2VZzBzwa7j7HfLO9B13rKLXtc6NMgnFzMt2fjevXhVSI
PPXdIuQo69eCAdPXNgFaPAfHbrFxj1K5GtvepF24rj1jO11KGB5DPrexlQa5j5YOfq0yg0qZBRe7
JfTNv6KGKz9xODdpwYx2Ah/bYb/G0SRYMgJYfKwSgMwKG259Of95qb74QnSOnPjBjq3bGtGDtT+o
qb+k1CoV0B0y0XbVRgNdX9ujAAPAaMf82dvD/c3Ym3g7LaNM1Q7l87R3+KAJNoJf8SQcBNdwAE2P
IQCaLoxFOiTFnvgJ5WPV0NbOOq8CpfqmyEVrMafMSYoVGIiEaIatgYA71QGLzhMYaJLPXVvCP9z7
CaL5aMkJ0RlNQvRENOuTa39D8qdBr6ig0xjf1DlqCEmtjjVmgavEkSCxx0zC51vPBYs+S8vqSndT
yi31nGswr8BR3Yf0FvdPXxm+//z0TXosAHFTb+HM0UU9b+6orggEZK598vMFbxvER7KdUhQa/GHL
vCFPeUmO2G6MKHwj1l6pJGt1ohV7dh3dvVl6dF7eIRlpkvRYMkttuYxA7bWewnp2bQ38Tmnk9cgD
aaJ0SR7I21jH0ys2YauzTyj25xL0kERfuwQX2ICpF9yX/BJJNPKjnYk6QdMH6p1dq23n2Yj1Xz7k
B3N84iwXSzZpTNV2NbiRLWTg4ho3kExW/nKiFCj9bBWXrlUZf+G6tKxR4Ats/UlfA6QHLX1r691m
eyIfp4kGv7JxnPHph9c7Vg1mn8kQWsWD+4rn0x0ubTaTyBr4TFnrSWqpZpYLtFAFRXWDEnsktJAG
cxMV+/FpQM9IkFV7upa8rKotdK0e3SGwd1+N+Z+hEN4khPzn1vgEgV4oYMt/XJoWQflNJB18ET4f
Z/0WyCW5n3hoWo0MZPzb4E4srYvCSS0RwikYfZAUFM7E0mp2VpF68g/U8HMVRzORbvRb6ECBfPtY
1EJFLSLY3TCugidfgPF+C6Zy+t4p/AwGyJ/tcdXfOr/ceQRyaYwG0EIEPwukxWYI1zRwLruYaljx
3trp7c6wggdJjK7IORHhk8aXnt1ANKK2bQpMgjo4iZT0eM8arqEbF5YFcAXxVb1u7Me91GnAHi5q
7ybU9pgoSD8AiG9O3vGX0uKknQzKfJVzYiqktpEFg04CZjoA5kAotI6HME7f0QoOkY54N+Fps3aG
zzO4Zyx8QyyLCVP0rl1ho3TK/HQbPa07GdObLRSe+fizWWh4KBEJw5nGLIzpjJAkqSH0hVJ0MigN
TH650I5TGuOsc4wZl71sAk26FZPhaIEe8KTAuXZfSxTOfzSnJrcGk7Gyj+ggbXe4PlSnLTkZP0Ke
hWgfaQIV4DJcKH9JVfwHmcWlJGQCCgtrZpC97NOV5bt9v/YIz2V82jR9qyQAVZGU7UOI69rD+pZB
+N9kR/19BHD60udcevXBl8r5juFrLHAr7kAi41M+PLML7mEvGdA61uNc5NNp0QbpQBvreg4mlAxi
ovCiNj9lFzjKyxtTS7xUYcjoiTGmQRavD41suprkcEFKs6flNcCutJmseokgUnqZJCVijmK61Ni4
RkdJ8D53dqTgrjGFSQWYMJUqqNUWbGIaIH8/saBPBrxWljO9UPEg5KHkZGirg65PL6mzfuD2r4bE
gppYdO9xex4BT8BRjMASXIwiztiU60/0voDkgg97nxlFf3PQ0/UqWiyBm69dVgUVweJy5FTZDsKH
riB9IZv9UceghcZ6n5qJD8J0efHX+QF84FICLVpc1Zd0zKGGbSHwfbZ8S6SMP2gEK7zoPd5fmsOo
X/y+oaPXmWDWvuKT1SmtP2vjYFSo7R8wV2B5m60fLrPQkYbF4CWJCybwKeGL7twa3LG1GgK2a/GL
zUaM9BWdzQtPRhvzACkE1Ys/OrBQhUVZpTqFAV6q2ccjCYNuE+MSRJniYknN7i5BoMDkPkyyN431
8MBrMvTz6wDQvnUhllsMT9PzleBa2OzOPkeM7NQJbi6+a+jRB/Y5dLU7stQ/v4uueAFJvkf3ug/V
fnBJoDhKktrPFP9qio++MeVW/ev51yOfPS8Wu0faXN1ECYttKc+/dZvNBOCQMm9fqFSC+z/cIi66
TVvgoCcR/NrDMUtkn0Bp7n5B4+t4+MTMiQFZQOfOcewNxwspAXPi59t3f/BU4PBrBN3PWiF+WwCP
Jgd667VXhE7h67V74z0BWTD43WUtcljwiECAhcyrnS3nPBI1Rj4anhOKDU7jcebtdOQLyaUUmFxd
nq6LFJqGtxI6/RIBofx7lFolju1Y3DIkP/JYe/Dd7JpEh7eZYccFIFo41VRjOmVAMCNBre1hLVS5
YbG7q6UpJv8Z2yziVI/bL6tRmJ2llZnANk3WDJz/Sl1uB8/92y0P71Zvgjfd/3dCtVeNoHF6GP4g
lIcE9WYwA0RvU/V9LeL/kcGtK0hdGZj6OK+LIrO93US5AGC23sHkBWls/KSNMtvH8+e0PNfXnA5A
qQVgQbaKhkI2wN+yKgxJnYZXFR5rJHPCJnJfxgzZvRU7Vg3XQAQwIxdpc33ZIzdKWClC3eInI2TO
OT8lWeGCSsfDRlLOAK76o+tXzZuItyejSyqGbcoU2IIepvnlHD8url1lhq5S0R4SAxO7SE8/oSO0
gmnG/0rO4EbWuVx2nYsBPh+VII59UeqMniSHyhEKp3fed3CBv5jQXIQNObWt0woLvWOpHA3Xw4HM
EuBmaaCCLxsA6Hm+nkD82sFDtyYHhkaKYIb9nD4A+hGJ89PCnAt6ZJWLYi9V+q+ageyITsAJ3nx2
RnGNuKDXVJRHpN8VQCXhUgSinGwaqtzlCKYv6IOOAO4kqeRd3mMeDvmx34M6XXc2+LUaHQWzHvOU
NmKyyz+KhT7rW39VWYhsznKMuMzqWO9kizMjJAusPGw+DeBAev++ZDDLmDVC7FMc834g51RYIZAV
ae1yi090u9pSTfuhNjxvXnYJVbkYU2Pgm92QLSW9+aXs0GFuvXIU2tVf9Yt4jzM1SgfDUgIfscn/
sXee6cvmgJ1oBLBByNLcpuJx+ipZ+jKqIwCMN1WXSWwItbUpc/Fw8+Sa79unkxVDDSD+fGiY/kMA
x3BIdpvdQhwK2CJJ04kX7pIhm65cG/qrdzpAJ36OkFZcfO2V33MV2Q4mW17Rmxa3NQ2oIagQISMx
zhMD2F5jG/2YH7Fg+zZosjPU5sSqQLUoDXwMTQzLgXn+OWHOrqL3SLdFoNGS0Ab5CuPD6rP7h3mj
T/IhVugGGGtQaC0954yzL6KqLnc4sHMTwBK4lrc5G6StUoEFprQabV8yMEb+qgJstoygbKYygp03
dAfhVmgkHo25Qj85MEChmBeYSY7vsUO990qkra4HC9B9UFzrGUqZS0shsjx0LQqH0WQfNESwa2WA
JNWVgeX1MxErL+awhjTlxOdthUC6lOzp+0eHKbm3oCC/dV8vwSTT1p5IVPg7iIOvBrq2kefGHYL7
NdikX8Spuqiz0ayTcxtFgSAOeYFiUrxWXVaLMP2k/bdiBj6U/zeTruLUtIyC7wcN1mF9GW1Zy032
WWA7lSQR8dmVF2eQhVtNhICX6nTSC+upzcZkCanlvJ5pUC39/434bcnkmNvN1Nqmb5/mwDFkR4U4
lOThvcmVSP2IONWy5FMiLBU+LX1j4gSAZbgD52LHudECOOYg81EOkzW697XFedKUKJLXYbFfvdFI
3ZxJp9g4KBR9a7Csu7sPEfDWyk5qiJSXqHv3Kp0//VcA9U/pKpNj/mlBfxdTfT/jLhjkvJQP6I5I
RK+8RuCwVhBaiAfMY98XqSnZSssX8A9TxWwhikZ/jQIlu5vADPK3WQzBydi0mV2hlPGXU3l/lnXF
iNkN8SKRJD34wiii+XVMbbXOZwUih90VSnx7a7/C4BuXhxjsOur9ZekDtxM3w+HW/BASnyfUxpAg
pnYX8qFGwhloKKuqMZDcd7pbMk10ywmRlrWsFh+fkk4WHV21Bzx0xRHWoXCfzz/vGN3ubwKAwitt
hwdBVf7Us9GySAxvIisqBLQw7ElWMkm2DhEn/3ZflqXIhDM95yIumoZpawwAtKpeSqECqxjOnTUd
ADxDHMqVswXfgsL0CFR+is5F5rbvodiBN0HH9m4LnaS4w3tW+o0lwxSfrZbmfM2nSKAxkux5ZBzm
foOgb7dyh01gdgY1sIFIhCVxf7MATTXlDIpEKIRY/KEoOlpbfM8ndIxXYiNVOGpe5RYHLg+iTBPQ
BQ2nuctWhjp9R54menBgP+4Op4Q8cHhIfD2KNdA1ljB8uv/vmNM8qzeauY9U4oYFOQoNxX8/RIS1
N9miIgl4UTUP/b/rNK67c6rx8gbzvv02o8O2blTlv1KS/UzcqQyitiukLXYpsFt9RP1n9zYUPSw6
vN0k/hdM4uvCmB6KRiEFXwLcvj2g9TNkctkHGqxP6010tNIKiHZ7jHABswxzOMNEqndCSpdOzVxB
IWD+JEO4C2yEiVaUqLuBJjT6sfhFwL8JG+R1XptOV6vlSGLZaAVMyWj/PX5b/pzJi6jbOArrO8bq
c6qya7oQN499gQK0Pd3UefJHQen2Hdc1kVYL0UpwOp1BceFAJ2Iq8stKcVeMwhLC18+OK4uYOj/n
1Eq1P2PNM7RKn3io7gOjH64XrgceT8qI8a/8OxX0VE+zi57lQzTsTOLOZILZaPTtxz4TzRMcD67N
CzFvpqqx3QyOedtKNrmGPwlVh8em5HBKyr6t31Mx+mW7HmGCIKjFlsaueDlZQyvpvhJcANwNwWe6
Wf9EEEElrw92iH83IaCq8+mCe/New+gM/CJbNAqboDo78KggZ0xc8F63HhdhYY19Z2xkJUZ2YApD
C2oUd7FHC5CBKBvTOU9tXADFYy/njcR3vSrom5rFsUFCUz+h6xpSDManX2vs1eix7IVtkPQazgOl
SCWmc77ZfhbcRWxReKHDQkAFXwfDewbPrLuZAMWt7Jz5OcVluT7v9pXk2VpI/sjCtkyqySvNCrzb
CFLxwpBe/oFJUIUIH31v7AgXg7EE7TMu204wecR0UkSPuXvJU/4u7jCVUdUdaWNYIYs0PDmYCC1J
2FCC0K6VSgdEvKiQJbgx0sjbziLTeRJWmvgvKC6wFnKziNi1c/7ZBxTVHMHa+rws581NrLWYpZ7X
LKXqHJhCUV2TydF8CQyET4rxzDFW8dv/7Sx7o8vHjQb97WhiM3DOh8YhhtCgJX7SqZ2f3pT9xAP2
i0UEIXtAxZGLYns9Dmx4j1B5WrGiuwjJEwDVMfwTYR9gcx08T6RpcgK/s5+sc7UKfChHnuuRmihG
jgm1L2xJk6B0K7bi0GedWUX9Eyhwr9Rj76R37VM9iG9oBLGNTPAHcIT7rj6gZHPLrDzkdCRHJTPM
GkY4snCftwFLYuuwnRYkWNgFo1aGwVhZkB4KfGzyhIEPbqwKYA1h//F/IGygBZPmgOVEJJIpdF+3
6kIcE+AIrvTr4gKSzA+Q8FBdMC6ajWPa6aQa7/zgCaiiXQOYNPrjVN0EfGu4LUstG6EDY2Bm+fNI
RUE5Wkxfksn5ThzcTc8V4PApv/OOJSM/X3nSNylf96FQzYbUW5QtOq5PwfNiViD028LV5EqgcR6m
Oqji3kQwrzOvAEtWmxUZ939T8Pw0BKR1DEHssWP1GuzHbc9VEPsIISdHddoa70Qn6c6SGCSLOdiq
SRyIbM/4O4vsmqjmNuKgkOV8Q9qAr447bq/rGUBEtACYmP3ympJVJXO9Xy40AkcQU32nkGekYHop
2WcsqWIG/5gZo18ypwMlJG7LflDAWZzGXXe1vBL+5T+SN0Nm2fp7/fd46adHZE4fIytFsMvpdsdc
Fx/p7lrus+9DuR8HT1brZs3t9CTXZPEsqT3FghJ0vdiLiYDpvd1MV2UXUZsoumiGmOf5d0OlzVzF
4z1+Uz4uuNzx3N+zIpdSMr6twsiVwg5p7eno56RcAbO5oNdKAFsVwlLlz47uRFB29FAbaZ5IcpXZ
kn6eIDKumkOc2kuNfFoCTqiM+a50vZvZ+FWLtF1AejcVESvEb3ReflJ6CnYVzV2akumNHFlj5oiB
4DgdzqHjhgVrBV0yWHH3iVxqUDOwXP1YQ6cWIOnuScmRUnk28QIU4wOcMFsIKBCvwcL1DeBLO4mW
xuwg5Wb1k951eeXAv2WdiBi0/vQu4VscVJYjFhPCnMjdpWByis1EwA3rHWjCV4M4q6958pyxFlxz
BiD7/GD4Ukb0vVRK7A5+Ier/4zCsRMajY/BAHDMCdJ4WFE01NOS/80zRV1HOiSFTSSjNmJxBQ50T
vIxVTUF5NNURubGgF37M0r5jHMNaPjqmLC8uIqU8hRULhRrljV+lRcKks/Zcjq/HXMLUsA4GKVjx
0076vi6mTa2XymsO6fdL1srp07cZN6hqxfaWGwYXgYlmupnEUvvTDwIP0irxE2xlzh1JHyRoEFsA
NFmYVoHDfp54vUA5+JFxJPgJPnEaj93VIeSfzHpKUTF4NVgJB2Oe2UCJCBr3fqw8MTQF5Q96fyiQ
QMhxuUYvZ9unFwQTjOO+PAzEFYCIOPMWc+meEimujbqvTGq/ppiriDkIYaTZEZCHbm7Y+FQAXhgZ
jf8lhzEYBi891CfbLHzxDjThfWsxgiUG0o5ns7GmLIj6Be8AoyXl3ZGBZIETaXTAXwSucVPbBnIw
SRs7vqcjVNkz2mDdrjKFuIda7akOejN41tFZvdAjB5Z1LQ1rf76QJwYSlbcBPlkZBq2OLcPZexGs
fH4/1k3lzKExM9aRWfpKolg3T2ckW2hePzL4YnKkEtNWM7FPn5HvgStYNLihc0M63BrE9fMbvkth
UetG/6x5n7i/JUjrgptVQUZS0WpKAVb2pL9vmPra1XgJmw/8Tywt5qZ6jQkuyDY7tlFR1wT1ofgb
fjlq8xmgd14DvFvTwEbOKdx72fqMJxkm0B/Msp80w2OiM5oebJRnDL3ruXdGKq9DzHEVgdJCklza
AgCGmueVViTS0/XTyehydBtodyHq18R6zX2GyS3O4r9jtrvTECzz443h689KibLnXJ4QIOeoKE4y
LvChE3xBkDsYb57ZClSSBnA/0Vl8/1SSC+jWPjayS1Y84xRV2lvtYQGciUYi/Vdumv7/ECAqPnNP
IwGO5recainpELa+ZkNyDuk4itGhkshNDNZijtZkKCQv6hxAF3s8ZV1VKuw4preeLa1Xq6HyZdoL
pizW83HusfKabmQA9w3rmdi7rlNtjcLGxXO1zzdBBXkygjpGOrUudbdwp65Z67dXbrC7PkfF4v0M
JDFNm5aQVelyF1uacSBRUl7dGeU1CPXyk5xhocz9FbOsX6mCp+3zU2qNOH2TWy9aVhVx9P/dwkdq
VeXAmgQ1Ilr/aHMIbjXEeEUt3F52MyR52ExSH9C/bUR9gpJ8MmV7F+2PZDzG24pRnCXPcifeH0dc
KETr+kTKsdd4pvEoGWJtZ+YgiIrNVXyuwz6MG5jHne6XPTrwG3BoLX9U4PU9dvzW7hn3XargrSM1
EmYXnF19oFGI9sZIeNR++4pEf2iDfNi6F+lei7ccWVez9FnufUi4+TKsgLNem49Nzupxw5hdOTJt
2Skz7VJ6nc6mowp0rgjCr1M7m05kH4EVeQPDOM3Qqf/C2FHseNaK8csdSIBbEgU6pcYrQHmX+owp
KbBps3YyetE5rLV4CU0PJktCW7RHf2YpDBuYRQi0Pel0yCHLGE+rl67+SWf/vwW5jRTpJXrmQHGW
UiCQLcpuM9N6KH/KpcGfNcILgw11Bi68wgG6cYgUGCIYyhXvbakBigg7UPunGv1H4bi8oPPmNDSR
zHqghLZLwp0QBIm5fZV2G/gmkPmwyXUGx6bnPEyFjZzKz3oDIchNII4kgD+rVaV1mAKS1z00qZem
Il2xOgWw7OxsgkE4+H8PQrEgICLKehfjrhZLro/XD9aeTb3y9BxjTF5YyF/e4XuGlJvg1A8tPVoq
3mh54LYTDNMpqgErW8K4AkSVeiZWLuLn/R2kBIcXlOXKDm1rIRWG8Mzl13QlAdM+wA73Af3hKpfi
9q53mVNrkJBOOl4/J6qLJUyHLltbp58PTWzvJamMLC5WUNf41bZAM0a1guL4mEHbnX6aHoAXtnnu
GR5WVak+HsPkVusFnORPJzlytAFFNfrCXuUPf4sb9e9mWetkLj81Fbu0NllBpH1+OYBt9GPd4RR1
iZz4YC4WgBpTtpGtah9Wkdy3P5O1dQE2IlDBkoBkDYqAQyEaSUAx8QD16Pq+Q3ibvAi+v/rWIQMr
QfBhZlKgu5XleFLVu3PJuQ/PciPDzWfai/mdhFPn/+1vIvR6HcUbQ73Kku6VVX/jr8E0TMF85m46
1I4FY62smGK3xEepdeR9NAR0ZX86eqOmwQvvnQXuQtqYRKhUkJRkJJyi0f1xpTJ8eE9r1bp3Bm1M
QuZpfYX2CLbQoIgyV8H8swOxR2O/H7N2Nqp/Ope4IK/+0BUYby7pgqmtPMdCIoeoPePtRuOlO58f
8C2Ibhokgdh1WlEvNZriLEL+C5D7euRUt2KwWxSfO05UPGKuaApJhluo9tKPHSE4Sq8lOuzr90IL
+7koNSWJArrM7sWz3dnZW51Ru/H3EbRuAYZPjNGAo/ixpEi/g3L6mwHFPMd3uWlgJtFPk7nT0mSi
/3xVgRyLwf/c+Hjm25UjlFkRWPPdrf+OBzY2Mn99CI+yjrIl6/aUSMu6oYz2uRvyVuhb9s0FGNgW
h0cCdBHseZ763Pl6b6mZ5Z0I/UvNEaA4sxfuoTE9kipkkwP8vYNcjT77GJwKezDEZw+FRFnJj4ei
+E3Ei9rIsdlFbGDYTy+YG8+dWqo0GXw/FgaxXBOUMCjmh49g1R/klZpUnnC23EHrhW1HSQx8Havv
otjw7wekUJLxX9T/ElLfAXsPTHHLzdhzbzWicFihB7xTkMEPDOdbt+HS/b9VYgzyB3ertG0cV3uh
CFyn/n/3IdwSNhB2zK68a07jDRnTJb4Y8gOmxlDY0h2J8ITuTFTTXpxeZilmp9wQ059t6oCMZXow
oqKtSNwrxSutmWsqiItbD5nIHuLnzEEVqXPLWDmm2ceNWb1Lz0P7ITUhkJrh9Gr4ztRGaAkEqtBM
dfPYzj3lscAtmQfzJtUZVcW/pnu9fPHPbLvVv5STidsKgkfVmW8eHx6+aRg5zwy6IIOrgoQiG7dR
D62UrorsQ7JcXwPVgyIzJs/ciadPRc9L77h0Hd6bF2y2ffIb6Zqr6PbTre3jurtQTRJ8k4PBFgor
IGolkKVn8+nGJ7aUck3G5JYRBrWq8kacDAx4//CbH4vDDM09WMmnwHNW3rakAe1IKXjtJxlGXgqS
ebZG2KU01NCCYUdyTqJMF7vlUgwZ9YzU1gOjviOYOUm5cdUk3d7S7kMO9iOclVzlEmMvMltxPoLU
hyMBo3PF9FzK41tyWbsb2eHlux3IX9PMbspK35t3bsWmJ2WlkVLiLLuAj2VWJSSx52O18AEZUIri
29YNPWJadXttnikIaI7U4AvCJshsal6NotOQZN2Tpm3CENmzr4PtFMQ+GS/FxedUHuNRz/o0LqcZ
VAcGiTA8BcdBMWL+vR0Y9DJLyJqsCsqf7PKrRaUr0oms7SGMXLh4qKpCA98sp07k/xIEQRYVkz5T
9TwvfrUwo967bA1AnB0uo1qsSOtlP9zyuZJCPeXlYNu2ksxbcfgfVFVbZgfLi+CcLdaRQXJ8ohmd
B1mX0knluTo8z0PvqjuAQXp4MF1haWKSaXEnR39zYMZisVrltjnv3PHQq+0ieJYZk5yyhcD/DWME
CpNkRubRG5S5o1c+Kb45cXUUkrHJHyUultUSPaWXCzfQddjneFlaX1v3nE8WM/jFvY40QjPHe2og
66ioPg+iVezhfCNMEPDSUd1L+NIkSTp2fhsMNgeMs2MYq99rEohxqd3eI5dYVDLqvlwZMgNgn0tE
tKK48HwFeBZWgTR9GytUf/4oSIKC8Z+PBfpI3md55QTG+lpT4TvmREkA7YebLNEaH28ekXWV3zN4
2zqLeLBDl/NJVnnT2U2bi1JJbdk2n4ECYJeI3PGCLOYuO+FwkT2PxdBgmX4ZlibjH3jsQHpZQbK7
pW1ec9t4NfC+Zxr3iVMjH4C3z8iSOjLwmIC5y82vJBRb4ec2UPH08sdYENIDP3lSCqDJ0AmmDES+
QcmHKYVSt1r94VExsgCwBkqVWFzecfdgoFw9j0JyxdIaF3Ri9VuaUyrD1oc+ChfIeh6wZHQrqFYv
H1KS5sHGa2upEClOpBAQcoJUytC07i5KMzBsH07+1PFP/UzGW+94TX2khxp0g8Q6wtu4yF3GR0/R
xycEb9woURxLJ6sAuf8FChQEJtK+tZezaOLGEdYiiCujXXCyd++TV+Fu/Ut1OtlY6DCAccXQUZLG
90w9L+FbDAqPYOMh9g+7IdIcpK67UgXzebFYwDWBnLffWO9xZhAXbmmzLTBZXtxCIQYnvhl25ijh
HxyLnrxb9+AmIoPm1NsJY8PvrmkGcaUYdp2cpoG01fGsFO0rbqA91pHwdjJcb4+RKFbtOuhFeR6p
ylpEBfTxgfWJyV8gZgPdtkhXc88Wba0KkV3WPGqW9mH0nzrIbhYYLpGqzYEYSVcOeTyaxCG1+ZVn
WTLO5s8zVa7zqfO/yivZxPkOfPZCRd6a+vbsRiiKYvoz0lesqjUtLwsREn59Lc0Hy9kUelXRq2y5
lP+XFSabijDKx7AP/gCzWaHM8v/g6Te3YBAUeYVCSM1jhn1KqDLxWvNaArUt+6SfYhlv1ZpfqDn/
D/9rkn9IsNLMQvYbIHDtVKszTNeLcvR0bzNPQZr7Yte5Hc16zxaMAAHx/7x3onuxgFIbOellkeOz
RPElYAZxZEM86Y26bgwXp03Uh+1GVvMP4bi8I8tvyxsqAGGB7wIH3lYaSTVuTtXQZ/6jQj263KF7
sOcrbS/1a/M+RLBhYQphpLSF0S7dDYTDNY3FGcgFIaTKkZ+572kAO1ZzAv4oYmXHhWDmLXT8ul7Y
kk9eh69lfg5DozPXPhXm+4OLH/mkOhsMImZNBvvftHrMaLOqhSgX8ZUNjeo5iD7/QgJUdvlexCtH
Sw6OiZGBRxLF2ecfArFFAgNUNAbjrEDAv6Nc9bTz+P9FgN370GmXDQjv68gsDK/F7eoOb0snuF7+
QA4e50DLQYUNzxD/YHeiovyVrJECGyxGvjdfjzWowHNV8u+zBoPThb3yQXrur8MttOiL+3OSn+bu
G9LH7aR7lER6CcKNsDbpyBukEk3Tiwge9sIsuW4ZrK0kpPcLfdxRJpFheLzVbAcGGZyJRh+6XDtc
DrCDcCYXLdL/qJ3CyTTgkgQiDgc6PDZza8r/kSu+JKh8PKj4/gTmN8Ed3MjvtYF90LdpUtvtwoT0
6F68zmp/nUTe07YMkAjKP+RPMiryClerPryqPcziBM5vFvodNI4onOqm904ricy7tEDlVrwOUekp
ytnx4Jwe6p23YHruScu1+US9S3d7dyCIK9CsTb0HNTCfdKMHWCLJo1Ham1NRIjfbL7oH2rM4jdVD
+7s4KbIsLIgmBFObpTPA8L+M8VpntRYjF1cAHRwnbuZE7gl5N2UHT8dOrhqJ7+jRKqHkUEbsF/9o
xR0Jq30FPN/yY10ZmCx9ssMCYZrFc3KhTOXV8DOz5iqRRt3ySyp02Q/mS9DbQ47NV6VhTHnSYbH+
UIHcR0GqP61DE9ME1ke/kuas7Snlccim7AsDng1t6YcAg+yVbaGCBkDfYh3RthP850fhagnpYtf8
6/ZHFFKmsOn/X03BBQwjmoYrj4ojajyLi983W31gU2cIqD8a3pZr3V/vB6PnkcorXSabo9Iq+kq8
eakeXL+A/hR5CBRNtn5hy8hU4gRngAMz5qLeecwEvnQ4PZoYCHQjFwzbvKA7YXtyAANPL5bHtAKj
qqAMXDODEt3n6lGpUznb+GObHxC7IiFJkoPqouF5JQzwWqhviF8OONah0mDN2bIecdcbfDeH5y7b
XpKzk2DW8tbudf6Fb9+imhI0qFzDZ907xyx+hGorutVADYAusiwQfR0YXA7KT91uR+HxXWT5eoZW
YqcHnHHoQHKrdY4L/MuQZJ75OGZTxsnixB95veuyEUujI7gZ3tV5DpZ6NLtysyy4WTYKDqzyyPe7
5m7HJuMFa5uZb+tu3hSSh9wuXOS+4uqMeLgN8Dr+izvi7nkKOswndin4KNtHR107dpdkf20xNOGR
RMdrgU0wpPZrHK1gRZqjp3RVicKu0I7kn1zrPSS2aMnnP7LJMwVs+d5jxoMxqCwFaTuXA/aI86eN
E9WqZRMSqjzD0pG8KT6iFqy4zsN66LL0O+SSPJJbuIo9aTAiyFGAjqddN3Ue59afHqcpxCwP6Kto
fizudZ7wW7m0y5oD3Sqnv+/UVMcRgtDe8Wc3HH4QaycrwtkGUyqlX1rXqpNw6yPC3+RVo41iGvPK
rq8HUJaiXFhCHi6QdQGI5aKovDo0lp6Ks9hHBm2sDzZuAEa/RB/3VTcdp5wtvU+fYZMpGOUog25M
jc5jjMnuVD42C3zpjJsTEurxmb7CHnqh3SC32NLU3ezUlYpcx/AtOoV0l8eqBimMqS7/ZbxZtb94
dUFHIbnpmy1p3LR6pIsXrFOe3ITu6vPeSCdAcde75okg+5LthHAyZeIHsy5d+fvLNi9h6R7cKy6x
OrU+aBBHriR0wJyLhPuN+JW/jonkw6p6PU8SnOxCDsm8IagHAkhBWunNp3D6LaihNNKuIFtI8H/f
fmELBkIFJw7AQBZYI4/RcuP1lXNn95BcKoFQYm3TX6cCCxJtMuJPG6EAl8+S4tgYXvJkEWs1E1BM
eMdJAl+cej8bdrQZArpm2jfG/sai6hiq4aTCWhahM02EN7wQs+lxhleGLtgpUKnY2wQYspUqm8wz
p/UL9JucW8enYq7CVa5cwKnuD6INIGlKSpKNzKr2uJGpUOLOgbfnrgnGG1YzuHFf1vhqicnnCPOQ
BDip7V3Nt7O6rR+knkmFyZBvczrFk8x9nm1dkA/RiBy7EiqwmslWVDZ29DIoQkCBUI7EmX4RaK1u
g9PjDVsXvVfGsZOcM8Mu9/rGhduny6mKoFvf303Tfp/A9Af+FINNu3bDX+NNcJBHLFOsf/Ttre9C
Ts03m/jabqoJL3arfmuPt0VX+L0H7y2TuI4e54EBEU32lGoNKT0Tg1mgStKFZpQB6zSqMybKFwzG
kGkoMkF7yZvuszPuGKNWuoAYqeaUibfj4EwWJP+7/ETb/2Ea/Puv/I00aDSupYnTWp/62WdlJNAr
lNfnDivZsH1wvqi31X18dTBFD9x5HJPztJvQ7uiu2sXqpipo6Nkzm7fnRCkR5XGClCYRBExb/wqJ
zCFki/JSsOglQUewOEcP8+OcRy0v657xXas1CvNVSaF36V0pefDa49hvLPZdgkKw6ss/bx5U4dht
xkcZNvBLPnGo5c9S6Y4RFoxAkWaHHWmRj4ojtBKmgTN1TDCGQRKEoRbdSikfj9IMBoReKmSVE4Rs
JpqqSvkzv/6hQkNGyYNnvULsFPdFXjxfdDXptQlSeNpbfw74i+4wwFIdaJtOkd36Lc9R0Ry3FtMM
ETionwRn3KAnFp+PVuAIH6keWI59im2vgpY+/DUii6jL/H78PQg6n5RDpbL7JD954zgJiX7TXneh
P6NbZOjihehpyImIDK4YklTV0TeCdRIZaTfhghLBLo1dmJvvWsKX0lVLGNr6IhajQ/I1Qpku0UYh
pHgyD1vAm57Ml+F18v8VLHa/e7yclcvpzPJcc36FfYwVNf/D4O6Reeap5vzLU7KGwJJhqz+uMi5h
iNNhzPyBlVobqRa9v1m5LT0cVByndsisCE+L3njbXipmWozQ6abMl2DAwkfBphxRHGbCK7snxmoj
b9GhR+/2BGysMgu2SpP40Nx0RWxshr8tylQ5KQyg8ujOTH8rtTdzYdgSEVc0tou3pQ6uh27WQujV
sFgVsnOJEBD/uXSdB9/VwH8EUxH/Sy3IT2A+FRgCihsSetHSsIqPVUGrUBDrtMCl6tETtclzBlU9
kYHNScn0948KfRMLr3ycPpTfjtQakw/ERVgCAS5Sp3fRcv10jUF+8FHc8sQPXM2QD1DYJp3zkVR4
o50cv1M25AwagFDDK6jdkeLUwe2rAofpiGNRX5jb9c5+2jTak1w6bRhfG3ccre0JFeg2XxeHT7VS
YHD/zuF+Pw7oZfDTTuk8jCz5nxM/1KoNyS+sLC+zWVEquBA8GMSLYb576cMQU6DGpHZZlDp1rytS
5bHKlEAUdj3JXmOxzOK5ea8ZbJMI3OKm7b+lelXQ1+u71qReJx62rxdBqA/kP1I2YEgShjwuZaF6
COInHHZ9oI1M/AfVRvdsUuhwLGVutzpHjSEIQUXWwOwl0KzPVk24IIZ2mvqnOC/jikhoteAnDJKd
Vw541/4wII/DuQDVo1yrr4ueNP5nC83pCFPhS2Kq0/tevRJxkLPXp52JuCIxPvPtxqXqADCkpu45
1c0sP7CQoP82leKsE9cZikNy4M2yZtwciCDFIAZCixT4CVoRemGae85ATXuyzx560V2Filk2Ua/B
x/tg48k7KOai+eZIdM3P16OvvYFMYUZBW4bOH+dDwO//xYVyEmeqoX5aXotADlhtrDGBJWQ/NRs5
SMo4A0juwQHytxvJgjQCnGlqFe6/3Mh+QMgu/Na98Y7f7aNvi+jZxTqlabRMGg6NPiQXlIUnNUWN
e1dNSrE+ymeK4SweEw11+qC9rjbWa//uI7xEyLlWzNz5ueRkUZZrrR9jzMeiX3Ard47pB+gwOCDq
Kjhe/+Ag7DaI6zb1nVVO0614Wc9+SRqSszK5g6UWNUD6mGEzbO6W+oUWAtqbi4L6066wCG5NHMzM
ko2iaZDhBcpCVz27yhqap4B7wBPjN+RN03FXypHrQaOw1Buv1MnvrDFHbtp0YRcK92edF2PCZnqV
Ay8r1mcBsozZVaveyciJBUWkeOZo1d5LsAC1FdjV3WbAoD0tJRXSnbr2vub3qIW+uGk+khwnnxM2
N47goDF8YmN0ZmUyZSJv2PaItLllcRHer5kbAgqBMRKlf+SRE0MlQ5o0JbHmTEwcdoDIY48t3wyh
6JKAli7/hUlgSWCY1KkI28duUXDVp007xFFvgxB/YVtY0bbRf+0SS+GSonhoNAQBYUUdjKcBYxle
6RvIqijBik4lNf8htGyZsLXhZj5ZptYSLdnQvvXSkdmU3MiUyTfs/c25x9cOlAlvmUqmg8jKY1Pv
ex4kTvraZG4XHf2OYhfjNwRO44ICu9cgbZwCAE0M4Cjfs+dt6gyBAdNYABCbWLJqK7EMHqJ7Xq1R
Z2RyhUhNIIP058lvEB297AfGw755QqKkSH/H8gs1SSM1ZvIZcaoSphDDEeLzRr6qeO67vu7FLlxM
Zz8UK9PzEgQPxSIBYBfcGFxx5irrK0hpPrCe7eXDq3D1qirguh7buVrDAEqT6uHiV1+Q/X4hEAIX
/YS/nk15HkGmlZOcr5TzcBURzei2MF/+AM9gXE2TvgUjxzXK3Ny5/IiLCk5iHBywISpX3nAiPQT3
igj7b5AZjGPC3lAxbym0RfoxH8WaHr4v5P0HrTZdQOK4TgAWi3F/8ZlqTT/SRIV2/aOavjHulj1o
DKmXcM2jy3+qCqGiDfnhymcGyc74FUwuQjOldEbqdrIhcMlicDJFIkrGQN2zOQajUNIkxHMrIvjb
kOLgNp8LTLLTTnBJgACLQEowax85QONNdaBhs4THlLlpMhNx604vQI8HoEYNzyAeq8DA1vExWRKw
U6dN0lcm45olfffMk/lQo1ZPFxo64YgjrcZ6VUkrL/m8mBH1f0qAvc/FGIe16YpV/jnHq3AiJKVX
D1UrzoSHnCsZFEEbY/X3zjVMpSgAOPRq58jVLyUooDvDEssphJGlruzwt6GM4+1B6F9DWYcY+jH0
i3o3U8mQeFKq4xLGSnQHI9CH4TRocpJtWe4vITlfioyznn2qaImY08uj+DH/gA67V1u166uLkSLA
JYGzT+N0nxV+Xu0Hc21VGaO4uo6OYXLhQ5o/ZN46m/x1wMndK/sIN8xkT5XlZxm2ewXVEWaBMvRk
kEfVi4stZOWqF4GMU/LDNU1UdFeUUD455jWZOSszpsoMookkcPZPMUgtiS/BdjKsv3wTyIIoRbSx
vMg0b2oUAFTA+iwxHPMsBIC6mSolMSP10evWJdLi1BcMysXIpzBBvFMnUb75VYRlkX7QGO1tAkwe
6bPRxadW5e9GD4RMKqtNWOp5Y/pyh3Z9G9SMQdQr8YtbS712ttVX0bjlcwzO0cMQCQLrMHk4JtVY
Vfbcj66g/45mHa1gAAS/fBBYpylMPQx53nmhoEUjDeubo10diYPcD2FBji7nBR/3MdFjGu1AlYxp
2kEFdYvKILtkHS930HK/DDuxNZvfWSAg8ft24j8UydZ5xTwVc+w0G5X4sZzmNLvNTyaDnxDCxEkt
itLlILwp5kjRG/325d5lW1wceoKd/4dOW0PQnmUDObExsmkTyJJjKz3jVyoB9DelEaXDhYJ/gtGF
0BSVL+WD/rqcqYa60Zpeof+69v+v5p+vE0GS2sgV3TdMmdeA5vLJq8uq+ZMiHXGXEATqBW3Vl81V
pm95iW+jICyK/BhTkXZmsLkaKgK1zNqPMCo+pmsk7naJAW6Nt7EUzCCMna4RvrcnUj7Fa/uFlsKL
F6PRHslkQLi18lNAkyB17+tZTESKZYR0WGEoRu0Xqsu215eJrudPiJy1BMLdmlutA3O+oHUizpW+
9kwrzVZLYO2mOw8Vlzdwzqxhqlf3fcAwb0J/3tdzGgKcqScPU6UVB+96vatTE6Py/KGuL0pLCpxf
TFU6TAjlw1tIpkIg+8t2rIJDb98D/47LLfCSPsV5XESuvg2vNDnpV49JcvqriQnV+bBo2nA6+sp9
QNtgOCJFpaQ8HN/4MCPSI8ZniYjtvQivNygVF1GfAi1n4wt8AUx3NCMPyzmpjoF3WeL7szAYxx+P
PjRP/zIyRnXy3u+txcHK+99BGYRdTDbeiQOWlTKQRna6UX3qYXBuzUgU9N9wMq4k8XnHXayBN7KP
wlL0O8mYs2axcuLmdp9vXPCTwZtsVcHVeCgJS2EiilkcmV5CyOzoTrSOi9Vu0ynSwxmYFUKc5bdh
avIXJebJuk/PF+FMEVV3H+OAiZwtzF+/XE2C5vi5uwhNz/nTfQkiYcJHEsuyh1MaGKMWgJy9Kr37
1++5+mM3U3U1mDVPf/2LeBtFy7JuBhAAoShXga0J3GU3gB723Xf08rjqh6fhXbUi5f5SBoz6LIHD
RnDKqX7sMX5GAZCtPoKKJmXeaUOfHYC9a9eShLoAL5/5FDimTrQTgKSmGxWtS4AO6Sb3J1vYpMxH
4LVlVsSItSgdU8C4bGyuCRBEAXk1pUjTc9cN9MKPeEMco2zSsLk1cOpXNHU9oUNib6TY1ZwuHHA/
CSp/eampLtuDoVRmDfvLx3RUWQDb4fsX4EXKk0KEZjGH7PNrRwYVfN6gehALahu1Tsr9oj5kL0cy
dZIcue4SPiS+KEWw0GxWw2fWCwHKJTviD+HfsleP2LG9k/PK3O73TGVSA9d7990nLdRvP4czlqHc
+TxC+/XsaMsyR+8AJYf4TBg6c6/UY7BP7M3hpzUfZPDMPyevpUUq5UYGYn16UIhJkeZ23mI4+AI3
R/u76SI46F4lulw3TiAu0JTf9pK7Z+QJvl8N5i84/9vbVkeORRtuPWx+LHGj4NkqRqsDXjMfRUBi
jx9mfZAV69zdgdNsu1yspwo9CRdflHIf+zj1DGCsopq3o7Tx6fwt+orhjEXRDyRPnpMjtjQNVSKh
nqsOE85lAGdzIIl+cKevzsONFgic9ExCyBrEaofdQqOtaLyISqqNIPN8i1VOLQpmR6EN0IzFf7WI
KU66WUumj42SOFsKBSQ/V4r/h28W2fxTgkxVE8trtlsL6gcwKyfnyDMnJiY+4sx68PGQBmrg29Sp
zxEEMeBqhwJfaidy5qK333OBUe9kVQcgVeBFTFBeC6oLTWJVKEvkVVGyM1r2ETCY7tF5JgHzTVJc
pgyB7mx4iOOpGzqRm7yuLrtVMI0pDSucCNS9XqpYw+NUy1Y19Jg5sdaxJbD7NiTohHHp874rKZW0
P+183QRS16A4xxreqKOrk27pfvuH9DouywKQrqhPLt8kLky9DGdbXg/Kciv9xake6xWiyGs6eqrH
g3bbe8pWquEKolGLQnc+dcxSvvNRjg63vR1x88Gg9joXA4pj+Slkq2FAgSegnX1faTzU0tKutshM
ObiASsH+a8kjcwlikDFzOB35XLczz/qHZ2q1orvm1z2p81ok/CeN90Zgi7PUp/xeCwHNM3MCeXER
CCvDHFj+l0PHZa0by4OUVPaAFQmp/BoFBWhdYjfvU1htTIX2RwnOaGI6iTniqIehjX/O9/7D/XZu
TYgQvmxeiQVdMo+jVF1q3AubkJQztScxo8Xn9uNL7r7H7I9H1Cx8h6rlsCF1HWLTqd/vF1KxUPLo
Khf0HeJoKe4zyck1xWPAEChcbjApCOhN8F3uJovksPFt0tzvmmXkeK4uluGeBnBKb74BK1YHqmsy
q9H1kbmIZwqq+yjbPMMX/08hBi+8mKHJ3D3vHaqTtRvG/X0eQCz07HTx1QlGhF99u5VrnJELye8K
Li9yDQ5qKb8VogM4r6T8kL695nmh7WrxdafHAualWLRclW2qhuHlpQT2v7q62HbBfmpTVqCrpl5C
y8UQ9nLHWLNUFQvgOWEKbzgfQI9Fwj3qZGeTiTSkBgj0ogbXPGbZgw/oeuC1Cwi7euM9RdZYbF2p
sYLsVI+w9y9M82KQjwuJICVRIzM7AWbq8TVtGPSV4USha0nvZSClf12VDgBxLS2Jkf0fmiC1PJAv
1lAAX/X87Yls3v32VXmSi6j2kTuGQdZ8XU/AwmqRdO+HuFpAfsRzSm9Qp/c01gin2rrJMzd3fa4i
6i7/fEDlF07xUSmIA20daGsZJTQjDHFLstB4ZVTASdorCOt9ZDAgP/TYyG063A3vb0/t2jV/ZF5R
9xvEKd9YZM8jaK/x7VURqm6+UBsSc/2LJ1rjZfaQpZiEsENX17zGjdSac2CyfDrBD7faxbVPE2fD
j8ymQ8BAOhEFQKXvdlAdyDVir8xgwD2iAeYklprl8Apo3asvD70r/z1E1RHzRkMvy3AQqROyLWbB
kaYj6Z0ts3y8rS1IcfyG9hIJZduRkVvq6chfM2uNpPLIguo/Spkn6mjG1385+u1O7UsyggYYGcY2
I+mXFUSuSZLE1BTnUBYQjfqwfnZ7teQRK6TNzeVyMxs60IZAijXfYsBhdsAM0K9ngp8SwgHPboJy
G1ZStD39ypJyRb1zN2JDJ7+i1L6yDA4BcgQEqcIc198nS3yvY07HSDAsTb9HGbvjk5U4aogUeW0l
UuL8OHoBtYuup/QkPe+jDPMX9rrf+hajt4rbgmTnnfUXRZxQS2PqWA0Chi0jkIhOsqkkVpPA3SVe
SLsEnCs09nKRSCT8R4Y+HcPPAh1DopuMGLG0XzSx/ZnHk+uEz+SxLAKFldf14Y5JcHGGYcqs+myl
x4P+m33/Z4DWYxF4fcKRY0aJrdLat1UIwCt+4TRFnrxJx/3hgsZfgTG2joXQL8Y9OSzpWfb5tw+A
KeHQWwNeg96PafUtWlgvoLwJrDXQkUrBhTCsXEIc4ODyn1uASEZe8KhSsKi8PkrPpgClEAhZEc1Q
aPbi9TFtDMM2C+AYKaZBqFJch8yiC5/0hJj34SC6+4qQhDVg6wgJbd8jZF4CYi3O3iaKS/hzsAlw
l/ExV67cOo5P/YOdwJYmQ7tI0dYDUKdI5xvfwf+QfNULn+psIcyIx36veo3A4dj9bnuyctKxnvZ5
eLc3kHYPdRSvBeqNFSRgbBC4gZtMzC3JyqcVPRQtBHEK9eLSq03XPq6N9IkQYEyDZ2stMydwh0HY
sKfuxUjZZADTv1xm4GtRAuFQCcDKcLtxZZNWUb0Ma7rkd/n/kBXhBuGhADC/DCU9Q6JrPUDbeSF6
sjZO07goHI7jWxs/xJg/iq0G/4LCKA6z+JCHdiUFRqTysQpHfa3KKC4TZQPe/+hMkEO9icxxJLdm
9iZgii8A/uVPS2ZdlJjs3qZyZbd97sthSF5Lmz9y0hfANu/VZeq3mcAz+tDHiClnlSTRBZUe+vmL
AqYNFXJsgRUyDv8ujL8XVoI1GjnIxABSFTxh/la+JXjd5pwB95iqz1Z/6GdgpVThZ9Lp4A2t5/Mc
1JXi+zIbYKvZbprIKcrK4vZC6RKEK130dUus6MIOZf4MvehwkixYI1QZr3ambrI9n1umH/MxNvZ6
E9EmV52MAHL6rdK8h98IQ/o2DVVSHQlGGv6gZcPv5rufOhj/q98ZX4+hqPuWlnnYXvlpE6RclFX4
kvfah4GzEiVJ1oZlGQQoBqc+YeoQnChToYji2sNHDl62TtVE3Q96dyR+AGXpky0kcM6vd0qngN/R
LKja4gStsbQkmSHfTs+Wa3KVJqodOe/yBRkj7wWBf6Cd7Og+aDM5fHF+2JZwNWaGJme+7ZDxnKZl
1JfterxUVzqwSiaotrIn0NhArLWBQlO1mh/nO6PmiaXPNDSRTmEEa1/FZ9NTuwpOr7u2D4ti08gb
2HHJMduexG1zJ7Kpx7UF4MRYBm2EaVXRrGmmyKuP5djdgbPqyhXH7Iwufh2WQhPLWsbzC5k0VWG3
Vw5o6DrPpFeYbD1kkN3c7y58w1kfmWYpY+5tchyGMUDACiRmroH2xs2ok7KLpRmbi5XzxmZ9rQtr
kzywf/eonz4bUdVWkTCISJZ94zErn4u4vh9/AFNbE7Nzh9TpidugkYSdb7nB9wPB+OricWkFQ3cA
iPPyz5T1nNxi4ewSzy9HA5BH7Enpbp/3R1mzXbhD4SEpargMAUZqab8zqcByJe6UN7d2kL3VeAx5
Myx7kpJqUrRuH2Ee/iaMkSEFsTmCI7b46eQNz5dqLxwu2uVQP7gjZifuhbKgVeoq2V7ZeWiHNdvl
+/KrDraw2Hr/POaj4oR8tBSY4j91PWPYG9h2VsfoIOeOBrzS6x68x+i5Fz3GoC05MFvlBVpVMxzo
dEfBs4yn8J2aLNJuXkQmSYH2yd9BZ6IFJqYFboyC9WqGvLV3UG1/sAIZwztp/PT6+lFA3cpA8Owb
erI9j0BRy8mobJEFf9IQN+5kHyp3o4DpG8HLenAIkYPCIA7vv09lKLlk1utKukzPjwyM53ijpbFe
orSOfNr7MugCBU0kwODGfWkksCiTk11Ts7TYsFQ3MTJRQ7p/mBKlb/M71zsiWNkvqwWrgmrOUrkd
CdmPSfKNc9M8n3NlTIsEC3wszUoPv9NeKf6qNlwGQpsZspyMSjpBc2UwS318cPL9I+OR4j2BaBY/
NWZxWhkgjH+OCX1+PDSDsAQrQf4w0FpVH4U/DVc+vv/GGrHJZv6UD45knLB0FqsE4+ZwiX6xp+Ey
d8FZP8HpQO2Q3CYc7OyAfT2j2eA0rA9fH+0YSwT7DnOGmNAlTa5thddEgeIj/5D0qLIdziMzhTKL
zZ0oSS4KAz/EPiIlNCJO1ibDwzfS990Lzz0gkG+1mkkpTaBD2dTPgiUhMPScBRHlkXf5c6vLd83O
Dz94LqowehXDb4jDmnGeGxdHL42Mdl5NmYF1VxmWwEOKIBEmyudYqh6M70qAISqcYhjdsH62mPq1
jFQY0k57uNEmjYD0TvyUUTdx76xyPUdWlyChqH7g4q+biQ2IvLJ8C+hP6WMRF5w2jO+nmxhp3dmJ
V/CzpkerA3pvK1VC3xQmyaeGnVFGRtpQG0rqxk2H9TVACwdyPyjSQ0bxGlMc9A9mJITdc/GxpAzW
1sZGynIWTSJzI06A9yHMpyJgkvgIJOaogCDBk+KJem2mJp1lWo4cku2aC/XT0rXphcYXYJxF4jeO
qeQ89SI/GtiTPynByZI6EV4lROmSrYyOgsmI5K1QPrz6TC8v1pKExv6FpZ61Fxjzlq8r7wWi7HnC
UvgXW6KpmEZEZFfidJf6etUlIj5vole7OGh1KieAtYVXaYoe/TYuFl3Hdbyqn47DmAryQEYbaEu/
8wWAqstORkoHd1zb5uZImcd3afyh/z4FCbR5NGLjif8sXnzrUhKVhESR2Oj50FipOg4dYIpXf5Al
JaX1hkWtIwzJ1lwb9rBb+sbVsIBL9x1VX1Sv9cR1bKyhaUuYX4/1lsc5FT6EoNbXW7PWWJM0wdmW
tt/E0GQKiE5lwdK7ZcvFLZOU7XAebkWjXr4uKyOCcyzYrwmWacK7SLH7mLKKc2zSi2XHQ0rbjQph
mIsp4+26lo1sGdietSbd2RFJ06f3aQFf48V2uvoBW2rXhcdqMxfSkdYZQUEs/KWNd14GPkHkbcGm
r0JPIxJ6wAyUYrprutRUZLQJ/BSHasGssCd1BcckDQ+iH6hFcw5dZN6KYOne2YkS2+BWL56yzrHb
i9R7KM70vtf6PyAfSmDBVL29N7ewouqsVjqvSpmoR7AG3fROIyYnOsBCXllIihh3oroMBM0ul7EZ
pP8uM2A9KHTNsSTxnBILtl1TpIa7Z+AC4DjzezBmJe20gshhDtSkAF/dBFKVrOa4ARfT5XidI2NI
RhX6qrdpINyaHGrMUan/0DWruqFmvi5hoMhKxD9oEWBnkPU6E+0+12BPOLPX6ZojAW60nq0d/X3v
XkxrvTUm08uHSvS88g70+83nnglUzID7Ujto+bnYIe+2llSsVHmzOK9MA15y8ZNjCMKK1rQ1ALDj
LED5ylk0OgqA0YM4tUpc3/xHma/pcOp9bwa2SzCHxBjHC6KMhzS5U2djG/LoBqdpONP8GrAn63hh
MKxh0gbbTQL791qWROYxcIvB5TWGeUOTtMHOvkTDwIFzEyCIWYUa3P/9vjJMpSh1sj4ZXAhHsw8Z
PAwmU7mHCjIjWWYXMb9iPEGhrgJj4fUFfgPz5c10paUUjq6Vhsfd2ZYCg2Sj71N0T2er0MCekeWn
Rz7g19nl0czi9nCUIPxSEre0/NFguvrr6wnKpTNGo8pgd3D58GIfgXfAIn0vqm4JyRbFlnBVNSHs
1MezqnzOrxC3KoHUnwAWjOORsdxqgRyu1LQr+NiG9aI9lNgya6ZyuT+cbb4o+lhvxKobjYo350vX
UmaI34WzjHC7W9o35gwgleDg2aXi+ocoj+dWAL0I/tkvydrvQSuFMKLswUKDrn3Lg8CERc7sJike
VXjKs+VGOrcCjDYJnocCiUpIUMyDUypbMUjvjMc9eGWtYNbZeLcq9bFgCdE2ulTRcKtqnK4U8hVL
SoMtPmUd9i3mYe0dLfTSnObPlX+U2Kw91WKWO9bP2690ZdlurYhSavCO8DOQy9SlU+5a1QqOjcj5
F3TxdPp+prqCybd0oG47Nkdm65N6eslufB5n3nn7Tk1w0kDX/9ir3c295bQAL52fuqXp9LeTARXR
aA8SkWBPU6IsWDSr4x1iEQG87SUNdg/1p7w46rm/X+QAsSGZ8j2DTjlGSCadLyJd1bN3QhYR8J49
xgETovg6VgSZ8Tc7ZHNtlw7QkoX0Y2MBWujqzObkEcebpa7Dkx4pLAiiWh/JFP0yL57VqaF8fmgR
cEOUJoYjJfuHmeaXhuODQrCISlKU2LuPsxe6EP0zzO+C/X8Xkw9MkvgwDKcTn9OVazBDgiv+1agY
drmaWDJtHOCHKTHM7nNGxxGjvVqEJh39nS09PJ4fjBYH4K1zA3fW/f2ZXovfV+FHBtlBzcbNnMn6
+RnSsXJW0278FQ1mUaewy5FxE4Fll+Nbznro4V1MbfgcmkTy1ULubDefGBY9yMoaSBr5GbVxiunR
wuHTQArSLZYtIaWoI+rsxhW5HKLjpM9RsLWyFBN+KMCNbZGvcjHOniKtNzBdvCuKErJ9AdbfAoMy
HOIbPPG7rMfWhvzcTBQ0snj9+6x15c3t85qm0G/2flG3chqw6aue8QZLgxVJM5Exlhx2yghV4wZt
MQKTAZLcqBByhbNyPLSKVj03CW99rShKrbKtTr0BjTttOUJvI012aNlG3AhETVImaGUwUEVyqMTc
/f3CyECnxsmr0FpiJHOtPTBxnoILg7RgR/kaFPdfxo9W/or05N9/njdiSnPy5InLbYoiO7UxUC2/
xEsHo1LlQV6moH7LMBihJylYLYwiI1mNR8nJYOy1cLpHf8yxHQmWwOGg13vs8JifZHSYh2+x8OhV
i+fSV13s3tMq7BeHlRwTa9WgXJBdlp4UfB0ieV2RyFBwAU8TicUZ1LpAHd5cwOTM2HWx4vCND/V0
30srO5o8OnX76SC2zm6Df+pBPHbB8HoP6LOnm8kWlNK1ktLCPw0njZ/GQ3SyeBgRXTKqKtwJBm1m
TWF0eVtxPy8ueeaCWM/jqs6kg87k93TRLoxOshYqzJYnMcClC/1GyKm3qf8UXa2ogBw6FOsLiBG0
2PPsF9Gd/QEgyzHUmHdmqGpm8BHbu++QHtdMTHyY52nPQ1FjOxoZ5AhLLfkXL39IcmCp+QoOWr4I
kGfIhPQQLaktt9JHEp07NYdJlFWi1euspjISjnzIE4YUvWRvlRqMbpGcEAvcXGG/ZU3z3O9M7tCk
j5kAiJ7kKAaoDa5x/rEIxllmToElSpEL9b7Xk6gXuHokL/z6giqEmkB+WO8a43RzfDEa0AluBJGg
yEsaqxoXGSknaeMV9TuYPYwFjVB2nBXtlCM/V9LQZDGtneGbRGxifrhiHWfVYxw9aQX385+8Yfb6
MHSsPFtgfREWW85t89EXVwPyfu0R8pOmiv2emkGQQ0BQ3q2UZoN1LN6dfvwO4MOMmy4+sbqg00Fy
xRO00/WxgRh33c56Y1qpwqQD5wAwRsOdJInAngcG36Ivvz31W1sRVEEpR2J12W3/8mhlFz+WuOGJ
6H8Mo1WZZf/1TeQPO9W1RSgcWCVedfa2DvTvVQCatp4/k3orIe/DWSOoMpM8nlp5NoqkTpXzopIE
hV8d7uXVcwHJ3o05qaoxeeigL9aZkjrHX/ftSJetN6JvLt90AvcaizVpsnufocYx133QrMBEGxEu
ulsvETNae4OeySI5L3J3sd0uALyGSMRCKVxBXnszZqtzp20CMgTX9cECogXJuzLo27kG3ot/UNJP
7MSwTpkxXGUsXMfgiTQCmDO/itxUM3n46v3+D6eBArUWLt8ThBt3kFe95e3YswwrbwfCfdTgGvcD
7/9gQchNNd7RIBBVufsMXt3ykf1XxUC0ArqvsglTXBzGrdnx5e/5bm+HeTIhdsFZPY1QIjNUrYPy
qvqfpkKkqZScnUFGDjy9ztKfchHBXfgokCV6eZQz0ItBIM3nNOHTCwFNvoI31UCYp7o4ZMKWgXAS
pllAmLWAmgrXwxMKdTtqUYt4RKrGmGV//gNRBB2AX0zB3xEaGbqWL4Z38bJQuz3JQ/z9SeAhx307
MHpuVhnzPvPPZBK1X+WbcgDFi0+SEbDx1Dv7WAEeGps+rDgFf+pS0bt15D4BPJma3nJG+FXO/a3A
aSlwVp9fiI/RZ949HvVgc7ZVwAZpKhtHsL9nPZIxy8dQoJJClfQAIzRJ5YMDkFa5I+INz2dKceNu
f8NLkmoe+6Uj7OJMTp3qlHGKPZCvxSz0oxZmsXoRlTIbeTOuRxjKXs2Cqs9LKRI5614ATRbZriVm
BOpo59C9NVmZ/Agv9Nf7Q1InuojosCuhfe78+2I9uTGzWQ69Gv/KPK4wIeX+NLKG7lMNprbq3IpW
wH9/iD6bCK5K8Oubtx6hhkzBm2UT6CtfS7+1mUYeoxTtm1M5E7wfmKAFi9Km7sEu2BVOEV+pQrM+
S9JyQcdnWTA9fiu4M0YrFBCvgkWjxWw5V1LeeE6hNQthnpLH9XX9AVuOEN8NerVAa5iiOqzlKBTA
nCXrS1Z67bn0sPy8vO3OuxHAt9s9IlkkT+5JdS8o5D6MZ6OV4BXFwJeP0OniVuS3iWomB0eu6kOD
JuNPRWerQFvi6z2DfuSO57i3Pkx4wA3B9hYiByqH+4rFhSaraQ7pDFvDhyTP9UdKk9tQL19K5IYe
7Mh55TaiTHkxTJOZ7ZuC/M19+2Cp4s+ss3n2a5CUy4wUTziB3dOq/n9JSeHrCJJ50j9HJtlHyuWw
Kb+K4PWZ7HBmGlkh/gHffDXnKIix3sa4oXhBQcaTorWQvs4dhdRYl1IRL8ot6/rXQLQC+MtTQOFM
4RGMinz+i7ig4LNFfWfnVWdKSjqBNw4bBb/fSGb6x8WFyn3duAHB6xDQ6i4+/YnQTfR3bD61Mw8G
g5Bo0a2UNdPrhJbgV/8epqQAdK7t3tKwy5QU/M5lvSYDk9Q2L6PvHzbDpGlr+8R1Mgk2J923jDZl
L9Lr5ytKKFeqFAvi/w5NMGvWlWhGE8ca0frY9swa2Fd4Y46VZBTMqaMMAT96vBtOQrQ2aXlSZvWt
OJZOCHzXstGYppb/QBPnzw7CHThVXgI18505pb43iC+xNkDz263uQM6qVASn+8hWD8XvGzeKfWyk
EF4hUxr3y5mYrnkMHXcW3irGCCnqDnVdZE6nc72lj9GJNC+h1ZQDPATtM9NlaF6ARylJZ1c4yIPN
E4Cf7JAl+Ngq4+9Y+KsgkGshFMu1tXy9aR85P6zCj2fIVY4w9Rpgb9AiFs0qNH7B8XVL31yDSVK5
3H3XGoxLpyxDV2fX41iAIVkvmY3dr+jLQP4uOe//OxCE5F+orbGEjg2QNfLl26RCU5JUj11dDSbA
WuO3jSwlsvoeU4zyy9lcG9P/2/UMGejJrSijiCKqdLl0cPON5hd42Gx+Ft46WbPQPxZM/hbPfxxg
dD/R+b/+mnlfQGb7d4IMawz5vuWlu3wr8sNgROQnB+r9xA2meZC2vc2yZBacCweHjio6tD//Rb/l
WgXzdPnNDENz9eT4SUk8p4yGsoxhBdp7DPsYePBnKGboyu/P8K32dxKQ2yjRwtwLUwEcRVi3vtmf
84sDvsx6ToJ3/b+o/0sLTudt1W+grTkVn/8NHGtlu5n2H7EgiVDavu4UPyX1WquTUNi9E/YL6KZH
OnVlz37Gi1xpI0Rq8UBEe7nXSXS5uNXae9m3QbT+t3cPJMrGlSrF7dzyRmRAkRxSrv81ETQMQjPG
NDuijRvHaZeoJP8OVMUdASy1FElO+AyDyRFFjZ3F6SbXx9J4jZJZYhRtLmmSnm7LS+JX918J2B49
2O3wE3IqtDxqUF7TG2Tfj7XwZyMJsE+alJZpAhjwpU1Vh43UUDmv8Oj51pGHb61dzdgngLpwkSnB
bjgxvbpq9hkZhY5NbsCBnmea/VA2d+pRy5jx67CRCfp5V5GAJFbFez/3sNjWxDl4hXdNToFdweXQ
SpfR5Ao2g8JOmB8SHZkn05Data6cQRgZEfR7tEyIyiPw5Suvu0k+tjhq6DwrNekhQs/3j7L7Gxit
frpgGgdvjtmOI6hDNFog3SDoPA2PVK0MnBsIjrL4ax5p8hUiESUMFZMK0soBT065uszis8tVr96I
dqsE7p7Dm+e7dZaCUliiiEQckZa5TaGU+hA/2a00x1LFIQP3ijVvr/vabotBK+6xLIvaxM9Ao7Pq
OmoRS/hCR/seTGNFpqEmdPNsiGBoNsAzgyzIa/NOLDq46c4IsH1vZs933zUJJdbUBlMDEamv3POS
hznJekrAc6e8TfXpGWyrNwddjzYhn7YQ00S+XDcDJYwJ0ji8z02ttkbTTsjpWg4vhoq+v8DKw/uJ
GoSXwdGjRizBKZnzDJ8KJnt4V2Vku9fGtlsHnYVcwofE+Vwa8oH36yxAXzF3d5Uzb+GcPEHypDHp
iU9/JcMXwJulN1Xbxi7Zw0sGF79xNgK0toSpNK5ato/joj/IaXcgUnpMPbxkb45RVD75jHPSWHB8
KIB+9J7rOajI4Ilp2f+6DBTuTFpL1GrAQy5buWkV9Gkol2vArPkvT42hxVjeau5zCxEyDBKnPlP5
MQs9aDJ2NMFzIZhdQMX45zDVrtTu3d14+nTh/3CxSEhRyTCwh6TK0HObzJ3SnK/VVlc/M5l/IaQk
MfyrR9wFiASGHX6qcwA6fQYIGGnvSHCw9l8Qc/jizeWwUnaNvKHA1TkkjNctUSGpBAh2ejvt9t66
oc/HJRuQWwYvth7OV4F2foN09ubqiIFnHAFuX6z6aVuhsxvKQlBMwhD/DRq7c9+nkJv7+AOz+NXB
Veo9ytL6DXuNvqC2MJyt62HPvW/qibjbYrkDIEKr1UHSCbEoJigdqAaKZ4vazuDsMPPY2EbF0wN2
MtsFue1/88g/UICsWQswX/AdBL2oLfxGDZMcX1M+M6Zuz6WSnQ9VHFL5NgOdDL9hC4qmE7Z6Ktjy
RGbbI95SBULqV/Jm2PKVHpSamEGE+VKn/4yvh9XgIRQjysLaFU+QMmInGu7QTEYEJMRDbUyjn1uS
LG8v99FPn2LtfSVGn18LNwu7JV+WBQGUqBB0NwL1vo33b+S/ZwWhMlWptJSuruvQTEnDqfadO8jn
sUpKqBHDvaXpXcCPD8uUD5Ar5o7AvFuxgjUD2iXU4zUnAemYrfq74YjXRgnYfFO6jKHnmHtu7Zon
9BraXDIUE3dKQwTq3h/PXnG10ZvJnx4Ox1Xgf8Kyq4AuScyX/UlO9EwPqVDdpgw0S7vRusFMTwQr
llJBIT4+WajKNp6E6P+dUjkBfj3Fr2qjukVQNbksrAnfYm5IDt5H1JzAcyJ04WHj/vyc2r1ycVYl
zVR/WCyOiCxgU1ysx/bhQjjN9Lw5/M0BKFechzJIEUUmBrEq9ccbAGG/lK0vZ1EINgJCp8FXqQsX
ocC4Cu2lhFUl98oLtf095MwZJqrO7x7BfakmCR10brQXwTqwkLmkYSt94o/0SvWg10P5PCzp0GEZ
EeHfolPYAORe4oFd5nN+k6qPqiWLYtv4CS4ibsY79TQiipqb8kVTjgXFe0vK+Gn6VU620t2AaFEh
pKwW+eMdYOKUdj07n9u1ITRqPJYTAeNyqE2qLFgWraeWYd8q+EfIATNbWMF3ezbfnJc7rg0quWHt
S0Qi9XqZ7VB+gAAkHU/LcGjnBLlP5TZRvVSTbmdlbUkNm15MSbYrkTHwIPrAUURJGQfr2hTtxDPX
OnWghs862mg7BcL+BpGFOsXscoZArN+fb1Pjywr2Utr3EX0uLzub11Ze+0hfN3kM8ixYDfdyDvah
yW8b7vd89zRddBJI2dKVsYlQmrJYStc7tPcI/Rf8Wfmcw8k0QCqYe6cllBObARWY4haIMRRjqct8
VIsgQu+GuRpgpHn9iGUANZy2g/ETXaVaWuoHxPgCd7gJmDWkPwbtG9VPbFGFXe+qMLcHWOTJUsrQ
ZMbWtbe5KR5l5I9B2SazysI8EavWHs19TdBj0EHt9bbTj+h1kI18omQOzAfgFYXXRSGQv9x7Z8ZW
iT5g1omI8OiS3mvCCnjipik0TE8Kc2pwEGlDiMBNF9jvzEr4ygip0l6TOGRZo/0rS9HZCYiqmZYF
z4alnKj6wBtVuWkmmy94KazbU72y2w0P3U6YF7dUqoXW32LbTqwm3JD6Z01nAutR+H7APXzU5DrR
O/I58kErz0RDuJYr+7ibhBB/6kY2O8glmx5oshcXb+l/klWBMNs0NDeyz0lHlPg4AQIvDatPu+F4
wx7+TSW8Xj3bLn96RPGbPXpCM2a9qKYob9mCiKhpVZvTn2aHkvC8SBrL58LAL5Y+VX9kqrFES5aG
qBybZ4T0kiCr6b1xqhGAQjeujJwVDccSTmxU0c2Xmjn0H/m4IFDqAsvL8JdBY1+rW/Z4yNnlw+rI
JmkHKmeVX/o0jm2gD7efaQLlhkjFE/oPrMBbFOtlvOTDyXP/VK8bqyMuYnFTe0KlR+y5SRL0BQKA
2xpz93eeafr40dQEK+SMxSipY+jBE/7FnSbJLecNX12v6wqDn9awqIDOymBpMjaUkOwJDSh+8uFO
Wyhmpk/fyzIc74zlGLZWjrMC2SzcSkm0AGRS6azbVi7hlePT9DSQpt189JrNmevLLwvEQIM6HNJi
KQu2WhoXcx/WAGtioQufWhSfzdAypBjNVbRplmhYV76VOrVex4QlyFmU+BhwmQkcuDExmpxm/JcD
+pFy3Xs+mETWeoGyzcYpPuLE6SniZht5HMOZqy7OofStRmpKhsj67xatusCO5J7oxE71DGepps3/
Oh/OxU5PuHkv0OemtWSNVmw6RcmFe3t/6BXZDzvc977cDLad2Tttm0lnBHgcKzvTPNAJpFzNwqOk
k+2rrehrgxlCzBoMcPik9Sih96mS9Xzg7hUdMz/mWCwHb9SaUeA31W9tc1S8nDZcMdXyoJ/5X9mJ
hqQmhc+rNTf24vRVrQDRwuYufyt21XRhH/CdcigB8r1+8iuSN0x9AKK0f2aJ7dtEct+8WF0sUiYK
meSHQGOUX0XPI94RQOHRiV8oeWGnnRT4jrYf9K6iehSxwTXi7JLkLFOj3pGavzArTB87YyH8kBUJ
JOpR54f74dDCu+l044m8tc29wGzw0siEYiFXkUGBXN1FZmdqSCAcF+fnxnMbbbsZeSRRzf58ANRG
08ORAjqmXEamAtRcv3HGD/W7XQmbvGTAkJPKHpgt+vrzcbwGPrazwu/cBN6dU+BBoA7fmEkYddDR
uzmrv/wRv/t7ovukV2PFR3wTd15nIGs4lspJKiVuHh6vcAXkcdr001PrvON+soFFpwIbdYWih9Xn
+/kmMOn8yU4wEYD9LEMlOZPfVcSvlN8z1Mnlc1o4Azw977wcgtrCWjRsgeFfLvzz07oi320Eywj0
UyNtyhIC7Oio25xJE1AWKLAqaEd/Wdwmjcqp/pwMAeVrTKFCGXF+IlUJztKbEbtz2ftq6szz5Vk1
9RynmIVvT4PWvqCjC9kO8BPQAaA0cw9BVLNcoM0KgZVoq7DPZe5f60b5qhB/wAXwoTB4tcVexiTe
icaz/bb88drAHMfV7Ap1JkXg5PUauW+/bLiV+wNDWH8cjj63laIFUvzSqPfC6SgIDlxySeK8nge0
5LTLzdMRchUV20+LohMHUpPMIuvfFKzqqh9iZFr63i3TaBu8nQ4ZKQiQe4sxYFoEwKT9SmbWkZnC
AzWMjfD4vxLAxktL6BYD4hNuHHbA/ZUaOkYaiV8V+Xy2BTgCmD8MlDydIayp1XAzt4LJL1HwHBuu
xqcEPKwD0IkRYUukY14kU76FNbnv3T/X+g+hFhtm8V9NBY7kyVErP/cTHBrb/irjRwQllxnE2F0u
5NslaFP09dDkkrqzEeADZic2IokpZJ+hKnazVQ4qnyF8eY+Cy/0g9FCW/zgSOV5zIggVb8Qjp7Cx
WDuX9Qe3RHZrNi6KkTVUqaKVdOKyyLcOHoDsJftK/+6CP5Pfj4qNmMtv4Y5U+2e2UTyN8uqkyw1N
XK5qpDKTkOEpo211+nXQKAlxF9mCSLg9rj91xpcgP3D6fjy3JBAWBxZ6hHTs/2X9VpqoywcBhpZD
nIaglE+XBGacswUM/l/NtPNysqmk2ss9Fm4sh+0at1fclMJaWPcngJy4gEs6AQOogVTEJdPqXq4X
BD/1hxghRm5qZBBBvnxYF4VfmvZ+c85GhWXyVCLMO2mGrg25lopOcFAyM4tszLg/2r54aqaeZP+e
5UDRTTNir5eazWoIc5B9wy5fL+hHoyqYxpej4pn3fAV11Mrs7rLvZ+axJB8KKeG3WsM+SQsW5V4T
r6tNbJHrPbawu2+myo3pgZTrfGBtzetodEq60pUA2XjC4yTPBTL8lPRZUTR9rNCTU1RlD7qnia/E
DDs6wNqfnmy8NkS2HXivrNDrwGz8Wg7dg65cM3MVYaThPnbwdXM3bYTGlyJdqxH3TnoNomZwXeni
VmpshF/d/ficEvpRTPxvVywopHBSpfmuURv4Y+jHHgTLslIO0c1SoPNFfRXE9x6jjuial/7rKB1d
9PoMwZjtC+/frpOu6xXCyBEW8dHO/Ba5KB9+OzmJ/WZWJqijrcOsTy2TjsY3qmylRxOk4B/xteem
yMgxZxkJlQqAyWXPzwX7eUw3W7MlYQY4jZQ3YDBjNnL2QmAx7wFv3vlJcNceyxwt28sAH9RmgvNM
u0rIrl7Ldy8mum4pMBub+mBQ/lbU6r8PGWdZ//P08EFlPLpPf8YDSGunnav/Hr1TuPlANyWUgO1q
mZf+WIn25U1pA8ac+wX/2G+oBdc+/E+Sxibk7d1axAmJ9AFbHIG8FV8nXDaE7xhduoNSnAn+Ggoa
HLgn1QP66JE78yeVhLI3hNMP4gFlYj4OhYd6pQjn5csMbn7c6hLjnpvzemb9xI0PDEeBil1H8T8a
f8g12Epy/ukQRd2JKREnpFxpnns/YcfWIrENExVNxfSbqcvRjJ21j+qJyOK+j79YtwbQd1omRF14
S6NsF5Hktnq+tSt4k+ab2JatiWbhcahJxjcWk3vmImW9/9ljELrDHl5UEtsjKpxz2dOVbD+eLpIW
c896vhKnbod3tk8+oYyVAvYHLJe3AYwEgyTm6DpxlL0tH/vmT0ogvd60EiIjTfphqBGxMSuW7sXb
Tn/Yvz2vA7ceMj4Ia91X+SXy3RxPzPeVt36NHMzvcyI8ai6byv6UAe27zXY1pr7zG0qRZ7dZQhgP
G1svyKKkClIM9Xv7YIkV+g0SfMHiLy8ocPO9b5EO6dLv8LQyMLsCijUywxZElBWD4WOJA1DQOJmH
1x9XyAkJYEk0xM+LVZ/kaldjYT/o3lzfVsF3VubW8E1YzyG5Kh+0+eKdiwQlFpUQOh/7maOflKpP
ZnzYkeTRaQbGLvZMXRq/JZ8iUXrKNxqTqS3Szv93vap1KPeB0IrZoGY8TYOF+8VItS1bvyn4XIxc
6M2lbMRP4YShpdVp6iqWMfFdp6YJ/zNSyS+OsXSwTE5n1R0m5E7hCO8JL41lXFAey78Ro+F7RH3q
24vohgLj0ZdjQ5apu4ln4KGb+iaOLFrpzTwFrP4iy2UyaLwkqQjjIklp8XwQr3Y442XKQ51mhxwV
uRdrUC386XMOoLdoRFz3264+YYlKuKo4jqNWUYx6zmtnkHmOlzelTlmWfgMKihxM9sX8ah96OBLM
yNpEiDcD3QbLYe5ZOPjDNlfkdEUaqwDt7qbUFaCIi1xehRBFnBR360r+FcFD/ljlanqfZxLzndfy
jSzdJe2hipIMafl/wlKNNlmLyAoP00WiWa3HPj1o3ZPZt5ngJaaLdALXtjf/bz2OoeOj+6nDCuHQ
LBusAtDhmJxO8e2MTGpn+P3IVXwoCp5O+EMvqTs7ny1Uyue48FrtkxIHgIBBm9EfyHmNF/eUOlhh
kXkh4LyCyrj+tvOg3svy5WEKqYRry8V63vbhsLeiQO8mB7n0x0WNmfotuLzNC9hCSh89QBSZpVmU
awYlkkGnLbtyVqGLZCfsz1llGzQhvXx3DJZkMjSLtgcVt0c198fmmcdPLWi3ceUPcqeHqy4JwgGI
Clj19m3MVO8OsRghDjt0X1p9YljHA8+hXQSKZuRr3xMEgdtv1+Mqj5eRmOV/szOVodNYRvgzMrON
SmteTsJAYJAG6Hd0lOkq8vQnDcwdqtAZF7jhBHyR1CVgRIT6bjrt6OYkZXKqe+Sl609MWnSpMCCn
8P8s5UEJTMTOklOfvcpNogxeE9D81zQs6sqIHYXSFHzMedC1QArPPrV03jSSUKxly4j1iPwtqlhF
PmBIHVW3WJXYvcUF5tl/rIP/mkW1c5GEcjyrYpf7Zp8v9v19oytSZuLrIY0OKRKOk2JO491oKmky
O/MOghZ5kkcDFakO38YaZw7k6+BGjW6dNBQmU0Ech7wEnrrOVT0gOx4fjydBrtQflmM2N8+gZSP9
7j2mZlpVdGj/z7FgwR0bJAQslfEN1nNjRUI32aTr1pdpdpaR7EME/dmavXaBHXjQf3t66l7Jk66M
DXmsTCvNLQzz6CgME3WW3282ADPa+cE45kbCY+9lbttm+WC3epMUpRT6NZoURCIDSyyHR8Kjh98b
Ve4yqEdQA0XCa24li7jIXHgPtFSxDL4+mAYgUx4LmUVKsBG62jM3wAu0pE2NDR1bRcggzPMvTkss
3uV9zuYWApJgebUF2ajSBkTWGVfMWamQt2wzs4tJKN6U4dfow3dfvxbKos7LAOwMwf4gf3oJ1G62
975kIhgET0xFGDJ7tUbLONBZeK+ovjyue2wGJ23ChLXmt/7nhO8fanyL5Kds24G20BVFRfba8uT3
xA3tebY8Tudipe6cZ9g2X06usvhfBzLsiLVeSgCXVn8IskFyG04L6Aqxa1JXqeyhRoYz1osOgohh
TbgdXEWeqTtGWwGIemCDdvEf3j1O1f9L6tKcEueVGl2ZQV2wWWegQknjKYI2YwxzcWadbEiLvYAg
2eks1tqX944CkdQpRwHD8ZdRNcRkt6l4ijFrcq7pQYAnJYsNJ4dhbrAFtRZTS/F9bVJBKHUlWmcR
Wd1pVxkqjhavhRMNBXc06ryUmHCfEvJMFX6qilZRwWaWEtaS2CirkJPUJsf4k/T+6Hjix7thY3CN
frjswMEcvtn0eG6pJXtgv3yILA1D90YqsecmSn5C0rC9AJkMljBYvRh64NDPoyOfcn3FN+oZPbY8
p0yVzKg8JrnJ3Cnh9A4S6rTOmSYy7B3UV0d4H7xsP/zwHP5RePvb5HN/+z96zh3FL63JXSD11Gq4
kvV4aq18Mvy1o5m3PN0o6KSnogMnbfGA4YTcgJeOpaOFlR7+RgWR6jtmLEj78eR9yYoIB7DhnT97
8OVBRgtGFb4MRfwR0+GS/ybjRNl2+eyVQskVKRDDl3AxmP9/NCMGDx4LL7QaGFWAIpHhqycNCPXw
31k/yGV7Y4eAGL/C0KUNTUQbVDZdqVF9ZduNT4QkLeS7lylWHcw3eW5p63ykTkcDq0emdOa/gK3L
qppImeYbc0Er74g+JEQWni8nCgT1W8Hv6a9U+U4XS1OcBUs1KqdQaaU26BiQFBbRYfdy7tw2YOR9
q2fskiIfTZK0xansvfW6UCCfpMB3csQdtx7gT4linz6o2zrxqRUDj3T5bEg/vimcgmyBVmWrbVdi
OCDLlarCtI3tYpxoyDeyjgAlqH/NdmHJKebn312ZxRa+4oW41kyZ3uB4swlKjEVzCwcn2OwT/EJ8
42cMvzXmrKn9jIUuVq7Gwt+JMhMg4tIhsb82pB6rE1lCE7ZG828gfKgCNNuOlt4MiKXtqeK0bYFW
UDqC7kMMFrn4dlyXHIEGtAylarEFJEwv67lEzzIhNu9E04fFhlLJQzG3rp6BH13wRvVFuVeaobqx
JyUSegCBcmMF6Fd45agmcPYx5PVd8fAD3oWis6KWUbAMzwcPf8rCK3fWNQEKCkQQIFmGuWo+7NOv
OmmvT+Yn2ioPvU2wj+pkmfTv6IhBBjmes1pQ7n5WqqZ0x9DTynavi52iAn7J+RsColgO+1SOBlYj
zsGiG2IrJeJSAwWjD0hcm0A6lsEJTTBXBpixzLtBfdKlyXDle6D4yAc/WX6hNDp87MUsY5aV0f9F
eKDlYA2qyz70g+YLpiU8WwvMGHQEj51hbUJCstoxkMy02J7zI9QlBu7jrLh1hVLmnW58+UAK2C6p
8/Q8jXWoDwUeDQKO1xuQe7AbI+/DYMdFDYGgcSIecgQ7aB5+ic3BSfigrHvENGddHzIfhvXxI4tp
eSBbBCFTSVDSJPwCkg7b6Lc1/dernh0yV+BwF2xHZRIWlsvbZ23+GK4EzKrjRQ6EdNXNvWbvmgQf
5g/PGgAQRApsZV03oLVjSHP6Hdwpzh8ENL4gagG1O1TirJxQNfMgApJyd6h/T62tjifdIwqm+isM
c/DJl+JA4mPNphwjgqBOmIR3xrM9cSWDu7SdAAldiwVt4tJ56c13G4DMMMfZd4ajuaQ9NWhZm/XG
F2iC1gV4F6UfslIRj70T+sO6Vf+S/JzFcnmSRETj8AhQMwmE/X9ZgMsbZFNuGI08Cm1hypHDI6tv
AAxjUq1vlFFUTh2cRLJgVzxK0gr8g6VtVs9n/fXoWas3q8j5lDtVWR3JsxggUlYIXgFEvBKIchAb
0crYMiFZQv5aR1I9Tsdha6vQgvVuM1izO1maftEvFrSrDwPcPFCSMrEf86AvGB6jz1AbtN3Sq4EU
osK94ZSQITzwmMVvichBl+R/ZrEi6P8/ZGwj7W1NxCrlMMijp1IKmr/srOWjpM3MFR0lCglebKf9
ZBvCtOLJU2ZyDwD8lyDZbtX3q0NiVr6q2s/lbO5x0xk8cRj1nwp+o5UsbmZWB4U4e9cGe0KSzvhE
hjZ2WJguUQtn1rq28txJmppOn0TvYhMqKOXAg4D1mPPel8PiAOz2737I90NsbflCbgAeVWvelD6i
Dig+YE2Hkofqqh6sHEc7mmhibC6E7SPNoGc4KlKnWFoSCrFHf9R43LNKgPI6L105LbpnZQrMFUdX
dEK35XZ5azP5P7GvTKjqZgGs7KZJq9DIAb/HCCnkTBnJ/liF8LaxLtnrV4Xtm9hN3nadEsecJjrR
kwuBGpUbEBS3eR4ZpYxeJIoDQx5c9VSVobhAQy9gGbw388ZrtNQb6I8H08ugPjExJtkSD6XjixzP
0zNIbX3kXmO+fORuvm6+qXm1x77objophHuljFj60V1qEkdxQ+PgeHsTGv/bYOnA/Iz7qZvegnXZ
LU8gs2TrOGVnzaWDLZwyClyEEYkiddpvQY4IAC4KkVjYEendUldlLomgSD8ET6KR0qc4KtgTYl8i
rCZuMhV0+zAe+iPIRxN5sMQzkAO4u88n7bu5lXu78KjzcHnHqj+sze4VoXmaqQWRxWfW1kkP7d/y
FvsRNJjKmgiI3SJkrAwEAIypdV0InFs6VeNnHLUQNl89uaK2e1I20PV7vyup36Ez1u1zSuht1Wwr
oYyi4QPMYpYY1ZbdbsdKvXwuXwHFxw8JEhCgV3SKzCZjb0G/ptohpi6liwn120n82lXrI10adElV
qXYsLvn47JzB5zMKJ5gbpZPfhBxXJGEqKwIqeY9ykIukUWPmfAN39w6b2BDJqP+8QZbRIFBtoYsH
T5dD/FZcxdxtpnTJjdi6K6NyaIl2JO3bR7n4bNP0yeEo+7A4TRMeUPQzPHJW/qfGjeB434jYp6Tc
h5pupNnOg8cYVNpIppNJhjGUDJL6Qx/NQzaO/rkX7NGhLTAdZmxi2it3dYcCi786Utk3jdiZP8a1
HAMtlj75dFzH3YIlkzAXeIWlB9vHF7YTnwK/ovABX46SDDVJqytEg7N3gi5SKfgEXher+s+YdpgH
+6mS+XVr9X+EM2+B03GZ5Z7DqrzSKO2zAAFa9L25WZV8ZmboUizHY8s9QEa5MDRti1kVyeYXXRkO
L3Jos9RYcCRCNj0Ddq1FB5RlpcYg/71kaYuQkgXhlcktHtMcniXh/qFbDM08+K0Bqvtxf16NDaLD
6fNsk580tvWYbeAgHrdMaeXSUMHlsPJTZt4osI+SwWKTw4FpOT+dXjvqYBxC4qyagpo7XTi4DElk
G+k+VV72jUwy/GkznuRToyfgRLwqO0eXZOv1dwhdbl+1lUhuerxy0fJcA9W+7C2UGkhpyTQs4DIw
ldnLyq8mWnm4ropGV3ON6W+l7OFKk2NU3L/M2Uo1qe8B52VPA64VL2i5128kcsy1QtgZupMSDetJ
tR3toz4sA0dN1vTaViS56B4ce/s5+F7HG1EUYf/lENAHtihRI3mZH6K+mizmPXrn2EqXI7/qMsHF
KMgbZLburoljxwVokt1Zb/wCAzgfcIb/ItzjCoXZaItzmxjZVrjwu+XyRK/PBrtdoj8I6MKFeTY/
0OuhOuTc2edyBU5THcv/rbHX5K75OmIPOqQb629atbvYhfG8MfUo13P6/Hco+CDTmP586vg5cUM2
Al7XhXX4eiLDAQugIbptpsdnx1RKmjbefBOSo2lzFMfgEB/YS1VDAa8alqyE91pECkB7k+2Mvllp
7RpmARM015WCAVkrN7E4jhvxcxV46Q/4jcfcKmmWtNC8x9iKSh6z7coDNxwpi5iJppJUq60sWhHX
LuruXwz/hm92dA1DkDf83HXOJSmMYEr8tl4jWViK87q9BwX+lKLQ2hS3kOKkOUprphkHcjHcQPg8
6IMnn0nrj5DrzpxL/1CSJ+zj5A87EZ1qCdel9U0McE3mYb/piMI5KchWo9VYtsK5JDDwBG0iMtuC
LEOxHf7xUqSL750gb4/lhtLrDdaYq15RtnqIJku+i8LMKSB9bl/FNvQrC24gkUyW+Xor1JSQEVcV
iDAt1DVOWAfILFHd2Yjoz/Usz1Bfph3T5CZ92k30xB+F3FQugNylomMoBPZoZqrLUHVkIBsZbZzD
XYlTfYswHvycc6g4xOZoa3kcuKMxTF/R8G/kMtlcKcx5z4MxLP5AGNMIOqYXbIdJT0x3UFi5jmux
+ki0szQ0XdmySkv8PaB3oZw/hjO6RhaBQE54kxhZLN/msmPDQCoJejStw4LaDcoUzdU3Fs+KgX25
LhwTwCfbQy9K2QkjJAXAP5GIHsdrX0sB1KZwhTWcYoaRtR8649XQvGKioJfEqFIZ5rNNsTcSrvyH
iv8p9vXDKAcghzOF+kYpES0aMPcCQKGonyJ3DD1Q2cVohoQyQ6pgnPVoKd7xyon/Cvhd1lN9NAs+
nvNdjzHK6UdQhevKmxcxJog2als9VD41rKGfsXgZLsa6KhQ9nowgSw+a2CpauEl6aZ6UtgSVKAeJ
wYD2/jbFXwStBFxPIhBDlxGf6denJWZeLDZPmbBIUJnTGo6Si4vgXnYps83xa5XFaMf0oYRNapPs
Kc1tG94eWmh6b+Big/9pfhkRJNNL9edfi/jHwThAIVi1GypNF5cnjq0Ii+3zvd2jVsy32o7xo+UG
BFyxRote3zNMgpfJgXJHWCt6UF14i4VtPXzbHmoMdpQE1vsXEunFi5HnxabjARKcxVjCIZHstehw
G834XVWiz+qBith75xSTuTmQAIsKMVgq527FyqhdDRCX9giFdastw5RT+PYcG87BeIrzhe1+qc8j
oFwPXyPiyraDx1L6WO4O2ngr/x4qYA/q4qAStGZ/SV2DJiKIyVi3F+K6OrRb1yTVD+5ktwPQEYd+
Mr1/E0YvRci90RmQTSppo+71/ITauq7jAW70yf0jKiE3x5lCgMeDje7oov2SMyQ2idvZIbIEk6Be
annQe01sNnWJ1jMWxTyZHnl0ipQz5KvOIIXpXFtAMHUcxnj+yg6yQF0Te/EmGI9acqPppfvCr0Ln
M0gH0iVkYUXva9MVctXQdZw6kUWq+QzidjFOi6jV2v6XysDiTiOfKlBvLreFpy1axOMIAsm+cFYN
VyQCw19xH8C/j/7yAQr16xKjRj2qe4tdzMTa0Agem6awb0Zg7EY32y/4HeSz49O7NOIdblKxYste
VvEMA4V6V+S7D8VT4Lwx8NI1QrvuY+j5DvB9pUJBmyRUkfPoJodIyP3iZpoeqx5LIPiAl+yssbJV
CfCOSo5GtIUc6hmQtA5z0f8eWTSpEFR1Oh4wpyWTbrcc3pVk4Q5rch3evaidy0qLLfdqyHrPW0QB
KOPkcopBrFJ1FAZd4V2tvubPvPu8puXyC6wWObeQahudVTqcYTPTqdk7/ANIM81DPz0m8m+celf3
ZTbM6aWwA83lV4h6QN0Q6wIXuVbgCk/zQs4Rj72j7F5Fel4d34/6j29qT31fsiN8bbCAUB2C44qR
2oUDIUzGqZQcX5jeJZ72QahiT2tYwVUySUZK6CBj5aKvdsFmpE+ObG4OCDOG9dCXo5OkU1qN0d9n
vpfEJPrRuFUSddnlm5mb2JQocbOvlGIr8kvmF824WLAEyElR2QxKfHO0KYQBZo2YCER+OGFc3mbA
wfbSVVO6kfIv17vg51gOJXOi2vmG9jmyvC4st7lFPjZJjlAFbvpZrQ/m8bN9OOIXO2fjN3bNx3X6
I6c+ZU3an5HGL4I/ioGJmHYeeWaoxcgSNCPMj8V1S0jB+XNC/bGyHReauhgxFdZ0eaagsD89G4xO
0IJRtxZ08ZdGuaEjxemkafh5BGeS7TXF0ON46dSiyZIQYWIR8Nz83jQm1VFeLIJ2bAuBzcqMittd
u9/CPtMFLV93jDZLih/ShGUim1jaxCqSHENo69oxsR8G5AYfM+CxHU2JfFDAHAP9Kc3GcCyZkYuW
9vwnPHfSe9ucIcFe77PTKLTYXVg7F440htmJMkSh7OGR9RzUydHVx5zY4e0jjQlJPV/5WJwKAYIE
ehvuYeCETR+wT6AtIEJEIz6oTe5qVjwtFO9iIHXaYTFSkHD3dr+Ko+68L4qg0wB4kFCBhqPs9Fyz
lgFdpZUVSAja6D8fhJnvKD97qYzGIorIkTrrP0+rHr0DKjwyGuLvS0Z/au2gA2AHpSretucKX2Cy
+hcC41URnZzq3Aabt4Dfx0BO9hZiGz4uoOJDYhjBajqoBSRrzYKGkpZ7UybgXsqeh2YFZhsnb5T3
p2g+tTQmzYOxi9uIfZX39svD4KTAuiWDTJPnZoMiRx/dsYF5nzH6oNk2rVt8JNaGbBNJbs419x0z
fwZQe0Kek75+Q+1NphOyTwD4YijvAf5OZxIzXVjCib/3t0xkaq+aiO7dRJuhVWCkb3PoLfDVO1RW
6NqhTfvclQ3abQgI7C5EoBijIpC0tEV9c5vaKFY0jvFSie24WEVQ+Zynx+ATYhBsDZ+N8jhl/x2n
CajU6xQsZQuIID72Gqqh+8nmMv90U4uEVLaX1ySHi9mnFQDw51nrKeo+RHTM5Hbsh4f3Egm3jtW6
NwJVvnCCIVIJ4K4JzTr3pnH/+8C0jgE6NLTbJsZTR+/FMCKDINXKhC9WHMYc7at1kPU0m16qgXgE
rEBHD0LB77EN7AZF1goOzd+Q0tccjTem5Ng/mM8XZfclZxWeJMV/UWASjyrb54ARh5eBsT+Scceu
1N+FrgK0Brv6qtYw2LUa/ZQiWrIdFVhPYUNt5TU9N8+d6pRGC5pWdci3wfYuCdYrObkgbLS3yV4p
03X52Pxc3QQyBcfm9IsZShVqyzb/5K50bl5iJad1tYvPnW8p9hCDtytPpJsSrouDtY66zrmbWqQd
aOBse60dOjeAW04+n4wv8QhUEEqfKESeDCbGQWmxc8AEQ9T7t129CdtHCrkvKs3mh1jN4zU0y1hj
7i+jLj1s/P7tT2hf331NC0GF/Wg5FcdUjBlggryCGOgRUbb6+hQ8pmHju6kg+/Dj9AIIw2WdPeha
8byqLVYXUQ66+UopbpJx0zZ2DNPunakOiAR/+xvu3XTGdliz5hmRAxc4tNVE5q74wbeVMzwb1gc3
lW9XAD5XuMi8IOYq+bQdAZam05LIpMRWm/ZFjtNNIHm4dSm7nGMbkVpAdWLTk7jlavOjsCoabguk
3S8wUFJPU7lVqzk0+xCsCPuiLQQRkio87FqSGcFQpRZ0otjdEwNleMNXCcL9lcoQLkazwR9Dzr+T
VBwkSU5sm62hSmLorzeYvTaqAx8PBinJspmFV/wXoCGkO9djiQ7W3vsAjQrQo8SDWF20l3XpNq9T
gA8g9a+P+rfGOQWo1BQzq7vUI4cF+XnLUZJp/OXbWG/sthlgRYBQofBrsA62lRbmfbxQinjoX4LZ
0n7eZqnsca9v4K09MyRwSw9shMU3xrBaceEuQX8c6EcqAZJjq8I+rEFKQDx1ynBBMWsrrZQzhOhX
JU2FjIRfRMggCcW0svOjxZIogv7ycL/5cim1ws5sQI1Y2lLR9KULu/VQ5iGCNj6qdhLn+4EMl/oA
l5q0I635dE0SJ4Xmtbn8SrQTEV2z83Q9PNJswgBoQYp0kVkz22Isf6a2aCcL2wfgtmowv3VSFNwu
28urd6kJJK83pXfqJNZIwiz/YzM3O3mSvVOEAXYCWg9GVClwwcR+4tpZe6abyjnPhwjjlvPIxLv9
SXT1izHPmTsVlmYz4RgJQl4G7MchJTRDY5ARXfBL767miw6fOOXQP86udpWRuvL5ToeR3dicu3OI
rPHcjBvRgWT/jEfh1XTWgyWUjtOjytXsEsauFA09p7JqFDGEwB5jrlhMzJCUm72FSnYBjBjEeeby
jpwmGLCecjkqM//KHYatnNUM6A16wmCi5z8pZ14jm+/ET+Szjm7KawdBtYMeDBRWCXzEuXfCbTIz
lXE+h9uWAsCI7q/yDrlKsaxwoHDlJM/LJIMz3xlNOXWMcuQLy3ZKlQKQk+DHBF1XeZGL3rv72VeV
hjslfEAj8BfSJIBnYUjgV0qzxQuTMsxtclXXQ+ZivsrYXUMVFH9UGsytmGwRjAOK4LHiT4WFaMu+
rxh1HWlJNGZxG17qGIv9+ToYY4GJICG3+kZQ5sgTdd9rlN5vSIj5Dh8cwJthAIlLKJ/cvHN1hU5f
FFBEegya6+ONY0ESLiooZezON+x+GeYSICHxyOoSKeL2iv+IWE7XhD4bexu/4lIlMG9UFsX+RLEq
+BYKdH9CyW3L/rQze2rPGooBZMOLIhN31JDfOiq5IEPs3rTt7Th/iYCRbzNo7LD6Us/r25ko4Irj
QUWLu0UVlkDHf+aRrVxuyCy70ZKdnSofnMAdzU2eowXO4vyAJw/foxY8eP/XWbcaexct3R1//pS8
d6Z6ZW3a9O0QRxk4T4bnXJw6oU5kMh/BKAaklTf9ruowZLVwuBvnZgF3XFwjR2LdBNqA9WKJkxwu
KXCKDAO63xCYwLQe4vk8Oy0qe696fN22Dw5JGHJB7u56s8aZSd96Hcp4LrHNFVs3FEh6BQ+Ov9lm
A6U+SI0CX+dcTeK8SjONU5L6/nDL8/AAwrWk9QZp3WfcqMvXvCz1L56Tj6FmT1q4XexPrYldfDHH
8MACHOcWtytj3Glx58vKb9sniyFzXj1b8wjI6WoB+2cPLgYMmKbvQxl6rCQQ/8YjysEIWkqC2VhZ
/hqi+j/C+lD2S78KinxH0khPTY/UsGriIkyfEq3x9B5iFbR0neT4Slf5hkgW6fDM1alMNlcr5NFh
+hSRW0Ivt+F7W+Mq4x0gh0cvt4i4jmhQTNg5Ez025QGYCsMQiXTIrk7s8ggkY9ZoaWwzJV1derIu
jwJcE24X4MjSK8ZFfYYOd6qfVQBRpQEa7BsQbrKJrYymnWy72AGsjjoS9jyS/Y3ZssSs4OBgKaBL
5b2BF7Ek7d1j504+OzbKbeUpuAZoS439/3oruM1R2mYIoBZmonZKNWyQHp/hxrdTU7t0iV9mLmeA
re76/9QbfahDWEtCiKtgl88yWMK+dxKLfpLIqsSz8pr+X1GlRFatCP7axwsvX8S6V7f5kDlqtEI8
9KfN0lnZ/YZUBnoSJYEGAKoujmquzCuLdSI+g16s6TvKggHxoqB6rYfcM7Q06tGNC/x5eO4UkUmD
Gj9FNKgycdoIPtVkviuXoSU49xBqdeGPRtGkKHOxKnuicTLUU4KS+CUhxTFVmhdg/PfM0jv62nVP
JXgbE60YgS8gvnD0htUV2Ts5FPyEw46gff8uWtHKpCxNxIlk3kSalrGnfAkjtHJSjOvA4uYn478/
dxvDYtDcS6HvKgXJmhn0WpPF1M8SHbDGc7P7P6/HPheLhJWFz7vETVxowTvvWdL6tB7Epso6RJjL
Xy1pOvIVSSCl20mIQcp80o2T/wXd1RDtYXlv8ial4ESfqn+aWZwjtQX0DB3UcR1m8nmfM+yZjbDC
QSODwUc5gtlEbs99qfBNecSXx+LBs72MoqsEVbM2OmbrwPKX8dgdh3P8ztaSWsSvv3cf/PJ4ifu9
93JeU08WadC9jruSKGXZ3I5sY1sKuBUJT/bTc1wHSpRcg5PoxkRu78ESGEQ+CtPUntuJ3Jt/kpdX
kszJSZ1pJQrDJqHjWoq05F6gN4KpHnFq9+gVSG4aK/80er6qaQsQk7fH8Oi53AgxlMTU5ZHwXRwG
TkttxdOhWVQmY35+auqHg0HMnfJq/tiEq8ohVYQJo9uD1D4hEatilXKU5ud/HGjnXZZXrNUW6lfD
8kIxNhzktRV52Xz6lNVI+QaaLvXtWswkJWGW2Iwf0jo1VNqPFUxYQV6MPvqQUy2EEvuJswZkf/Gr
ghpifPdKr+7+58pW5KdUpCX0XxmrMDnBwET7dz6dQ0n6hneYUHZqvF92LWc4xtBuUqxrML/xi5mJ
Atp+RLt63QM3is0sqFydkFR7imoGCYjmAjPgI4mU2dlf/GM7QebemFqG/XBhBCtUJkUBMNFaCE6n
VL/b4SxCdQm5GCg4DhgFCGfy8/zvRL8O3sL9ltBmlUs6h0A23MSzHv35y2SWTKp5Jtt2vglc+bJZ
Tv9KGGbHYKkDrpjbDrc/6S5oW4Slnkqi3RpHoYI5JxNn0CKHacItcCCvVZAjMBKxMtu/4WIiS3cd
Y90ko65kaG/H9ByIMxgPIXII+cZ/Ha6A6/VlhuBJReekKBbhCx+vb1yNCKcJ/ApqHuVvDZikcaIn
G+5IFeg178ljOmq7N+kh1L/l38vGFtLSVk+1FLhm6m4QqR8hEL1Gu0K2fsyBf0oxg6w4YTuJ1DZn
wX1pj2P/Uv4SvUVTGa6qpVVQ2tG5eP3Qdv3yMxMiprrsSD5rw3e2MbZ3xUMCL37yqkLl5rhPmr8k
mJymEg4cyxWC8hV4cZ5Y9yp+iHVSfXJsxuvNeqF0wuXrxMoFLAgPNGb2FIwCLSqHtU4HQjlDrsub
bfB2S6GQLNKE3w2ZGptwiUQIvCnv3FWQ8svV+RbT3OFup5O3TUNakH+d6jcBF4yP0b4oPRwrFw5z
XdS9XRXHqpKODHHXY+p91FXbOIoDO4ZOp2c/sVcvhv2ffIhhxxykGUET2IIXHEYzKg89ge0ZPL5w
XbBPW9vBl6wGLP5Wq7B6Mtg5oJ0+P9smznVVzH4bi1BEo2p+zXhjhkgWEcow+eQMi1Hk34r+fEFj
nXFWkYQFa1X22YuM/Sl9Lior8HWpqrlseq5MLnhDoYVc2RJKcS+TE5hMN7w/A1XfZMVE4ZNS1Z3J
n6U2torkcAC2IV+DxUZCLv6jroBDvYZUQyEBjubjMFrDtshUttN07BI5kLfVuIH2laZ8XaumcfA2
Hkw6JY1WhXawaJu/H9UN/rcE4vAK29OFc4TfyMdJafKN3S9omDE9jXMuH1ZnU25YvZYc9qn5VFHi
Kgf14bSMwtxP6l2MJLEr4G4RkUVKK9UAfIQR9nw36rq3QNyTPY0El2+ldn2lEGQnK0FwKJ1G3SU+
uz8CiHeUGX4p+b2UQaRdhRtaoGEOhXeu8rgO0d/JWvsXHkFHSwR4TU+pUhjXToihyYHqt/4qIUJo
tJdQJ7QLF6J/p/LvUUtKQeHN5PDV8s1eVglSoQO5yBMqOoAI5Qkb/9wJcDxdihJ9k4KsmCV6ozQi
nfkFs0Kkgj3Wtcp5z+zMf9SeGCbY5fHX4kJTaoVbmAw+xQ5mwh36Vk7HzJQ1vRjFiYumuPWEhVMZ
f7ZvZQCJAvEzNr2j+MQZ0Cz9py8n5jaJC37gzk389hAotjMnETKocyanC4B31Z4mgmTPRQe1gRXy
ZVrMlS1zhxF8T5/O2IUhuVwbDTCUkXjYMk8NPpfFVp9CA/nPkY5TC3fBgFkBvjGE9LWSUKIYqR31
ZVNHND8qVnDrciOa4GxjEq5Ma+SxxVz+EURWObiDi1tzJw8A/3D5zHbgAlctVIYEt+bsnIQnRxwZ
HHbW3Y5VWsYQU/CBXD5ZENlWUwHW8dGGjiCmFV9Ab7M17N/YB5AUfxeVpqaC7oZNUqe38Z/UtJG+
9swMhRoDZWduDRYIjozJ98XKgtTge4g6AfmONEKydGFhEjYL6skzNezGFZaBKqDFz6RamrppwHei
xKsHaUZn8OR0Bp0XP/2m8qtRZutUQ5YHT0V0EpY18MyxQRdl+UK5MdnIZ3xCYsosjHEjNZR6qn57
XL6GEIlqo9way+Cw3Cqf742eZnOZs2Ch3RetFgmXoZ5ejEwsb2FSpRjUBYfOREN6YvJvLtzCkfyo
Kosl3kX1bpG12HVbcWFCZkF2uxDzbJiyk4UoduHw0yFX+Q3WUAm+DOhGoeLI5JJlYMYjqVG7Af8z
myRxMKVdLLQeTJV4eO8Gs92UM7nWPjO3ixrxVI74WVHjtPIb0XXL1L++7x/dzVE/2jovmU5CrEaZ
m4/P9/43aqNPIcKma/5jwBr3VqOj3ZChyKpQk6XF8fqxhIt6ClErdBMZKbSjFz/N5tHPed5+Zc1s
4dC6Af79FsEmUu0jybHg9HRSFDMLPyAdZkdTFe7Y9/JzF8CQLqS9D6V3Y/QCuaY10sMbE/OPOtY7
u0AkF9OgWyq/E7rGJKbOSvz+zsEtEVEyKdGxc2DOQOGobBPN/MBddRCwsOCCPDH8KbzH3C4eYVxx
33q5LtBbUoTvXk4Jti+MgQ8PbS+djeRt5H30EIFvqieCw59nCCQP5gnqNrTg7YVW5AK2KDATItEC
FGlFqbzK7ocR1hgnDNNFbZ8pN7AJ3JivthTK/1pmJ5VjBHYR1lfy2oyGlwPyGXlov7V5GLvN5BZS
WHuOUVUoENasOZ88B8BovkJmloctbcxElck518uNz1u1QUz5afmcDyxZyNwvKKKLhnDhX6++cLNX
/e/VSVVETjVfp3rrm8d8ewHtuhK1C4YRIPmOqRw2CX3b2BTBcwo1QLIYirXFQT0kdrbFOT8X6qsM
kuf39kYFzXRx+U3mqDEZJf5Szts+jo/4TOQUlz3UgOb97B8hjwL9cke8HtTlHmt1in4ULYd/SX8g
Utuf+G5qvZXzTSeQnNcjYAQefHF0eixCEohPkj7cmW7CP7q6UcwYTTaMbgTCpyx+wBp99WNLAmPd
gbiQWfFhW6pXU3DzCUOLaNl9hug7aLmhJ+6wo8bnqnUfg5sq8CfOm88u5wV28h0hmyeHk8UQ8+WF
7wWHMDBf3JOmxD9wKBkuGIGhSiHe3QBkFHfWCTbo/L58BKoBOgkG/HIUWCfq8wW4P+vk0FKFAiTF
c50M5N/HM8tHWM0BYz/QuG28rclNrntsBy7VLMdPiWzremQ+M3c0/2J3qFxLWc1kRUPqJ8hRLOI5
+QMTPrnG/16zdJLRO2mvKYI0D2gCgdvxaVYN2q06WnPz0UK6v/FnEyw6LLgCizJ0EIJ8FfWe4npT
wvsXUF5hFs3Erq5GY8AxEvj70f50t5rPkcwd9dIpV5kI/rvm/3S2Jr0p3m2A5s/cE7LUjf8M1cF0
76q5uNUK2VpWQqLoHdRDdWZ1u9vweU1OPYfRGAnsANzEGg/6JmxVdSD55+1FkgUEpw1HaX9bndUl
e1fNObnv0S1wpkvFXogpZePXFPeQlTVPaoXew6ZBQ3C0LHrobXGWfjxgBa98smFJetW/wadBiOAw
u5RvpQgZXF88UWwR/GVVcS4kdJvAuSXOvYY2Y4fezhs2OHHl622t44y1iWuhwNOYctifCuywuJkK
3BuG8d4ss/bBHG63f+PVNl/mthwGECzjjgUVKLPV6S3YhyPdZSPI4bHU/jhJczY7FG23UgDIKFUQ
2ng6iZ0ud/xaYHxd4fl0unWJvARKgX3nscUZuQZSypfpGtk/kDjvClGzxwrqfV/C9XSfkp9lmk/g
wqwbGlr9j8NaqKRulyEIqekV/OhHIdQ/1inDd2NShin9NihHJkD8EeRADGzKTU7DtR3kVVZyZXQc
sTmtCDtrS343sVKB9z6TPTODmO+dVkf8gowR2ymE4HFMVGELAkxOfvY12MujrtMcjGROvVYHdWq8
453rJAfdtDPM623OkJ4p8n9WE8xgyK33ue+hXcFZ9+NZ9+yIzQHW3qTNh9py0Xg/IhnG14c822Cn
H0dRLPuMBzkVvC4Kbig++GGRmoKwNwRxCvxQY3LtmsxEfSNUutXzUtVgbOv5aLm+qRRnDRJ2adu7
/YWToEwogYBMt1nZ2eEbRGn7BmMXkteA4BTNt18pEKb1LVPcDPq0xnEotqZDO9m2omQeJzCRVjh7
9Hb+XEk6uF/V+i1VhUZa6LT8Zefphd7j6UP4CwzZQvHz+WYiBTTMiSxf9RclErGBBZGQSgJn+d/w
3O8XppuDGYgyvVIpto31KBH+NlrBOIg2cEO2a0YdoLxLjaJdg2iHwkTbMvZFuVp5v/eqIAL3DOxm
MmIq/l10oTZ+bpZKSoLAg3urDHefgWRAXLnFREypyRdg+m/npn61V8+2i1i4v1w16Iz+bXmAbbNg
NohRWT0khxxAb7PybYXqUxOJgcfrLFyTJe6PzPizy4ePJ9NR6N1oAsSLNM8/NBUwTYNRHX1XKwLY
pxLPYOCkMX6nY3cfmg0nkKDIb6I3cTPH41VfGvQWXmIVUoiLczAnNq1O3JYKB7vPydD24Qw7Glq7
mgFOK78gnjH9Ii67DLaKrmyObIrtFmWTcAcudNSoQXB6gbjNYVc5oNhHQSHLeud7QkSLKCS99AZx
yWwqtORsDnsNYjEsHg8R9eK8MgT4x0xqq2WBeY+NnqPxikRLyYHPm6Aty5R3waILcNXMuGUTMHlD
MLsIg2pLaM4rIDxdlKRD2Bsmnngcs/q4aL8Ju9f20kDQwllhjDgU77wsl89dnkydalnngx56ySdL
8u5V0b/bN9zRz84Je5O/s8dik/Hd9RkyzqX6xaqvdWo3wdeTZidxX2qajOYbnMYIZLcj8geHdWy7
27kluazhkUWfmsxYu4nWmt3cKt/5sXOZVCa2NlpejVNfdZQY6/qy/zBmfsNaNowHCm+8HI82exLm
F2SNwxo6/YHXFONYCPxfKHci+wfIPZFJCzA5NeDD627fFzt0J1liy5IbJFKWiVl5jqfdlqQyHd4E
RmK7Y/FtcqXFg86yestoWncGteLJB1+C+Ufg4K0NMBRGuXNnBXRQjJPRZNQ880yIcYJy4OqTXGRS
KzDi4WaC+StTAEb1O5v0v2QCtEyymOXLaYvpbUJhTDmXP3AkwXB+jaz4yTIuBoFvXVTty7nPDNim
sdSqjZ82CwQoavGg6CVLGQTDNWBMSz1rRhyOWHwdXyl5QL80JT7Bxix0C3UMveLqooWUMO/Ul9te
QWvFxjn6UDwHfUKzs+kjPCDgxaTR++aBPK2ejJ4SboZGWrHrnkaNu8rTSkQ6wAK1NeQcNjWInWow
8yZXXqyeHvLRbrzbjhhV5XH9KYNhrBhMZm6IVQ6FU85ONUpxVUKs9HhUhPv9BbxviL4iVPP2rNlQ
4XzXL04rPVKbO3Ppb5qpTnepuM6zJdIsAUyHxNdOaB2nzWyoBXUDaltqG+rzIY6GQlt9Dr1qJh3m
H5lGZU98zXmndjUSjLi1yYVj8qh1w6jVjM/fMdltsANfF75+6m6Krg1dF4Se3ZGbA20WULRPYMcN
PW3rw4zQZMFJvZiy+g7kvISOiAwU1QqkPbMwoB6sunkO+MmKCLUuHl22COFQv3t3ICskIThOyVEr
CRe81E8JwYWOa4/8Lh7ZXB9h4uTFl/tA7rRbKlDPYiPcvgaFcy2gG6rsFwnsRnB21CTSoxccmoY7
rkr7PDbS9yMzDhy3KLFv58GFzUKaCZEYEHyUoPL+ZIPmxFxn4aT2uan0lFrA7Bi9Q6SMNzl/Ntbs
swhdp3Rg6QxzRo4DY/naWA2re66Unh+A8LWZGILSubJtrZWqLSAuaIB/lACMakRl6twgr7YAzAbL
eKdCpQAQQ4dg3A7nw9LWH22EdTQ0L2qCrav1DLAed2WZucfOVBXmyLP0lSoDFwMY0mPvd2Y2bb8t
CHFoAiDtAbW4d4BMgydPt3blWAo/TthMO7bL2XpijHHA3RHf319atdjpv5qHG+r3r2mRMmJoKPK1
EDwfb+W9dg3JVQKco3W51E7ZugN0RIMzVwFSAlMqWkz7KIPXgiNx9WJ85cPO6ISo6cOIsvkCDDTm
6ZwtDYED8PMwVpdUY9rRzalaKIFjLRRWmq5tOLPu/9KidL2uZGWIfzqP9rf9djpIuFEcimZ20IDz
EE1txj2drZ7xoffGNwCaXxzTMWEn7m3bsMChu9nlZGjFx9VPDMuQOvyFILFKBLT9BktNNtpgXgc2
WkHV2qDHqiMX8SVZTOciSW4J9VoP7vErlOUKlpEYM3vZrKzxGb6YnAP1IhJbP0EqDKfkwAAElgAs
3wbuIqqckWSUu8MdmU+Wvw5u7cTkqyEgssTdJQf2tYcmsuKpN/urZ9z9tmkD9uWLeI3lP1X2UBih
MzPhAag/fjIEx5Gx1D8w7AmyoHM1EV0ASIlJesazWI0/KNWXsRuVmVz2tmUwl2nrhL/1h8wgEF2J
MJjeq9BogMbHD+7SS9237JfX+OpeGFyS1iNp+oRoWDEacVrlt5zmIDDnkm2OLxvuKkV7NJ+BCulz
EOPLrkKT1+deEiyQ19BRgoxE10QMC8PBp2hgdfeFURk0A2IgRzYg71Tq911JSvK0XxUO68uGzGZD
nkZVBvTR26EYp9ciQTIO89dSgO0bVMhFObX2c/Xr5OMPMN8yd1hISwO49azNT2D7/50BYqF0Pn7r
xExzx5bWkgEPOedh0bZHvpFIw/8DwUkvsKo7R+vNDmcIloHV7u0VoWa+rqxfGMPuZ2iz8tkbUmdA
X8UeLCHgOewxGnkMDBgFJgbNFxu9bXpnQNLXWSxjmwo+3HEfdhI/y3loTXKLBtiEJfTM7/bX3qE3
TpbESNOsTTmq6K2hHl5caZxL5YnG83x8uLLpnm75KoV90GzFDF5Y6JvadPrFqcuYk1eT+2ZZ1y9O
0Po2c8T0ZqDKu3tUSb1J4aIixZ2+wJi9uQrCwBL+gz21gsGP1T6ky9EiYWGhS4tEbQiYhI5IyEQP
UNxUK1MN77mX5t45ydSEkD/4o81FpN+oysNLcrnpx0G3h8axTvAoa8rUl/vMZ3zfozESQJ7+O863
3bUzdA/Sn6dQiNiVb+AXqP/X2/THHEtvHGRo7DfAcEQXRTkRUsjb+ef1aSBRFdM9OQZ056k3ZWXv
8W1SPQKWrGcudO7GUHb84ijKhqVmrjgeAVWy+GCZr9DOtzQ5l4RUiohes8Y+te2wmlMS6lKq+xmj
b8p2W1LtXKwJXQgJudxXZuK2tNuBajV+k+I6Tk5batlpcOkGZz27D5bRIxUBmeNvnenVQUfuaaEu
vGiDaKRcWroxV4uun5PoVpBiucMWc890IWjMY4JgIHp5xZGmH6C8CGB+uq4HoLuHp4vlk1t3WxLF
Xn0azhFisKpNMz19IYkIQgT4g9KvE9HpoejY53U2NWFCPOtRdSPlPyYADEaVNJFI6ZyoA6/5PPqm
J7zCC8lTXWMKD684td2ssmXr1zoQpz1aHxXpkpclHhNwMQgygPjPOyM0jrIgk+lbOXOyMUn4EGGM
oBjSVcu0sUBf7Bm8+JhuaS3XJ2lgEdgmrwZE8rMDkC64rmbg0EEs6Jv+e8MAeW6F2Y/u0qaeD3Zv
MOjyRaeqBXCJ4Z9+lrhnN6J1fFVbisZjdK6mj9LfBxNOUxMCbZkZYB0nSdJBY2eNXGm+c1A4Pk6g
ydapwqhFEChGr599N/S/bkuwHw78tveNk+2Py47TzQBLC/TjHHPnoqXKVhVqLSzny/RkEOFJGuxC
Ds99yERei9DcqGIg+MUNhrmYMpTO+5HeO5HITLUahMKcP1pQFIQhQFuYQHG6gtQfBJTCLAFkPXNU
nxPAJKmp0GQIwD6sDLWlMRpBcuN+Z0hWZQMWzTe/LPzaCy/vFmj+4MHSW1YIYWamrOrasIB1DiWY
t2FRMcE2lcrUJ+wxK5igys71VE9mNcrKEw5ZDFG7woPIW9hEm3HIDLK8LQVaM7VDmRsOzmnxh+UX
nfXB4xAr+XR+RQ0yif6xVqqhAe1hB3TfZc/TjZvNDUQv6C9f3qDSoTx8/PBVBt+6SW2ZdGs2tc0g
SL5yuzYpb6V6ICWO0SX/wTvHqlj0UStTz94iReXx7E930ve0PqvUvolp67gIXI8zrzvDYx/NNl0U
bov81GYySBri8AU3XWa8eUrDkj4gvpnWiWD06IQyDeIrSWYAF7ynie8BuPLjDsIVkXMDZW8wbNDi
2zdLCl+N8B6TlVnwNXn83ouA8gucp4L2JGsJHlgWpXIlIGaPl1UKU001oEtWb+r4B30AacmuaWiz
YyDqPBAtYTcyNuk1Iz2fmSR4kk2/YrGRihqIFiN94ouFUSRjKip38waIaIptaCU38dvFbSQNNGUS
r1wzop5+b9aiyRBjDgbN7uZRZSsRFxiu+Mbgzf3v9KhN2k6Q3IFej7DD0JsQ+JCOWxfPmHNcuVpC
HvV8GVTmVy467kFuZQKpwrc2EL4Qw79fnJf6lfUuLeCFSidwwskG6o6pKKeZxp2k+L3bCSMJx47Q
Egv9UA9p1Y0YVgbdsilkzLBJGhGuXlMybNSyiPB7K9CvpzRiN7Edy1ha3bma5hIZhexnba1lT8Zl
LftKvfgQsYN7u4ui6J62nY+2m/xTyAjQRavL4ObHM72MYGTY831zmJo5JJnAVK0IOXFgL/kIfqcb
xprlAPMMxLjnBSzeC38VG11XQAEajMoBR7MUANaXxfAqT0oiOVLEIrQPz6W+uXmswCIfejd11mVQ
DyNG3To0Nn10vZmEu0+dI16sL2USNelFkhccRR9cQt8v0EX/R2eDb38JXMJIMDsa3Yn4J/uOGS3I
xpHWTPNwsqjvlbX8IgThclKxtONkvsiEKYSreytq3OfOtPEsCSElME+in2lPqWR7j6v2/o9r1M9B
4p6+GuTqAd+iW0RIMj4fOGrXC8hRMijtBSdqAmELss/tvQn+cCz+sJ/TYc63w83ytXq0Oo5c55RX
N2NryUP5ujsWMq8fQZmPjkkQMEpB+dr1bRzoIOf2Gvq1/VtM7zPK2DBogLH4OmsOXsLvNEh8kvw+
dQgzpmu+YB7gn7P7O/Bn6XKKINDPfdqLlW6QAOC2WcOO1FuobBP76EmRgkN0Q/Xd6ILdGjfFetpg
ANmJVIM2vA9luoieOZ7uBIwYQoaKTzSGHYIDP54uUYU8FLlNKyikrPxz35RMi5D9BFOs54P4bPmQ
/E3L/stXcSd47NRwbzgtH/7Y91y9ECwYPG5dGoAirgHJd66z6UpJZL7ZfDfT6X2UEct4hZbArgeU
wZc2iCUJ74PGll8dZxLRtpNb0Wc7IilukKQMjqG3HzvqsPFGR6fo/1MEwKrsHv/CL9xTmkr50o6p
uPGpMStGxuD/Ogv6vBEyrREEM355GIl8HcRJ7anUYKItUGAIFHdpVvcERAzjTuVlUQnOWdlUVOOK
eT3TtBa7YUuQCQNmSZRqRSbGnx/3f9NMRDXDyp43mZH9fDCg2mHOSmxC3lfmYXWmLaUgKP3rkDKJ
MgBAhnxXDnBcz9oCS62hUm2kiGiJG05AczhXZ6CW9VOVNUAQ+7DrUPiV73m57QIVcS7qSxzr+qK/
rCIG7WDeiC4v9n4+sjt/Lyvll8XNGoZJ9VRZ4nsrKMtWM3nihEbwE1Tbjhpgw19kd9jKVTvlc2eY
JxfmFGAXvyOgRT1clBDOQN1L/TLU1JyKRm3ImbEDnBvwwSIa3WyjJ7HvrEMUqExPN1TdSUSC8le0
4iYBBYHMxqc7ySrARGqiiybmQh9cs+g6SgALJtK0Ua1Q76utrbQ8d+AlLYRFoY9KFRGm5Ssa6RSZ
oEP607cV6bvN+Zjr3D8QddKacuaAxNw+qROgHye1L0UH7P5DSfWimMNB7mdfHbroN3w3x79elYlI
aWMD7+jpFKzhCZX0MjYXk0ye7otYiK7ggHfa5mF9Yvct+oiR+2pwk1qlKkoUAjhR25lsvYUONRbl
qompid6Ce2j1VU/afb6fBBYR3gTUoyW6UuvwS6Z46UZoDHipXoKoBToqkk2H0bByXogmZ7iG6e0d
mZbPJX/OL3GPESHLf+PWZGMcUCMmz/YwXiyqtt0alMxnOp6JyQv4bWaP2w17RlYdEYqNZowMaLiQ
HhHlfHeCeDUiRN7tf8dHDJwqXkH119n8ZwrS5yjAcAvPb+J8xhkFi2jr3rXmb16TTuDS+9nRA4t+
duim5QEFLaPnGUb6xFiPBVc/SFGUTM6TSKkBObJvIdABkfVi55gHHwmDhUeQKhRHZO4noBKX4eZY
H7BKJcqoYZw0D5fLqhn36sEmsXGYirIZ7YcQS4SItom3fdd2IYYGBZXmkVLVGTr0bOAXzFOkTSKl
CVbs11pu7t8Pky9xOXp+7K/JecgHYIZpmtjWT7WH0EF1trvkQ1+DVG4kEqmnZ+CmzP8LYTb7x7sC
OnfSV9zHDQjjaCAptTTl+c0Msa5xS2L/zqPhL0418GTduQOP+QpaLNCR2uBSQ0e22i2Gwm9y3FMx
YewvdPWRm21TPPLGTp8En+OO+rLNJr2xDA7Kwj35zFvIgvajFuze4n0ebsizSirSCl/cwsMI2Egf
0q76CLsb+jtuRMuwP/roPzZ0zf1fj4GxV1rgNBjXjF/rmty3ZXZUwTTpQ0gSYB5FSLbd9PdY85Ic
pa0IXkWb+X1mqx+ErNUNMnWQIK9JXLkj8FpKbX6uaCKXi8aPyHNqDJ+QsFyMtvKRlp5x9B1NHt8y
onPnHkfjLgaJaOuwppoI2l7FPAPWg5uFCyRtuJzq7Zy6bMVXDD0i80nWpwuS9VPV/AVuKWLscerP
rSi21FEVvUsY9NfqfZvHmzVs/+CgFMA/Xj8XFsLvf5ng1lRyBuGUoOtq9p7y2dRI9vCXochcp3+n
PWSP4e7N5gMbHvxJ0H7+t+tIR19Y3v4tfaY4r2V2Cz705QHWUZAGz4GFRRCOVBb4Ja402D2D+TMt
mWGGSWBzudB+KiiqFiqG2X/0t6S33iGsE9515an9rG57Aj7Vi7z6wR/2k5sb4H7vaQKDJHJ09fmo
I/tf5SdfGFNE+q5y7/iFeIyBT3iCiisdVajtjOGOn+OrDPVxKh+vXCBQTL/ytEYxcV1Z7HQFW0ZP
SEy0L6XOdcSVgb256mEl8Qp0FMj3j/ToCsZYHGvKoVaE2SeKsUtrW6HWZjYYxlHenEVV8iLjb0CD
PYg4ZwFDKplW5jc4F40HS/9KIyqwUGxK9+Wyy+yWih9N0ycXLfsal24FPoVIqW2Y8hTrUlP9qSzr
5lYSAhzA7NJur9AQv9bpFYrMawc2klECFJLydxYYmKy2ONowJxQZz38UVIpmxipIiJZfb3Ej+txY
XhVTl9rWugu4HZGY0My1LnnvhpBiCQTQ2FICyzPtou4DfX6S//wHFqtL7hPCJGfg3uWXrmU3keMi
gXwf0iAkrszo/sw1IlvAexAfM2Ug9oYjhS9plYA43oR5hjmlwRntpbK8YLogRgigLD4rySf6VKdI
6uKvo73aLF3a0b4alb5ZDeA1EzffSPweWuMQXWqKka+mpgyraQt53tLhdDuAd7qyUfXh8gE/pfLH
BjkBNC11B4lcz5MIhLxKx3AJz+N+yzA38Tj9KTUVvaoZJUkn/tFH7rbdbmSk7/060fBs+5/HONMv
Gh3NTnrNc+DPWQfRQrtQADkp563ID3V/3GMahnOXRpt5jtFJBh46YfRdi3BiivUuMDtzzUZIaeyh
fxHUVDPmZ01YMgC74vOdbPzvaGJHwIwVxdSundUqQ324ol22KUtYRbGg1HmpraN4PafyJFmAdQhe
Zpe5LVHpLL5ORD4VmU+rKgwExdYZULimQKsbqoDn5LMKOx1TZScEKPRwC6R3LVRkKbZ4gPlZZi8B
Ra5L5wRCg7nAR0bptMeEvflx2RX3ck/VKWUnLTz9xHm2JjElqKbHkrmpmGzMj/oqCMtO8BscpB2x
LuCs+V8Z5oHVp6jOeD7yejSLTnpUt3ZNCK5XueAKwnOSQoJrlrwLAYuyEEYUGAX64Czyhf4rv96u
jC5BerR8hZ96O+pM4yUM+zBwaSiy8nEOzFx3u8H1TNYRLe6K4SXZFkoG7U4a1iin5rRgJg/h25iF
IUEsiZ0kGW5fa0vtEIQj8gFIFHwvcZNC17Hpow5juNik/orabjS3vxr98WHRXACAPr0Xn/5HTt1l
3imszQo6EmWnoYZUgk043zj4n5yFcNyGclgx+/YW5gCJUo8cBR7XvqsMf4QKUWmnh6Ag/nMVSzth
bRpnl7q6/i8gRt7WwH6/ENGqvcVEN7Soc+MwU63Tfbf+0U4GMiF0DVjGcIYg9Xv9XUdSv1eK6ew8
kGS4A4D9CvdjcKPFPHzHAcQKHE7jS6LNPPlIHoA5TxLuOEpXmKw8KIhggc2L0q0wWcnxK/ZT1/U7
jALv4DgWOZ3dNe9S4JucFAipxwrop83U20PpWbYTMz0n8R1lZYS8iiqzcFxVOUuK9vXwHu8fIXLg
8w7fXjFyNbpAYZVRxfZXzwC5cHceeo1pAL/ca2oO+UasO0rk91KTUqjlOT7i9G9iYqNxJpIxQkIw
g/jkI4jKmVqzhsIXXmWfufL38oIpkY6LjkEDnb+93C3g+O5MjVD+DRzg2hlkNMvp4B11Lp8wu9e4
JUNxPJ16bfTFEIMiE+VlbDhakXVen7BkrPAc1r7f7ppqBrdqJzACCnYQ961Fsn5gcYXkRhi9dBRb
IzC22/n6b3hNADbPBfzGOtfXO0ZrTJgSc/leEQedlPhfWJEGnqIiHHXEBYux4xzt4/wE/fjvrKvf
zBJZ0rVJc7tLn14KwikS2a9W9m1NB0PGFjw1+Nv4TZV/8uiQXO2b1RPvZqq407yJ+BAChJBm48KE
IONjl6zAiBU4EkAb0VnKno9BuoJeuEjeWJWPJTPEbO3jXFs469hBubGzyYwaL9Q1YLj6P32+9CQV
vTqXY6sprv4JwtZiMsiwCAPzKeWRn8sbem4nUKcWMED0R/p6VDTjB/v/0F3iIE6CBQjhuA63lNPZ
+1KLwl5J0qRbfQ221Sf3UQSyiPzqModKHJayqr58DFYH0BVmV9XwW5HD8QIW97PZ0lRd5bPs+UN4
qu11ktwnG+TFMlOk2saCdhiwOcEnDWZh3g9LliV2Tf+Z4MWQEpwVKd8lUaSYYJRut/zoKPPYZG/C
XFppcTl4h4xddkEhHJHkfkICJe+PVdmNNaeJgCUWVNoRM4SFCWeq+PugjD5BO2rhnloWxrsQAWZ5
5ksMptxPYTnsKGlB3QWcxeaqKiQtSfGNf3yu2d1w4h1ntLBQzfKf2oix4VJf3AMhTB6Vn85hNVrZ
M/pcM+LFXs1FzaTvwwN9vTxPY6vxlqK78UFI9pA1Y6Tjbg5CbrxI9qqx/iZt6I+Em1dlEyGbe8Hq
zJifQrYKohMzAY//QG1WlJ4xMNpe4i5hRudSHWF2tIIef5fB6i+Pgnfc3kkVbHtv5m6P7mjyV7Ix
FbqB1oWKq93CGxUUi9H4fkJtbFiFn778GChHVVQ2invmGxouDsZVoMPNqJPYANgvzNUKmWMtJGRH
8INFjHRq73SkjuPv+mYdy6DIGh+8hZX12BEYrNuSJBhV5GEjfO6zSY/lTpuILvy3v8iitUypdGGv
R1MGpAEXkpJ2QPWoPlJtjgHpf+XaZggkZxo7dbPbzzw2skvG0C57S+McS6NRO/XeyP7UdeBj5zLg
ato+69OdOrBGGj+/3IQuF1PubanS78+w5oPTJHxCCgqOsHM6lMNQp/+dZStIzu5M16vmaxcDHmlh
Hj68rcd5CyJAYLN0/qEFuMuTPsV9oCMoM8tts7KBdLiEoTN4sjuWZT7qkydcl04YeIyvUZ9RmzTl
aJlAjW/Ow708z0XAH1ytLT0qCw15LOBgJQ2Nm9Sb9gAQOl+0I9NwWIBC+aXSl6Us7sDfB0ScPSTN
QIC8bMKPF5LUAbWjwGpDRvy42Vo1aBmyeeXnCKcdw6WxF6R+EjBdaiwTan+HS63r3XePJ8gfQpUg
sfMScF2ebCLU5dCyyUl1vGi2IEv1obbkF1gSKAcmJQxDL/9RhaL+qfoMk5fnZEzmjj1w45O/YTWV
nOOaUd4TeufexbNaeIowqarXBRhgV+nGCc2n3V+zfZgKEB/bRKDeWXdtRh+B5UmU08HMsHPC/qka
nmV4NxoC596vGsfcpdKVU5KrlJvx0+mqLzYAjrnwkBc7ArkcmRSdQfh0EAP8xj+hxY3p2JcZDlZC
rxXAj6WBdWdINOvUgwN/OQ0hYsu4g8B35coFe5vZb3y33XCfZCE7yer5dCpJ3tHsIi8RF9kg66H8
GohCVFadVU81myiSi1Si5d4WlLNXzT3aoR/cctl9884YmwQ+MQKXsFnNREMRHompcb2H8IoV6pc+
vLM1k6dg2A1jptIH9aCij1BWLH/oUCAPVV+r8fnCfc4js34yZlke2V6PX/nxteShPDv87seGklT8
Qe54UoxLOBhW9HGo2qk8ptKgGteU89+9NPgbft3j6fCkZj1UERi7Yh/LAclPfZ9RhHffHTaY3mU/
0UqitOYjrolFXcQdstVXt7jfrsG2N82vw/b8JaNJarsTxkJuCssBFPfWSmw+LckVBb7JI5VZvick
7eR40EwQFTYOpYxVpFS1gokK76ArTM0n2aE0q2oLW8K1wEgHd2fbnE386LaJrxLdRo+Yn55cLLhE
gQdOZNFDk9jO/P41KeZk2ns5wHFFQaBALpR99TYd3CuAVgcBtC5wuQ42sMNeaE9bVNAqYkDY0mIv
5ONAPariNLCrXCuYDU8kgpFm/qRnNUTaVP56lZNBjtQSvJVx/RYCYjc7fCFF80Qoolf+sHcLBx3u
F3S3MpRFDNoGSo6jY1TSNDCDw+J61ScAoiL0D+qWLUwz+Ma0BHyKkbZSM/dv4yDazNWD/QSM+eYt
pjKC5MZU2Jd2aKV8c3YPV0pOTOU8yNKm72icMarPeEyovi/WOnpiyCEvyQGWzIQu5pBKEpgit71k
In+m+v576HTgwfknxV9fMtV+tZZiqij88FaM64OoIEbJNbWfpos0PY+lR9ljpWtBz2mwgUbGcn2I
VJmiu+ItAIchWazQ3sULG5nMiyTMpsjb5ZEHRaoVLbFoyGZ5KWKKYq7FEEKnTTenpKG4l5WlpD95
EbEH1UnlFJ4WxvlrkXmlpw9LPD2QC+siVX7jsxNlBrb2g7zonpAyyxlcxgfpCZ7YehSZp/hkDxsz
RbQHJGFewuH09VQzNf5mdl5Ajo5JbRG/F2hQKGzDhVi5UUq8BZDLrTVYgNmDFcSiP578LUWJbpSz
ENhWlXx28TZQi2dK8tQl3qHm0qxEGDNMjm0deZs3yNfhEgyO+jctimiBfe12FhIOHULfHL+ZqhL8
CSQ/YneS7uZQsejL4boYx4XA/5RLZDLCVVpLSHWmxClrMrvq32/HPQZhZcVoC1TKkqBAJNesjH6K
EvbDi37NlUsoEyQ7sS7ryS2IASwKxhXJRAmn8/mlfDmiP5tgBbZZ/cm+FyJdEj31ZzGasF3kBECn
MhQPdxsaxfxgFoUswzJtuyQgoao2TOG3Mprd4KDenumYNkdu76LLFsiIFQuCe+jn1e4tHvblgeHM
6N4X956b8pZ4vqyi6o/Bkr+ifcrPtpj8EfqGi4Z99wZK/rdVDPvc0vOcvpoM9UIQCfA60+Nn15Mr
tjCxepRPpr2m97VSW+aF1/fzA+b2MJ6Cd7o7s+JN/NZH8rjzsUPVsX7vrTbZRRxMOQGf3Dp53d0u
T+FrFYwQlUwum7TifPDYPTprzH0WlY/rkbY0RzNaBqYwpNQeW7DtUaxg7Xxdv5LXzKTiGlIN6Uq2
/59+DGlqS8aTZK9fPl+BTEVE9rhnbPLD9H92wPg8GncFhIq0AS3Zy8H69R4gB9dsXrAGua+6JeO9
YZU1o4foujZJ7BZRI0IolLXLDXeD6QVDNFNhs96y23WgD1EeKN7qQw3bCDl10FDjN8L2/14vQdJ+
1WgyGeSXM+4D4oGlPqRPq/Io3wwPiF8yJrrvS9CNdmPlaEkwAuX5VarDLpy9D4PllsAqY4BQd1fL
ocpqZonAvJHWARjniuleaz0n6qw1nAXrkpsPcp3V5P6OfPRuRSvBN2kVmRYmd5dvYKN/SwMguf2v
Hdu5p7uIKvn2EKlY8GiR6vbMe/0/Jw81TTLpfcDWtvY4i1ZxRnaX1CEaePzFBeIEPRnGuYSZwIyJ
zZq0Om/UtmRF7Qo5VR3X/1jJiek0BKaHsGLBUKxsF/SX/NIsYwCljaHnNcSjxV1alvOcT3CWQMCU
K8rwNW37Ep/GZatJnoYcaS6llsNsM36gm6rpf9Eiiqtj0f9hGjS0DPWX+aZdbdpCuypwCfxFCXtd
IdcZ7D5yHEnu8JD0alZ7CkmwNIu+9/87fEIr4+DM9Rl2nwnb+W0cOcwDGqpdAGqufWLEvXOJGjXU
ehH8ygpE2YG9u0rgAODB4y/F1iNrXHJAB2Ft5ZR6JvQardwk4MyGwx7DJCVXC6ePtc5qIXGlUx96
TAjTvT8KocFSJ5eXNA9PSKy1zUwszoX5Kb81SvIfvM4Xrnlxs0buksWZDPaHjGgqDmilavhYP9KC
lJnTwJsWI1X+gUenfSOdxUiUb/+AD2kkQwsS2fSOuv7XMjHtN2nAPxW+WDDkyIQ/EoDJeMA++v2p
SkLHBdxXWaWYBrnddvO0eOllt2p87eU77WnBLMc1h7c7SuStUKJVzpKmJcqcSmOo43x0f3hRCd1b
4iGIzTD46X5jtoJAsfKB+oxr4BVqMwSRGG/CFQCp0Fh7jaHKHTiXv+ycUV7O//5Fg40eS9fiqQqN
B4VCNFJeyDzOS7M8NaHwD/hGgBom7rvhZP9ZgCRbGlxcRQL3Dm7j/AJuM0IqFKDWpB3oWQOQFM4M
/qG+cs1TxRhJ9rxZhN5mIx5SEOncyYRn5Y+Sq4I9joXzMowvKQAti9jnXrjFNJUWUJ4dJ40aRDJM
pnpaGzBOql7bdc8GhA6HHUHShMuN8UHHv6GSTb+eie/M1fyNJ/gQrZ/wzJXKkxy3DqR3BdZLgHax
+lmv4JU46PbXUtLtZ1PQcthenm4HkOB3fHByB01ZH4fPwPRL14lN35g+66l2v0H/mIhK/BHRWGZT
5ixapAzEEGR3fPf98yaBFL+ym/zIjkamB/ArElo9LRmdoH7AqK6kbWDZP36p4bIU4AgAbdgzsCQK
8uBTkD24RZi625LQGqeHkJyEAHaQXZ4J4TyKAb/FnbbjN5ccSTkARqVHdiaSPkoZLMNnYJLOJpHr
fyolUEt61oMLPqmstIVl4B3OZ/D2B911m6D7wzmO1tSo/gn1d2EoOPrXuCACSYGDEh3cZhk9vs+5
aQAp8b0ucJZl6l5KqK5AfXJj+zTLEK8yYzhF27mtQu7BoeMZV/TTOU0nA4/huf7HdlpSEOd+Uaqh
ZcBfDRvjObF0KxJA+R8fcgc4wEkO+xUH5ctEqRGpYMXCvBOKGGwGtuR9qzfrEa1awQnkAQhc5Wrf
OAO+IvraaG6IphhnH6chAPZcb68NCVSQDgdtC2uU1zZyg48DZefzwRSKhBlnDSbSPy1j8QPHEaOA
CF7S4abEs/hIY56CBOyZ8KXJWxqtMOtRKY9I9HB7ESJKN3HfOZS9IaUEbUWKhLnX4Q8tDv8m5UCl
T/xj2sool71WpxjwxQh24PG9A20M2NDonjlrgGoMSxbKK1PYRMa7zfxePYZDVfZlpHvFSXgnjd1V
N099zoE/S1GBfdwOxei8ZTv93YmqINNj7e98xjACQ08LSb7QclMe145DeNSy8ksxnKa7aDHThc8i
Gojw98jLlFkRb65Y25cf7I3tCr6FjR+0ZZ2RiF9wGozHdBg5kyOUTAi1xhq7pBxTwbtHhirz+InV
EkZLkqp1VpE8OY6m7Hs9ii15W2xFCh496rdib9mSJxejj1baFm++Vv1RAB9Mx7vZVE8g3ek1WFUN
MASs4+rUZ0T4qDlrOFF8L9AaJHN6YD87+rOKFE0hroUXhEHz/xqrDefhX8CuPdH+X115iq0Z2hnp
8sWttXHXSXxXrEtdhzh9aOBENykDwy8AAPS7t/B28X2K2buA0hGJR2AJ4G7m1tARAEoxdfuBy5K+
i1EjgqIeEU6oK8HtYIIY7y5c10XuIX4gMwGdd8XbiGoPz2B1VY0RL9Pv28gqy1OxnsyfD+3o6FEV
+CULuhAYES33M2HNuJ+hnRX+dF0JYYPc3JkwcYZHbInUSFUV0JxKFKDglXngYfWcn6XMm06UItdd
tgfKK3Ex5ZzIRPaAQxn6zy5TvXy5cSbWLLMLVO5xru7lLLUIt/7VRDwNJleESyqFRRYpolX0tMhh
jgTL/X2m9fRnhjiawRZTNXs+HAm/ngF4MHAKmnIvBuixt8SfClGnUiXFZzKMmmXjP9tz6cKf3uOH
+p4KHDmyqHEXk8QQpNXAnYvPK8j4FTk40dJ+wSiTf2PnlEj8iGRrRHAXluNOcwR7C5+C2X3wTAxw
GLwCH6oSFq1hfHJeHJ5YmnwfRNF0X/Q8tlw8IoVkg5EcumBjWoOR/IVG8gcWL6c8AX6/GHEDHYxX
L42o1tLR8Z1prCLF34hwqdvFasd6iSpYvjIEtWKhMpb2h7BjV+snLRyJNa/HYe+Ccuc28KYoNIOZ
vq/TeHOR+oy/aCcd4MGR0Dp3g9fnvd2NI21gDKglySAG7KTySkniITWGimsAzEaMNaDvFGrx4Ejv
IoWMTc4/FpZuNa13Ds3pTleEAI7Yl9f6CbPYQKFduTX/zwSJ4Ke+sChDdDy1F9fOG7+w3ck6lJXx
0sdwY8LOMzbOoXq6LENzAdOtycyznoF40MSxqeZ86+C3Q1/2EIDwejg/dt3ryu4wfjsgwEDvs5FT
nARDNP11JNezRAICI12ny65HMNGl5Fe9+/WN2UfnF04PF5xMW+e6SCKqiMlwkGlxeBBR6bX45bvL
aN5uxD6kJ7Pf34+xDY/MqzsYmi9VNvA/bxWfIP1Xkgi3s1KSIB160yQzntpfJPt0xlUKZYvbHqPk
QnpX8oqj+7Kv+YA02Xhg0QU4Vf+VExFkjCxw9nGaLnErQ4t/9EXv3FEq9m7HntAmdOmb5iRg9ALQ
5EQEo4hhPHSfxSVH2tcbgWngGqEiEFDlFmZft0TtTd0rywdb7E4+vKDRWvlaAc8HW1BaVr/5LSnd
9NjIQFVw8PzOi+is2+bmArvr82B9LPz5WbmKpt2TbJgaT5tJorkrvJmmP1foQGjv5zgbr4pUNRqA
QmyNqCtTOysFs4CPrbMTW14sHNwe8ZcmAuW0w/JFHAdJhVB12K+3UZ3l6uPmS3SAgLgtORasnQyf
offpMaO7yemRimxReJ84RatTGt+yYEvMznioUv1ul+xQ31zwjWdowPhfp466aP9u8H3ggRIoE+IT
OGqVHVJ4KPGmMXHDgXSYHqxFyTuVJFeJnFsJiwEIb7PACnr9NXFkW4NIoqtjLNgJ4VQsY61InttD
X2mz8kbcRG78rrQuX6D/z5DZbgEw23JzhBggZ4meAyL/PrvbzD1YR4dHCRWtjxoRbryuENuyoDf5
/Om9eFj92dUf1ObuE2tNwx0U1cAZo+0pmZtP3en9n+d+Rh5qynermXslrsEXQGM2q/ozxNe7NjIw
SlUREdCYu0vTGwQOIzoHXQf3mpFsUjjZOpOqWhpR9QAXoxqrdb9Dbqip3VI9C7Sgn9qDBMMqhHK7
ZkztFYHsA9FtPqQChPi4+jS7UmIaxF3lD6P5V+gE3dFAZ9Af2OK6X/t/FfgYTt8DYoKDgrcCNih5
kF/AoS/PUPzSCDzX7w000F4vtZEKDtMKSxg3Ms0yIhIqR0j5i6xz/LdNximssoqESkkgJqad4Tg3
mJoQTVnJvxbyw6e8oee3r11EJrOtlqzrthJ7GByouYeTSNIlX8iSdp3fwHTtMZm5QzZ4x0uO2Nwa
osxURa8j+JB00XcqeZ5RzNY+z95rIz3yZr0Au2CTYM4SDwfH44s29UDgFbc35+YUFsTj7HuO+EX4
2oYd3/yt5LE+E05JOf1xym+NWeVOlJxKv/sD9YI3apmIjUjBb/p9rhT5ADK1PQWgQF/pdCHDzESG
SVq5U5G51QmFjiWLYCdSp8KNOkoDew+ie1s4lenX3DfHJuV/NOdKwArb3eHIBpmLTyZu+Lrwx8Wf
TmAXU8FKorX1TsAe6BkocpEm29U3hirIVI8TKZDv7OK13lHn9XZ/t2V20IEtXak2oclPtTOeDT/Y
O1ujLdK6VZPOVJ6Qbcya7kXw2nxWIHEIGmEnPPrQ3//g8KXdmJ0hKHjqJl2ZGlcSbz9nENZKMI74
Hn28bExQN3xa3eSeNVM/MLSggRC88mHtd6IHZblPKPomsem8B05GYt0vHYote+hJ5sydCF3RfOaP
hYvBEp86uaj6wgoiMYXKM4tRThwh3IrfOB/0A0v+Hfqo3CAgGRdBOpm1kodjqKcPD/3h8ZddTbac
RCl0JeGoEMGCXrCSgNrbaruLWuXbUxFAzW988QvHY5Ftx2+pXWJCibw5+gXeKvIQshKyP8njegb/
lO9YoBtAT4PmV+2vG9JIv/nQX2UODRANXMRq4vqZB93vjP1Q7yjKsWr55031iyMp8qwN/yRQRntd
/tryZjXQpFvOh4D8X+mc7D034CnitDmFIneuk6ZktTptf9nD6E0WKFUS2lKgfwHsWN+hrovI/GYk
LznzMRYLqOWeL2AZ/J0kfYjSPNYXN/eiN5aPbJKvTyLFxQ4MxU6+iXNiZkVt7yWfzTk8Ux0RjTBq
6mMsKK+zkYoPg4iU//LoQ9SOgM28r2JS0XQu5o01xmPFsfdUDzANZuTi3OP9/eNCaNF8OW5hDWCu
MEfj1ax7S7KZ5HRX8dn77/V9MBtiedqgCza7TMROlnSoSUxjAl/VefxVOc51OGqbJryMNcc5ke9z
HlT9wrzPZCNK/n3bJnjGhVWoZYV49g8Z6uWB3BAZehNXMA0i0xKHHZLZpqY91S1/kxF+Uwwm1b6l
EovA9ILwFOli4xG5kzhxHQMBGRCOC7kIGeNmjGAzO5HdGmGaNAQx1ndAislpfHot8GOcr3nJHk0A
IOW81UT3NqsTmldwxQvIAZ4CstFXM9viQIPi7MHkoVYmYnXL1xJVVq9ycDOrTNFz8iNIThSveluu
dStmqYJjPN+XHxdEGeQTG2itWxIUIPOB0yuRtLEqTwPCzAwitH8yBi6e3dHi/r3ifJCWVZV8vtAu
U7JWVyhuEDm5dRRaWm8uo1+XUbQbWHuNPjxNg4NIDd1O5kmdm/KHmFa2nb2Og656oErbQupI0CM3
NPpa9Us0vYJnfOJJur22kupSgyADIX/MBwag032oteZT9SLKAhlodV1janJhmT7SFUasSTFVCzz4
S5KAq9jPp9ltYFBCD9DCdbIB/DhLJhSg4oAyLmLnXC/i2AnIzoIxwYUH7cf1Q9LHLf6mvCIRjpVU
MMqdDZCG/1lqCu6YVbOtevfQEPE1Q0ZMVcZccYC/oBJYpg6+R7mOox3M1/t+6/ghpF3sw1x5+q+5
wkEvX0h+IGZvIuZBnJKXHGH4wIrpXLBJaouE95avnjlJrL6sQ1OAc23PAxl9FrGWyD+PZXEJH1Qw
W2c9LeiS7wyW6o4ZRGs/LSUBpeA51MvykEYwjhj8THPsU0wlc4w3T2v39UDRjP//GWvPZhmeSgqT
Q8TZWY2wrV2jjJZCq9CikwdCo4xyRtcYzUsrBGfnS2V3b5Dbj4c11TVIJC/kN3Wwg+5EZ0Vh+xEw
5dNn9yT3Jlk33UblqogVGBx2ZichXdMUksEhSa3wxMF4ltGNmuVOnQsOuqRFTSI5KTCobgZ4XOu0
5EAJHh/hcFgO6Mb7v3hcaKSU2R0V8541WbTc7qQgnmn+eW1i3j8qha47+vLzvm5GCjnpqmo5a+r5
gQTE9EmL0wESeE9wFxHWo1x8AzxJJeBSOENUs89klefb0RdKe/pamqQTQXt4O3q2tDLAp1jHoKgy
QfV5kysH3Hve1rbtsBmmbdmOU/JiPz4VMPogf13lYmqFKU/tcPzdXXJcT8g860/4iZ0tf+jhCuhW
N5N1KEe9p0QJu3ZYeZWx3gMTyXYm7ivGc2Ye5vguKhG1Fgcsx8trT2/bRm0aJL7oMy7FdjW+UXbs
kVSA4dIXZPbu/5nTvImT2eGFA0KSy76t936HD2VFjV6VZx0uxP6RhV+CKd6td3UyFl9ZI86Du2x8
bedn7AYHy22dYl3GfHwXFDk/0QjAJi5p0s1QixI21zOJdEBa9gvAlK7DoNkge74uivxDqOffNdEB
fxJ3xkg7FQSgDMZEe7wT2Ibhq4WyyPUWyMu/Bz5IxBgyEFEvaEX0rkYe/dHXEUgoFIx2WY+l9k0I
R9/saONc8wvEqhjYb28oDh53AHXbxTO671rTUCji0YWuInobf6adtS9wh9KIy1qEZ9RFrObexhn9
oUm4RkyEn2tGd8T8Hj5ZQ7u6ziJw40nHw5ihzDpv2/RjGhrJOS4/452wh0I9nUKPnf2H0wiQFw05
G3Tc6d1/n22xZxps3e/QBUajZfUghKehrzAzeLza+fxqrfSBw/W7I7nnJ0lp4f3bMiwzvpiTIUwH
ck2x5nO30lQjkFzO4jgLAdyXTVVjq1D0d9wQcQghxm2Xq/L61+jQfx3Ui4JfloeLgCWWcd+LAUNG
ndk6dwdmhX34RnKjVauAG9iu/mGFOz0xhSyHJBhL28qWc4vJvggNyBUjTcsapsVFgACdR5fHy920
4OcipS0v/jDVt0HgABf/26iWpYNDII7SOuFZv4CmwbTBbgCGCnMf3Fn6In0eJE3r66k5fQ+QTpxG
+ZLsB6/nQRUAccnPuD30k7fzwn5zt+02DTKn0H+6jz8wLFvNpGmiKVLG6Jt4ksYLHFnhZaiXsG8Q
8Zg3ztbblEH0Ak/VAsq+CgQ5mN/Fu40vriG8CEour4e3d1TrdieRCYYC7LRXqjpc0aQqdEzOOgro
EKpcZdT9FdL5DwzpdGTdwBZsQQCUsQgCyWngAciKX4sQKSRsO04IEx5lCfoPOzi8SRsU4PSIdV7y
56ZstVb7Df4B61bQBm0usMwt0shjtvqrA1rr1C3Dq+vfyLiwPbXqITiHxqF/f5ZNZiKgeMqIzXyE
pibM3JwwTy0H5KQ2ufJGRZqYOfIV8/Y+GXL0bfnm3rlha+fx7IldNxsidX0PspwdZrZK4/oa0/5a
6bshqDEzPwxTCQEuLuAhJuiZBLs2SdXZxlIRQTsJBHPP2K3UYx8ycHNmgtMMzmj/4rq/e8Sg4p3u
rRmsvJTfJTKnfhM9GiQBkqjzKzW5UOKVmX1a/xQ3CqDD7jDIkMrgPdMkuqWZOPip735WmgLZlPtc
ZY37JeZQGcnY3oLj8bxxNUpQtfU2S8qtA2Ltg8pPGIOsG1krvkKTVaBbdq/gCh4G2jVQolAH4JQn
Kt2X0GORhqJnaLltSVC/SG4vJmBnk0JF0KIpr099JIlpuDDoErU8DSqt+8ATv5BeE4qg6FPX6t16
fjEDouxrUMe9wENWu5bfEFlOgjvlVkLidyncZVUghkTM9S40ZijLnwkoUSsRYKPMNGR0TJ5x9r1q
kBaZTP0j3aq+ZQN+MpMnsT7V0yD3PLi11asPIZBcdb7CrNRkO7IhdDuUcn92+atBNWEU3sHO+8B9
2dmEWSpbBB2EdSSs8OqJ5J+0QnUdJN7YrdJ654STawdyd33/2JuUfjl5nqNs+Q8gxNVBFVcrquRV
LohUX4k1faLqTmEe6Q9c7pLJNaxIpsp99f6Tc2YhIGiIzh6biuO6GmsaWf1xPv46GzYMvh+a9Mb4
ezyF4ZIVxh27gP6bL2/mRlajmHevPvkJbOa+3G6duRlB6vxImcCOSSaj7xEvJdpj9rlYQomatMOC
LJ+CjwpckL2F1zUGkAsQMHynuS75XrfTBWxFijJrRTSj52CroaVHpSohFSEZW5ZbXTTabl8m+wUY
+aCxBAUt/P8df9pxcdvv1Mt4/SZmSeMQqwj4hykScGZyy5igxLttfJqogkItdtPvAMCKOCkE/TrU
vMQJAXh4XRrRqJNYS/eFW+Dw7UMSN6La9WJBybCj2pHBG56m2bSVHxqrXMUop8Z3c21aT4bwM2NZ
saYfT6VhzallkbObbQnsVN4tuYbpOBQ4oMqZwplOOw2afC7vgUSGwww5F3yCjwAiixaMNKUWdaLD
JXeiH88etu/Lb2YZ/EHjgWRMKSUA4jjl6Jqzlf3ORqigyHwprh6rAXbzJZi2+L9ksVwKobb5tRoF
jd07/oADdRinEkvwMqxprDUTXOb5XDip2tuXUBObd7m35CInxS2K1snlZbwWCX4eTsoQ0Js4RQbC
ksM3BBsew/NpW3h5a4GymW80reXyN+u4DJ/b5s2Sj34J5jjdumcDxUtkvCv35GquYKi25q7hv6Eg
vIinyxou03cZNaFHNvianIkS8BfqLSBbvDE1fOURUnjdCRfiwu+VuZBRcWuaRW8PHgnJc0VJQhMU
qbTT7DvGFd0Vmk0BrCjsWF7sprPpmKUuUyxf9/+IQ1mEnw/0/JpRccDDJUiWqPfLZzzNsyXFnMko
ldTfrDOaWWzOVc/QDFBUhkrjWgkt9scJan1q72wAUVSpiI+BnrWJAhg7iAXMa8FL6SENPMaZ51fx
0hqFw0SDL0TVDTir4kV1nmpf0qPM0fuf5/3f1abiNOM4aRq5CTDnAuhVqOUJxED/d96/TDR2HUwD
/EhF9qJGECiXanZkDFr+nQAWdgeGQbTMO537/2zW0CANXuFFnPYRVln+uaJzBgqdGoqwaEVqa6yO
VzDt57vHL9O350ngvL/Nhcaeq2xcD0+ZCGsybRyKAhsoUq0c3cqd4UQaINvOZZ2SMLDmp6WlgJnd
R5QCTkkTN8cPdzE9SIMypoYpTwMaFX3aayAmPno6iHt6R9TkHzHUSVNzKvTHaYsY8+3EnvCCGEK7
ahxpwmVK1bFC4RLVYViOGInoP1lFOE95/4TFf5Fr4r4BMfZadstHUvGvWP+32tkddNQkve2krZ9K
imIAp9ZPpR9VvY1+Hj7gCfAl1c0vMbLgAanmLstuWMJOCfhkiKGHRnYej7jX2IXKJPiXyxQSVVYb
JvEUK4388ahBmr2ectLdXb8e00bQKvcp5CGL+FXMl3y9KJ2/Gswss3PATkRnQrz9oUrk2bgkzXlx
tlm3Fe2zADyMunPj8sBlqAezeNgm6GWecHyDhueOGeiLmomZWovX+YnBkJhAKmLXnbhv0Ykp8Jlx
U/TIyY55Dxc0x8EHAvA/tZfW399mOAFkL6eFtjGTk1fnIQsCmR/ZTju0DUnVilCx5vXsFYxsR+zy
OOwpnf0zGrWpokvXmjjWJ6vs3+zyTnTM6fVo+GVWasH8PkYLqaY+e62suPhINpyatkdpiSO7Uexn
YEWql8XGk1saFg6yWrfFmIFAXIQdYFMpLrQtI5RB2kTxgv8VM0NCNXzEy+4szeifZzECe3Ehkig/
XVhBfha947xHBG6UR6IdeagNvXTBhI3egm3BmqRGL9f9Ifxc9y+Bdue4KadIfc1lcWkb7Y1OgI4r
r1f/A5QK8hAakys/BV2kA2DujjdF4KjW+2YINYaZEpzlhddMTnTFmYJ2zOeEj8sTpTrZMhDzUFB9
i2n0K8J8Oxw6wYBB383N74j56D5nFzL+lIx3/FKbHkW05j05vNjABlUtOfywO5BufBeDhWFGe8f9
Vz5JLT3Illw5AADa2mSTCIdTiOSEsAJq3YCAviDH4picKjnV+MZn43C4Wu71LkPzkReTBvAee8kI
yk8F1vr7Uw8Y5NWAL/2CPqZT7AT2aakTndETAfOcucagnDmLpzhHmPRuUhlcSFqE/ScwgyBymz7F
55Svj3WNoNkSJ4vIQTURph94xqezg7JJlfaxDn/cVE7wgh7G1yMJnufVudIZVv9nWJH/0YBXfsbk
jiUXRoK8ut2+CsmtLx2jZ1UzuwmAdsXQcX2eE5LJkc3kNx/hPfP0qGzYSXexqMmTFHzUDfQa8hMK
napmPJ8RMYFzDL1DL+1JGYTc/PiBiOWCBab0+T8XQ8yMF2aWP35LX4Y7rFh6g5FtxtJ26fcQZFqz
6tBRuwDiYoh6tALT26P91j3ZXcK5+1ggfWiUTW2mqGM/8u4O4ZfXbGO+W2gBSnmPzac/rp723PWB
YOxA4ZJk7ph8SluhMg0zErLthnAYV8E0MXk40HjoKNM93JILNdRjnJRfjPattKA/VviBNAEv1RWc
UgoFHws+qwLpjZn0rG7YaaVtHP7bc/kBgEvtAljF1bw7h/DhWWuvpvJmCVSW3JN2wTMXOAwTyHvQ
BDSPmYBILnyK9oLZc1VT6F6iz86OgVPZzyO+G6ZYn2xaaRxJVMGrY2jnU256yr57xcy5aa68BuGC
NZ/PMGoQnl4icUAPkzDEsCJldW7umTkv3vXg4ESNjUXs909UP/IhJLnDHrlArTbUhwPU92A/myyq
3EyJPk4MNElcyLSseJPJZX34jXo4cJnEoB7XkOV4n917PLCk4oI35F3KiBWNLkqd2lb8Sc8o2BZl
MfbpIM2ahhlXi7Al/vnjmo74F5gmP/J7Q1tDlQcrz/4oizXmem8C79VB5sVRfk03BY+XYcEJ5KbX
Rc6mloO1szrLsAYtLcTh3Jq92FyL4f6KeF0eiQIVvKsrEX6nr0jN/ejFVtUFmV7HvRpXEH5C+N7k
Y3+j735KW2OyW5FFN/d7ZVJCvUYBh301zK0uo4ga8avEzFzK8OEzb+hljR28h6tiWryu4k9TzgLU
M7QuMNddlsv3c1FiEKsQJIfRgom7pb0yTdnzTu98Vqx0PRsTQe5H0ahstJuvMn/Il7qGVNENi2qZ
MhxIyCUQk3Q4m58IQlXjfmulL+w9olpW6QgJDDS9XbQD0aOw+d6cHzahTP65wt6BOumAVVW3cEYq
EBaia6HQYYMszCCGXY0d54qhpI6MCWqW80XKv30vtuOvcO8M8YRtKlsWRBkClJifjtz/FgpvFhfI
B4eFLqF1R5i7ldrCrh+UdeAHCIuIkCSKgUIiswxVG+SUxPOhv5NZ+e1yxRBZrVUFVXOw5LLqpudD
C5lh0EMbFrF8+M2LTi5nsnKzWy16xIsieOP7NxydeCIwcucYFBtRzxzcVbkGn+19rCrAOXTF1QwP
94AIRzdQ8krETTB4eb9N4nuoDbB753NRCsBZkH/frvByq8E1apz0Mmbd1zw7MK1tm3h3jfvVXAuX
Iws9/YLRd3IZRklXGLIURAZepdl0xveZW3DOVv6T3V+hVzPRYiHsZJeNqtH7uNQBYY6JZTVQ5S5/
7/+dm1l0YyHv87EnOyhoUoreKr7pv3bu60TMrV/H4wwJ1DNa6hV2NEaPjHjI6bn8y1zn938Qdt6D
x0MzdeOFyWFYzHtTsLb5vhFX0Xcy/VGx9wkhuto91mqYRPwIcaWNC9kUQzGyJm6zzAsJQMnb/nSD
wlvhbaW7cfb9xrBP+rt+QJu0Rcf9CtLP0X1E57fInAFPui4R4lOQiivBjNM2Vi2nZiQeFBOnzWVN
MKBc/+ajdfKAtElNeVOWlrTqRn7E7k5cF4rf5gh/w/4VdCDhnwlEhWqRNFWDJNwsmj5UUTuWKcDa
bqTpITWj+1X/pUCvbnZaodnpWUoWrYpDeFdfotQy3rCE3DjzD7lNYnXsyeQ5/CMHAWplajfPekzl
y1+NT280xwLtboPOqur7E6yiFzkjX+Zt9X17Sctf2wXBcqV88zeZHoWkkrsg59Bw1rezdY+v3XW4
oCy65mEVwQSp21JVV911MNlHix3F7E8IL9yMqFgs6fc9UawMd9JxAN4h/RSSm+4YibXazm0E8R4b
BMtclPoHfgSI7JbHaK0cvhXLlvIjePyi2N37e1MBa09sva41enZMkzfBWgs8e3xsHMm//Sm0NXsF
kqxy60quokK+BiSaP3aPaOYe+83kjDoKVoBbajC0S2xDU1h2juW+m2w3V/tGg6l+v94rbWqIRHz6
/HGS19LKtGe61WOEvFVs+zT8z37jsRQnoK627eK7I4rPUgNhdjOF82pbrYhQlu24OHTzE3UVhIxL
MhfOeKuSmYis5qsjL3sAAia4J7ppHso+hoOSLmEmswf6nc9dlH8KLjgz6kglQm6L5f/mDuEdsya7
3lIEGxuWNYiMIJhF1mWZihoYl5nnMj2rHrv0DyG2ZEnSfnTb2YPYHDGY4zfBBD7IWYT4xJIS8DOE
Xsj+1iHYqrMpmDgfGXw1u55xRYwUx3OdMZdbXfozxMhqyq6+vHJpiu15lchSNH45a0AERtt4jF4w
mTm/Y5uWFN1M2OEBFy7z16/6EN60+6irTNqYjkmRrx/McBPJVIO449xPmnaVJE6mPLT45MpjkMwH
jc9yFSWmDVa1nYHWXyZLKc+/sVUH0N6W1AEjNCbJpATrnNrD7ozHFUBjYqaDOKriIqwP+BLMkw3i
mKywn7ZP3gLTZ2RDHYehx8r6zwNoJ/AHb8XTfb+IZaG0gtV7bks9HGR9w0ZnjzqfDs4hWHf2/KxE
Qjg7UynZ8o8q4DWVX8aUG+oCYHtaNkV2LjUk0ugXVBWgFPVtR6WTXaDa7lW2pDecgy6rW05OsJmv
FckI+Jp4o8uU8/OpMN3OwaTuCrXcbHgKhKW0VmLrN25lYMq21bMd18tMz6wF9z6OAgLP8MXok5Pe
NEMRpYFrSvK4I/A3txrFqPgXfZ3LFW3P7nRt7WVGYzkQ/WkGYCgKykgvwf0lUSL7pG09w+INFeJ3
RMpxSsbr2jZ3lsHC1+oJu59CUtt+wJ2rQBkixaXIoQz96kCiV5auJrPW4PpDq4uBw6M2fKBBsule
yPSNSg5Rcgp7mO2KEjoJfdiHLkyhfjvrG5tXGHhFba7f6LcV3HaChaTzilFWe4SHTKbD8AdSgSjY
wURM9ypoa4in/zm3N0G5N0DYpFLuMS+hoZig+BhIUVe7iC71Mq+mmWbpv8354apwQnhXGZzP2f/4
XPai33tQOPPQ7GL8PFSlueoRO2/s450wlAq7qs2SVDw+hrbjg2vG+dx0ShA4XN98GkIoXus5p28H
SLmXUnbDEAySFUpnLPSWkCu14+bqcMnQrqAZfBnbXmevko3uGAWuHNMwKqjakavONeqFEKThVI7q
Q5YRze7qUEJm8eOmvKSzKHcVIM+/QEScoa8UmWUr2Y1qEwQGkHDdFpQn2hxaEvooKVY5/Mcge0o+
twE0XHctWm2lD2RQdamvhgn17RDWcKu9gM4zZJcxThePGGNrlMLHQtF/5JIPVt06ifKkssjOscvF
WXlkD5JvK/9Ko8flTqbeOL1T8UoEvEeI99rhzfzRleNKNZdxyLIry8IP2M4Nk/sQzxV1FIQasOBr
6YGHJuikPSGtx7TvPPctz7er3uInIqOKRznZs9AW6RSyKd4E34PkH+leicmj+lp1gJtCY8vSM3+I
/vLqvMuH5apwSk+tWKDXoWr7hg2m5net4HF7C/o/vp9ih5VmKb2GD3MLArW5+XzqCtMDh14wh9pb
gFzdT/3S6tzH+dNXK+qbzC7DEAtEIOhE6hPMVCfXV8J9xywxmn5b1onaEYHhI1i2YPbntHfG0UPi
rHVAtxqejmUJ1z44iGPn2qEc4y7FRYnHRadbf1d4iLF82yBuoJHxEpE0hd5rK10P1SF/jIKGsWJ6
nyVbcdGQg3huPSjkXa0sjIGys/iGrRbR/O90PoMe218vN6Oxa6sc+762yG1XTfWS0DW4MX5XOPas
+pei2ResB06tofp1HXCfH188tcNHCU57ssqJb9LOg4ftPcDclwPeEB55C6l18tiY+CGe20Ku6XAH
ZNqcn5WP3ibR9oNDxfw3s7X0CmW25FApcphvOMtEo3OV4TMsNCNsuI00TrTrPkOfJBvATu739Wsz
JClqA7mObm/91heQmCL8ZexDW10ECGHg/rv8ExYU9NTSzGiUx+o0U8LUlhA3qSjAsp7jwmn50QR7
pMgEP/9WFh9GnVRbwQ/Q+Aw+otOl2n1X/cy7PznrBKljwl7adX4B5KnAMMZ+T0DeqDfDAXB9DXk3
czU7Y7nQ8ypqT15L9X4aC5pwNF5IJsFPAhB7xbFsf2y1ncjLSVSV1MxPVDJ9T2fTAwLFXCJVHrwM
Q6DsShxfVtYbJ55D312nWMdgcb7euoC6WIXIIRexbGuJi1N6BsdMsZ+6pXS14jKx1GZhoAt8pzoL
Nq3spizYzEdwDvbzaGUztUyH0ji0PEa350fi0jtfVfZqcKM/ifdGDePZNORgPUhc3wt5TTTKQbuy
hDO1nITuBa8Kh58REit/DIwpQiX4I3Gyx/noP/VlTm9f7VgVUVwjB5tPbSCvhYdlJiDRBOp2WNY5
6IM4nnEYqPsdllrZ3wfW1MyNl2+l0pl5ScX5neT8T0dTsOoK9PWLHRVh3ARXkv1sBmot3qazOHhA
+0ztLNniNpjcqHc2ycsIb6K0I8Ejs1kECx7ZI02LzBiCcv+1akq4yWWfI+5fiELYj7rLNhWHIaIk
LAznLz0ldKC4YJd8FY71Q1edlxFk4Ain3TgWjPO3rHZytGQjXmsDhE0ZwVJt3mFN0Ag20ifFLNSZ
oNvya4TsKKbQRzo9JLwQxyCoHZNl7vVj0/eiefSAIPNtEz0NwMJAtnl6RlH1ILOCECZQouUxeOoa
sLloOLuE8fQBNzFYtLaYHSJR/oKcBuhHKpV2ttkse3ZTgLNGKodQm4ePcTpsRRiNuXmxL4geEBIg
EXTWMKMm7XVnBmqxenq+KZz1yUemhq8LkP0fNoEL37tOviTAGUY9FaPJpRTBc3ystk0ehygLF+eV
fuAbJqSUDPc+Jc2nehtfvoXjXpwoC/Qf7PcIEJQK43t6WrQv6cvG2iq3P5Ob+8N1c7xCVlWTCUlk
S5/n2DNcf6BRIbzAY4kD5QKBgnEXfKaCPDXfjUtPPGJGx5LTZLX0qsPnQj/k+LO9P4jbdgPeLZRt
AqOFplsawzeOpMQPG7eyY8zYzCHT+X7B7OuzouVuJn9AFSgaNncvv0kukzqYoIwbhGN0t36yEMYL
Kq1kG+0VZZ1YTpH8jxbnDg6qC2cC9Bv7/aGNsauu4zhlHGKUqWZcw/pVFT+4U0XQa10rykjZV7af
rWQvWz+3K/1hgyFWFqNFj8HpwFw9Chf7rMr8KtbtoKqOLiHhJnsVm70XGVuwYnht+s6SqSp4/8xQ
0K0AgAKCeRO6Y3eXP1M3isc9Gj35hPWIXWK8xZSkkbT2JroS94J2VfDLZT2wkt+9o/DIuVIIpWeV
aLRqkGUswFqnVHSvc+KHhAIrZ732AUM8SIrNs14+IGZ9OuU5mYYwPPDgDFF6rZ4MGKRImCSYVkOh
0ZdB0or2ZjIUVk2Hs+HKvUKSCG8/9fW0uUCO/lrBngduQ6hsaPgVFGyVKfmCL7WQUxlCdsN1kVgM
Tj5bWFSTNV4AIsZh2ei6BVehQLLZ4WkTuwLQmSpFLihYcDv3T7M6mMyadhKfDE0i0VXUAtseptHa
R3O+2L9JZjr701AxurGEqS8VXwXuLtlMClePbow4FVc+CK+5d3iw3eXKZxCNBKVvVbatWw0T66Qh
7UCJN18WQNMDTcAizKPpt4JcfN1MXkqAoY+TcSAOtHkPRNsIY3kvPMU7X5Lt9H6J4dVVd2M0F1/r
eE1HPc7V0RRrV6LwAKcnPKfHLaFIg9azt3ObpaS++x7EHJEWBcwlnaLYnHHzLKw6DQ8tencCGLTL
i4rl1Qm7a5orR/cn3SG3KcTkTv964NR2G9dvMBjO2aNjWNXGxwdOG+6+kfBYlY89j4kfYnjow0DK
czmYD6u/5wF8vGdgTGgiEgj3bKSnSbqeHHCaA/6xVUaLdxym1qFTa5VUrjj29Z1190uZPdL8NMpt
rotKJ5PAy+Q/q4/C1GV+OKQmO6hEw/gnhknpv20noYaD5bNVT9F8LIafpOqG5hFacSQvfqlOX+6Y
lrFIJOiLlYAmeo0vTNT9B02nS8sptfpqBd41eeWkv3kZBfjauDAm4ZT0NO/baO69p9lxSyPPUD9M
W2ILmOzWwdLI+IClr/02jGmkMGAmnyvowtC1PUhEVg7+bdVvD29fiiZtlii5TgG91a2gSCzYwl6A
EBDRQTVY7shKB0qC4Zk54nTp4z/GgWeCHWOySjrrrZSUzfPKNMwnjlY9c9CPULwSMCOKZCJXnNHn
xzd1GCu+m5IT6so2kbPJbbUVnfKU2lAsqumpAIhnrLMrNw/IdVIP+Kb02FnBxMxEYux7f8bxxipy
H1lNkGcDYkz4lvVh6YWVYp6G0pXSteoDkg3CE1D/NdMhXxrGU2od8TqA0oo6ROBZOSI+L3Jo4OVr
sZKFFkObWKJtsKoAW+V5zZJDzgMSIUl06OIwaI8I8m0erUBu0xtCNRuMpcqcc0IGNdYCBVJNlDS+
HnAZnQVHG7uHojyGtPJwjohUBuchqFQoVZJMU+rLV2owO8DxwdIkkqgQVpAQ9TeVqTecEJW5Tzpt
+6uRS2ywxdjldwRx0eJjbIoXvtfoQllGmMT+5N6Xvl6n5zk8oxJDvEfiKY0Bcgl/zQ2AM8cfgTLr
2rCvzGSeP67hneXrGhSRS9N62Ui88rk0MRzGB1c/sP9SZLrNwse9OEoagQbe0OGIwqPAZNm/QyEq
GwkuLNT2DO2Ghzt/o17YMKo06ZPtgjg7AYZWSkj2aufG3BOrLRBUKYEK4nTicG7uP1bqZc7riE6K
cSj1iPPh9584LLTwtkVoQcrmf5bEH9BlsoxHEyxM2tvmqiPsnkYswpguf+6VmoCvUC9xxcOU/ciy
V2baCczOwWdL2ADeWd4mSZOPtcP5Zex2uvf2nop5+8D7Dwwk4MHBQkYxPqQgQkCnpAkaD6bzghBb
FFecfN/a0YIRAIeT/xTkjEfUbBTFc2DvyK26hPwKCtFTIK+4AzjWL2PACRf8wcodgWIvEV+1RO7Y
GQDcboNNT1rSMnxLypb8EeVxHDOgdvz4F9WbIghUwogRIGZcjwzc3zWCXxjACji8X5Y++o2YFE45
vY93OD/7r+uXhqZwffzd2ROR2jv7i7ayQQP+LJV9kA1vQwM9iz2dEsJLPJif9Qeg3Sy7PHN8g1wz
miethgEJps201WvBbMo18uEaHYeypBYRWp55JJHBfm+Utqf4x1wiSvE6ARSkgoJBHVy9WHWfSMRI
FCoqNHFNzvVWVLj3ndadCrWMOhpvAdZSZV6I9ZY7lDX+XFys591pyP6NQmjqm8AWIUBE4TywlOYw
LgK14k+w4ABUKI0Y9Ez+PbzhByZrS3PA5wkZyilW+Vb0TO/P0tHvNR5SJ7Orf4fbhmDcOr4OsxNm
4ZUzVP3cbk0hBTg+pnPYaSmJm0rVbsODzHmApzpHkCxFJjXOKWc7bSezu9JNL+hEERf7QY9Nmi+P
pRQXYL7k98RkFP6soPmRffVbjLdm89WUysqkaGxZFbXXqf7Y2YHHbPzQR4lZXkVYKTKzUSPWwqUm
34Et9spv+ajTMGuoNFSzJMgSehN9sQxpkL+Cp1fRn6QvYxL2kpuqOiPp5I6wJ56ONMUWdds/9n7Z
QcD55xjnuHpb/Ix7r+SUGs+QmdoONKe18KcpHsADoVzBtpAQUIBw9RcCZwmWsbSoNG8bh2P1UcFS
ToJGKzc1SU2dXY6Js+cc3BifSDh2OYvi2QdQS25oqMykpCC7zOYUg/zTQfvg7m5yly8loQRhb5hR
9AOjEdQHPBWkUll8fmbwMRsMxzcGJXjO1UVaHu3XGGTQsjXOGlhbfPAzxTngo6RNRBpafuev/4cr
YUfHUlXM+pWQD3XqRGdTSdxJ9VVuxLqakzWpQLzd8fERw4kUTKCd6DpP/FsjbjLC+14l8iOdOhIM
lIt8llEohex+obYjUSVZK8KufMrrPlIlFx1O9du9DAJvmZNA1ucLOPYs8n8dGvWdbUlNe7XAPP4R
ZzL45AiOBFdYulqjeLp+3kLp98vjHJMeU4a4uaYJD6oYlKLELdchyR0GXuvTFxaRmZKTPxyPaWCa
HqU83303B7gPEcqVDoXCynZxo5n6OFyWJsopip3zGB9pysXu9judfthHiKtfXDwDLGECQq9W+U/r
TycgOxgudIigFRZCIyx11OnSsWMcVNeK6tgd7Nx4h8lVOCpmLKHd/vZcy8r45EXWU1jp1XcM7Ljw
30+zSlNfKX10y7ky7HGPyCg0ifIffZIT3m6XevR+RLJWwJtGjgzgdEvx6LuG+58xXnbv6XNr2IAi
tXqYukLL+gsPDIUGGeThbSuh87JoMfrDepWYGbJYRNyHxBQJd5LvxASYoI84csf0x/FHqU0zRnhI
uJv6BtcWcKVB5JuVufVJiNXF3A+St4QSwd0Cnq0LlHd8+XGaIcq4YUDW66gka2nW8oHj6Avk2wPA
FwC4FcoZIVSqVBl5cMro70KA0GGU18UxILNEl2VwsFk9Pb7+h0akySC6+guMW3lKe9OEacF+GV98
bOQtv/D96He3WHNEn1JZHYyMgD+Qt+Q7zug7N3dT9r+bNC1bjEzR/IbikZwf0qjRGcruDf0F0bBM
o+4uG7QBa7HVdtdKdAEHtb4HuzZSIxxnJrvojjN89yvWInX7N99r14jALZRlR2qLeWU1R2Jnvyec
Eir/83/LsFvZ38eZffhJE2kt1zc6Jgk7GkJzIEKBJpea8RrXBhtAiCRhgEOQBtR2cmafDm4J36I3
eeefCSIlvtqyEJAwa5WfqYxIpGC61LOTKjrpBV2PadZyDSq0I9o4NXnQkET9luq87Pqzcl3yaB3Y
hCGF7ajx8cOCFObcogxV3qXrtEFsEhaIKnbF4FwcOfstGBTpCx7TLLfHXxbAExOVTBl+yVJ/ibsS
e6ldEd8P/J2qWfnO4DX6LTYdn+WE50pBbpYcFY+enx8FVTe/tvyaCNIuI8CGUDffVZI9mWxemwG3
CHJpiz6cHHPmUjKtCK36gqY1ydneGb+swt0TIBrxoVzAcUHamJZKqdflWtmd2mpGfVfKahTBOHkx
TOc2zwPeJpSCj8jfnXeRTMIZU5XMrtY+7MA5ulcVJV9vyD3jEDmfd/C37JN3BP7kb5DI0vAhgvbR
aT1g6R6NfB21+NSEYBKIV5PFAzf2dIJMOa7Y5fI54c0EEDKujuZxRJHi2CyvYIeEl5PFreDABYf0
W2GPQcejux6riqHhN/8HpPgcH8JWp4EgiQgTHXQsN2+yhT7BGZJ5PbjO4xDPnBfLZGOtTJSCv2gV
suDy/DNAHwojgzbiGtk8x7crs6g9bal4jc+GNRxP9LnCF/qfl0RzsQ9DCEM3Z6Sg8Ki38UsRBSGs
Xawl5LKnMr2T89kfhyVr0Lbj59cil+XeUDPls9yzqlkqW3/j87wGtYWDNHt7NTsVHRvO0zBGVEOc
XYzmqOIPti5tH3g/YK5VOV1QUTQXWSRNRmAY/iW/PLz2prggJKpEt3MlmWOwIZKjzU6lACoZFoL4
Sy0UgbmvXf4ujD/TkPEA2a190+mDe2wtlyqfAwpsFtLZjjycNM0Uj4l7AbyeSEx3FZUFhlz5CFr4
dxThKLBaRDmLYgdDkHY3zGLzPsFdg1S97tXiJSE1W8CnPakDBoUHVAL/GuvKgGlsvvtUo4oMK0wC
vMH8ISSzUFGGzqMuDmMUTrbDNMGsqt7r8CoVRpxLaVTS93ldF2KW7CTVxkyOb1mr5i23WpH9t00v
QZNqoSgBinaQbL4TvglCqMR1gjVWI0lujEYQlDPT4l9lHdeRCr4wi/nFyV+LZzTkZoaSJQ81PP8g
mfcre71W2Ts0/hHzEVl4vWbzSlRErJdSk/XVXr3HouU5v/8WlR5SJAjiB405c6uHv02hxwQettjK
DWiVUNO5P2WNWbfR/BDTJlc2qB/tGMhOC3x1WSxdGzo0cgv7FDu/KrVkwqcwpdNpKmtMxoIhMOw+
7vLYDdewVdqNRGh8LW0nXVrIkrQTlWpk1LAMSh9K2cWIRKzZ7oo9ZP7UcGeIBvxwuPCUWK1CZfty
B5xQO6akMuJJIcNpu2ksNsFdfI0lRWaFgwSVOvbG5oLcpHU+sNnYn5G1d5dJuYuXk8VSMDG0Rz/T
5EKVakZs1E4v/huvGtycs+KGqyWEuKqj7Dcmn8XmHZ/9BJCIv1cUeE/ENFDRLC9n6NWymUPLrLjN
JGVYCtD80m1BHROAF5QYso1T6/Vef3URNMHZCHday1VUdy3DtbAJuGCdjtOQSDexgqAMtQeyM7Oz
eNok5wraieo0ssGDl8PWDAOSvJoa6iZWs89lasWfh+y5uGZR6ISi7HC6FonCXWP/KtZyyU4Z6tNl
czpi2v8jsNE0SzXdroW0VG90xQvGo760j5nbLJ1sqBwCrepfo8c5e4oHQML1ODhLf/koOe7jFn03
cMpqaA+owyFkCUigHkHKU9Fl2ZU9EM0EdK2hxmjbg+3lFm7LprGnDhBnBWfDhmpgKlyTq1qMQ7HM
VqVk1CKrg9WC+46aYFaYXKg5vkTImD9VRQN48i4yxYzFDm90IYTqRFJSYv/qAuQfd83RHH227ets
jN+r0IM2/2jiOttKXDGVM1GUex64seNXLjbvpxHAnqHezmIhNzi5XuezXletnCUQwJ7HDQE77/0B
QFJW9duKuDqhzqOG+GzxiHoaiD+UbTurr+pjQUbErzwAHDiMohwU/ju/EQDpV2mtR/h5U5kvVV0i
mKBLXJnAX1l76PxxyGiSNXcZtqbUKWFw/OBP1ZblfPPM0G5Pr5Lw3PiY56mW2OMSAX7XTR9i2dS8
ylahlxnV5v6vcOrMnNujjNaYoIxSpjvRdoetuUfWKnxVnU1bDYQIfbLuNDVU4Ad1QCQXAtz3r6pW
CRMuKZzFckXx4ZP2duTjgFvZfWG6xifAXzJzKZVPVB+Z7c8OTAcjVuUA4KbxpJmmjuujlXkZHj8i
O1RoYdktLj/TUOIXDgel4/3ThvfRwXCo+iMm9eh1nkd0+PR+nU7JT/a3SkbKs8B8pL/EbiRRq70i
bXSIfhktdNKr17/aDt51RZzrcCtyZzumJs2JJJGDELexDhAFVNp7L5pBaKyQSXe6GU4oz/Dwj+iT
UjgRJwTiKjAFUzdBJPeaE9CJ700CyycNgqs2uYh54C461rq3xcxkXjd29dzeyovklHgG3pTKalvW
v1WT7FbvZvpi5+50rKb7F4GYLCFgRXvEXcRdqRyKveTMBsrtxhPaXC5ZH3bTq6u2bWj7CVTtFtF0
P2YuITUsOaiGaOJj7LLdaRjDi2hoYSiYMPIJyPUGsQgWbnqw4pGVGMcTY1818R8KereF5XFXnvbn
twbx/f1usdWyGqrALnZU+fxBDikAY/pwVqY5C1cyg3hoNLfrZAD41SmttsTwq+kmPA1MTE6eqAqo
7H3XDyxAi7dFkAwc/F6YLHJhlo+WuqkReZ+TZuYnGroqzo+Dj04iabbOtUFlV8SCheHLD9bKrjiC
spwZoo2EBorcO5YJTlXOVIemDt42JPibaz1o3RVc5iLiXRDJwis7W5bGBCrKrZMn4QacP0Uw6TNW
tMG2GI3+zaRNIoW5DNrSbmh1a1kSo6ogTlGbeOJY/3v4H0iP2IwN+4JSN3MH5bNLzoA4K7//MCKm
Gp7vT9jJqtADlVu+Ajvz4KA9BH9WqnUoX4KE+V/MM24PFymirN1UXmGU6N43DCNm2a3Jlss5ke0P
W7M4egDc6uAJfWQORZSDw3srmxBFFeUvHeFcvN0904A1k4h7v6qOh2OWGmhX/niG4bi1wcmHHcyz
dlRzr2LB+hPy/s7GPeDcO8aXF3lnX1ASAAukGr1Th5TeWTmZY+c//9jyFpwRMfG13MKwgqLX7C4j
+MUcYkzRFP3vLrJI+zpdZfqKg7Ssfhb7uKqypVl9af5XFRMRf4iIFqqSvpEL6qmKO7NWHZXzBNtb
5/RKSWPgMrwMCrABewTt/FQxH0B98b9h80l1slGe0vyLnLyqo/9mrRPZlW0BGmDfmygE9JW9rBMK
fcUfHlq1lVHM6PB+6ImBzPbBB1FRn7DVHMhXBT+ni2TevgVBAWJLqP6zSQ0jURJSrwvwN7YMQhTO
n/XIHvtMsLpS9yAeO3SnRJqOWRW+WsL2a5ReuwCMCna5xSzFER/keH9gjAvpS0ub57VPhyUajH/g
b+VRmDCvaYxF6UjCCovLdRNkbXTg/qRFefla7ji1G6/bFssWm85TuzDhpgngp4BOgEkWBjoKvHua
0a3FGmJzOW7HBc0jZd1RSzgdx9IBkom3L5Dw8vcSDAcItD1lTzLOkco6bIkUNODVBLS951WXf2OU
lQq3QOt2IuWX59VB5D7jdcxUZND9HmZNj96dL1LA6hpau5pmFiAfW21KMYMYlHxIHnuiFYYq9LZ2
Xhs1OWKWEOfiVJWoAVnZI9igB2VtcP2hGgqI2WeXXwoFvZ5gnpbcVLdgENN4xnXYppMNmRiXyh/C
4Z+jQw7eErTec8j6pypImPeMHPdn85diO12UfEEdj+w203RvWAEx5La4EQsKJBeE/YmahTbvU8/R
cr/0S2f+Pr3dLuymU1v+cueMJ/TgD9jloP6pzMuGRETn1Em7lji/Xcy/OsyVeZfiilWlPqzShlAm
4b0TGbeoMZ1zx38NbjIV2YABoU3F53GnancL/20x6RFxz8zmCrVdooV2u9u3dWA+p5YlW1M8R/CH
/7e1BPlCLv0sl9rhZghvJyxf8Cf1DpiTTPQ4E4OHERnAjXb1NzfTTRJRhlSYLCCCEtE476gYXNSZ
THCXN7QwspqtPI6o+UWHgU2fevT/DsPcoZughB9FULEtVQE6gPUFVmurP8GCubQfg1UxsJNsHPJQ
Tg/eZF3xMggPU9q5mr4XAZVBIhISB78DCbcfY4cLecOaosd3Zjg/vBcmgzK4dt9p0I9eufp1G/vn
Go+JnkrdsntURrmLrPVzEjJrZg85mfPqVsEdxEbVcICD/LvWb2C+OCSIUgQhRKpRwip2Pb0voGX8
uoeLwaFguXnhUC+iRRzw5yBdzDk+YnM4Sv5jbAP+EyguUQ7p0+OMnw2rRloG2ckH9+f3cTa4CV0M
2fOYxc7FURv0C4jfjX7d1XvavucVro3m77o3xlSqk1y0d0q3emr6UywRwKUzo5sx2sUK7Iv3Yadr
SD4/vB+JIucGeE9SzIz4IJ2t18Vauu8wsr2DCRnNXmTgJX1A8ntjGT0F6xNk9q0tJbgXDE/bMEmP
Ztnq9tv4VE2fFHW1cK2JChzxb7Ua/WFV9gN4rSSzEkVHGaV/1MwMbm+T5ObReA2Yc5kzkoYMK3s0
puUwJSHNnkS9mYa99YFSSZl+mrE1mQunnSD6ZMyNxcCPtZ339OSG4DncVr61OgR8jJWMFqoKSlsR
DhT53/zYjU766uU8CM963CqjNqGti4hczBy51hbZbQTkEx6E1KnBPxFMj9rZ4oilU30BrTQ6eopw
bzVYgFkA5DBn5tWiEcGdmCNAx0QelUNGTp3c7YQOBqe5PKRt1rf4bcGNVEd+gQkbWLI9OY2JxLP2
vRzVbKMPvdyluUUxZlZ4lEhWlPWSVs3FteH/rZJEqYOCbBZTufYBN1Kqw7a3OYVqEOl7Gf5APN1S
ObR6QibO7n/KSfGCBmC9hUu7/i3LI8qe7ow9EVir5ZVQ4Zq3NcZ3SFZj1eSaZxhQ7fcZA8JFxwZa
sccUzZJHWKzfX2cB2dtbVz3Ga9TtOLMW5ZtLihz5emyKwMHPoPK428ZSUjFl08LOvSJVpV/OasHz
wh7RywoiAOcW4lBWJDs6RJKkMuRoACdVb+YD32IgVNJ3PlWXAvdWYl2XTWxjVY5Yvy0KALF4v4+z
YLiYcxAPZJaUXesK0v+5Bl2LiVsiJCVvuFtfGEJhvMfEFDgi6TCw+t6Sf2iDAJo30hh4b2cBTc4Z
4MZJCIsQctH7zOqMeUTKY1ceOAzXWWoBLWaYV/dlR8xPguamn+G+3uTXMX7lKvzBVHGlTwteqIJP
vMrWY3+wyobI7E2jXJ0Qn1ECvJhg8seO1Gh5EKWCS4YVyLleTYQ9oT5DHgBhULwzAd7ZZAxIwufj
Ahd78o50YmS7mODg9WzF8hEOdSRFHSueBK3QDZQTJiLYuu0YVE4doj90T4MXpiGONSfVRtH20u5v
OzaUpbSUvwyqzEAkm78oeqhS0XiYcgQ8IaQqzrP7Z6Rdh8MKTNvRbVJ99fvnju/ehSih6LpChV85
Va3T11cDG/uLPw4U/8Pk6xb9ODcNAYER111LBbi5gfWHTUXhh6VVOR0myyP1F6TPIMx4Wk/pDPMX
Ln6URZ+Lldz12h5VOtJfnwDo4Nlb4DrSXmjoHoVUESvqKzV0/213zoUaypqHIERdvSL+IcqZ6O2s
e4UVwFw47qfTmgAqs5Y9+uw3c1SqXkeoxNA/bswleLaviYYQ/gSRFMsRHpWOg1ew0Ze0cVfgec7b
0qWdVSAZvCOv57j+7eENmkA5IwZMdEp2RKBcCyweAmjJ+RDZ7K3WM53rmWf7Q894QGupzgfh1O0F
vDPKJZQWcyHbRbnq0OQolxtxcmNwyqN6SkKUO+0/0Lk8y9lNCdjYSSW9H6HupBDoBXYjzJq4rb1k
CqNe+fLDpWRdmfFOe4jW7NCLBMWnM2HBY8EX+5JB9lsofNlOPLv6fHHrpooFiCj8S7nHKA/12UOh
e//IVwrzaUeUxE682cUqTgEzQd3YvplmB6sg7A6jmbogmhBPW6M1iHU/GL0XbHsSB9YUs3OkNy8I
dLrkiKHz4lwo0iKwXC6z4Rbx69Y7LThqNXuo18d/CXxgKLXkcu5nTJ85hcMZL+knpSVj0lgql3yP
/5PuiyvAjIGaqemksdDhzPk1Vr3/tb3IljVkgZ4G/ATuS9jXXY5+UdwIymVy5Im4HehFvMKceTPL
7P21JektmRitGzBiXW/j/KxUjZp5VqiUQzYVE6IttYCI3GSaYJZnUtv9URVl/29510dePtkEZX4j
XbUIRtM0oQWUp9Eefe4Cw5qCNK9FXUxS5i8GgDHHUGby4tX7otxNcZV/q7XUouI9HBqHidT7ixBf
2UZYlNLEyCmEvWBOgc0oS6iYT0TauAAUVq4Ac0MaGpq9x8O74r76OV/SMgIdV634QPoPu8QS6i20
Zgww6oip5SvSKUhIxSaeqEY9RDOpQSZt3aSgZX96L8Q7199YQocLfWV5LYd6y9IaqORdL5fy7d7g
VuEwbPVcJpq9fAiEkaPB1VdY47LqPHVwaDySyotT3CQM8Z7r1Uk3qvn7cBjaqzVt53tblwyBiv+W
JU1jb2PX6t0oXK5J+n2lOzP8PKmuj/JAZ2IV2H7fJkrqHerz29NHRTAYJ7v2lSuvRz0R5bJ2aUWI
39Ls48NyyHkuy8qDwIG/+3GEncJHrK+zq7/EK9niTurCvyQQ+bhb3kjd7X8GRGfbDMCKIzUkVr59
BwsaBOIfUB7B6JVFWoBxfqPKznqeqwcqa/krAEV6B5S+VgNGqd8OJnZGJ3G/Ehv5V21oYkbR9GBr
g6GDvsqv64MWllBDJDzpX5Vs36Yy6zl9naV2LLTJs0cWwR+RljRLiOCuzgHY2ahfaXDqNT1ybf9V
o2aS3EKHLjadozKGP2MndxiRaPx2UeRrcGCStDj6YR4hBCGKmAaJtSTUrtzkdMyIWOHs+nQREQF5
16SbsCuxInnxJ0k5XXp3rz8aYrUnCecJkDtuKuE0RXt9iDhniErzqUTWuLE3uTKNt675hIy/Ib3N
D/uEcnLWgAfMSsM9COk7nt2I1lHbamp6+nw2w1tToWChzR9P1u8hVGld+Afe+c23xn9W7LsZXo04
MTi4/VwFEo1XEFyyL9pj2QI5OWfjECt4bMP2YgbyYmQQL/pJubfW7GmFd3xAgDJKOGWeYz8GWuQx
GUH4ZE1ARYF7eVh325y53QVggke/gzjzCTReWbyFXhLmRP3Qw+QaS+tFxgMD5PfFEgO1q5KYAFjU
VOReYihs99VbxYRC0ohsvFs8qp3EH0cHz5YsBGNP818aSfr3bjVSAqaPE8a6aZDPa7hlCb9ciGol
ZWBCII4eCxIaZ1fxm6Nlj0dAZE8caOMMd46R03POu+hL/bzulbeplBUCYBtMq6Mt4L3QjpTVD/Tc
PJgSunLA8dS+oWnoCLVdKzBoeAaXYKKLe+he85noUOuuJQK2w2Aen4n9YxeHczNBA1lsBYH7goTv
7d8kwNOXi/E1pEgpAe6brbK4S69KqiP8aA/VymLk6ILs4gS+9SBNIk2PsGrT9i1zcX27H3CmfiHA
oNCw0hdL8ZN+nmTcF4liFoO3l9fDNMbRfcHmcE0FeWf9jHFzGyG0kDDJG/FtIqxHoR9YElxnh45P
pRGw2vP9ttyTCcUevDY9ZQv+RbahVRhTDg7PG54bRxpCBNpoJjkqSapiqNVjKQMx+3G78e9LisvO
tA0JJBKuVIHa71ja0kagHHmA0TiT/qdZ2otMdUDb8QgEtyvp39Z2nSvvMUuflo6UqJE2e8pRfyZh
BfHspfaEU/WLE9UDTPLcBY0S/8ktQuDuYY8XVV+4+xT+XnKrDNme5huREB4ZWZePXuB4Bbvz4wNQ
0PePbkET8AW2bd21yFxTDFzcJ/05H+fqm7Q6PUjQYu/qmJ/AfzaYC7bOFXfSY5WlPiuMy8SRn/D0
9TWD92t30CfplgvkPljH46Po2vS0jl+LAhINIoeXeO19uoWcWPDCDQWKe+bXxWg53XrT0tKyocHp
K0GoNbfQyxDr7Rl+Cj5f0riHUmY1CTpjZ5tYRUug+ao6m27S9xk4I9Wft2cR69L+AEUUJo2NepXb
F3/cxGOQH7Pa/+tJxaN6Fh9ED9354c5zOwJznvOuwL/QrC7FIsOHFIXG9/VnJ/dc/+fGlUXKLiC9
O9Bk/vlYwybkXM9cavtoEDbJTE5x+cKem6HBzeais6RyGEKTxilUEVZoFF4ZkdcLv+Q0ikYvuCPU
oKHGnupzR/Ma8kpshm4+lIsGQd2wpcm4tOWAjElxAnBgrpVmoXBgMvab2FhQZxxPirvpa93c3G7Q
E3O9kNS0QVaboDF8p3ET9wOj6qU90iypmEVyqNvzkIQ5saaKMlI15JLPpXX++TlUlHheYg7bl2DS
KoB3SI7I9OdBtVkOtRTT1wT4SDQo54B49xdRcR54i9hYg9DxA+RCJDI2/EHB3qQSLpKRDP5U1vpe
SWly84qIX47GYyQgwo9qYkKb4J+OcJiGDeHAMCLEb/a+UqkzVEZHEtfCdBQei+pQMuR+cEb4LdK6
QmdjkcnGzL3UT5zMVyWpAoQhG9yiqXvIzxiFSFw6yxDca+ZneUz+Ms+VyOnnIENyiKpU2CGS18cg
fA1bPODJ/iYltAihvChhvjW+dDHgwGFGSTMiGEwoROTCFGeUGcJcBplL+bHvxWAxrGVvWfIv27Ip
lDu0Gw9PzpFaZLK9XCLg35jjZD4WnLRls7lHQ72rr14shrGrbCZG4z6ltuMgwl5uV0hfb9ecFZZi
2yypDrMRVzaoNs/HChdoT/UWXymiERwMgK05BHJjdb+s8/CZJ8mslqS8IRCBKVweSDqQQhN+cFJ5
6vZpeUUKgHy/tuBLAoS4UTEpAhR+w3Helh5Q4RH8q/HgniZ6/3HauJZTb1BoNUyDonYAKefj1kyW
jY5kSsuG6DE4WAZPxr84xs5PDghJ71I2wPw6Y0mQ+eHpDUIxfCoCCoHXI0ZaRWLBlnR8JTtr46+s
YLsC7VLPOlIIvexlWUQ2cl7yd7+lu+UbSaKl1Z+T928TSfyGtrlyEFeG33yG2h1YEVUsvRuKzkC4
WrXIcoVoJ8YRKRJC3p2OdnUzYv8oBUcv0KqQpZQQ3QILbYz2pC3pbgVvKKk+wJxi7YwvI3CAu7EG
swRJkguZ4eD0DJu9sXH5EY0fCNGCoMqjc7PLRHKxplypuBZl81O3xUDbdn4FrXepJISiJRntHff3
7nibACZ+yrtkq54vhpyeHwX+egCVhffwIPI/DYE02npfgoIEFBajaDetYYNH8FHs0MGTfaEVtn/u
AVi9KllAbjYEBfIKfH0W1NROPq9RmhMx59HEcK7nqJwNgpUOnEhkAE7xiSByBm/JArkJ5PA6F3Yv
r6zRXcSmQl7OZjPvK7z3djTeaZ8RvERG/VN8KzSmBJdwszfdg4iINl/z/yLCYKKH/YUXirBz4pNF
dp2nFDA1HFWiz+kpqyRa7g52/DdZh/kX5PIcRQCbsGAQ7QoLVYMD0unrEpj/ZcWtu7Uya5utnzTG
tghaor65a0UPcQJg5vwUP9pg6zcv+G5lBV6QMk4b1FjBDm9up7PjORDNxNfBT8dVMO5taQyvDm24
hntYwG3S0FhAIcTEteq5bREuLEbX/z8oDjeZaMt7keSMpgkJOHhCWS9Dih0P8rrlyqYWxdZ6jz1j
MKrtbkRBxuattlG/ZdB/tMN4MgXkVO1HWwLei5wo4eYCqTKSzU9Al4d+5QLCzwN5M3tCEGmrZA2p
Cu0pGodEgRMIBJn6LFGtoBXDlWlbZJcWahOIOxK7MlhfQ9jdczYUvlVmeCdfoJYRXppJvs1/tOTm
ODSCx77TBIPCgYWaNauQ90GvwDaa2VudNwvEZo37UzGjmDpco9GdY9ypgGovUeC+AK4bAODI8ZxC
MdAJV/Nsikn9pDB6oWVoX6tTX8DCuuFeC9eKAhYHrHT4FlZiy1ebZSPjJTVWWHvOd40n6vo3hcpG
0CKUgWBj+dG2iXA6RBW+21Y6DBzsaG3PuKGi+C5coYFqEm9zoSTMjaGBZnKo1fglIT877OPRbjPQ
X3qHy8HwawA1PfOWUsKRj/JrV/cYeftjz4EWlspLHJmUaxMbKYapXjMl0iTBiqhLp9POnNhID85G
873dbFaCa7ZIn36jkDDlLnZbXEpG3KebgQp3qo0T/r7IPMUp/DzRwcOlPk8MDiX6Q5KbMcTD80H/
rkGw8NbVx0zS/lOSnCcfYfCW3fbiSasYU1OaX477C2nZFS75KB920lGfV/KW1V8Nc6pVz71d72Xb
XEODOb52XZW1SZ0sdp7FVBIxgqWwt8OfL9ot+DUCprOP6yPATyYiHNZXIVmO4CWe99fon89e78tJ
CRFVkwi9XNH1agxrjw6tmdhFfXO+n47XOsRk3F2Ji/MutEbIy1CsbXMLLMQ3ZQ7luaZNCbDlyXUZ
S+0fua6wcdI/4F0RLZcoFJR51xLSC0d7Gr4wWresh+Fon3XowKLMzUcgI7P7G0LBhBZsmhjJumRG
CFdt/JEO2cIkGBXSCmaoNP8NPTaR9CObk+68ilwECItbPrd5rcJYVXfbBkbggbG9BMSdrLUqseTn
FXhfycKYdg+VtI2SPqol8l0wkWymbAx0I3dwN/2ggRqN+WKVycmsQ7K2srLg40xG3k+oWWBenngn
rfNxqaLG8UcfoET81Ipvgh7EdLCF3fwXgwHjyz4BEtmoKUIMh4Dwm3o0y3UHMLkvMY899MqDwnbp
I3jR8B/HDweTE+T5XTQ7mwPBvVi6boir2YMJ4WBO22Yae0r3HyPr46pU+AfrMcoSUqI/t4SxONrc
wbs7fiS7wV82Me2pfQFqKy6f/oEViyuCzwQF5oBWVM9p5tnm0OzYp0ZaXQPgmMoIjlgYPx71CMMK
TOz4jsVLjNEqPT0qKPvsLCM/COtjX2weYTZP7O7vcdK+gys11uNqF9rOiO6uNC1wh0GxAzwSGK1M
ytBy+6bDPT2NZyxMzvKxboKPFHIUIKkIgpWuDk40h12qTkhy4tUU3BKK9edxtPckfYEtywg721oL
WRMkvj2k9Vr/6jc3HDyAyHe5XaBaWu2trIcsCxpYemQaKQtHoXXHG6HLo9HWdAfMoh9AHjAipshr
kRvp6RlafNzthJzBdHkibYbJ9k7CBTOaV1DYxPkhwWbDFZvHm+h4wgTov+Fk2vfNaylTPbgS1kRE
JWycAGF/tclXMkI6vsdFCvBghpU650sQ4D8HF1zFUEu90E/hjhRKI8LlbvfMu0RRuYaynhUUlx33
c/VLNNyrrIIlQx8yJPzN3dhhjfmR3axLJvxMkKEuF6JTNgOhh6hUFf1iB8jqD+d4XZfxuFObMTTF
hcVrFgHaiaWqnOS8VqMHNM/t9Pljkj6+ULhJXjXRoETXAzf8i1s+KPIwJ6ChBqNUfPLYQIjS9kVD
6XzksVp0RmwNAWe8rhaoEpSpWlCtlQugjNU/tQi3+vjEhBYwLySCoNZvZQlbI+PiFir98oMO5a0H
C/tBIfnWITrHuiJSaGBqCEjlqb/4QsJnobCTNGXGc93M/ryET5GvUCn55AKrKTwATEjvTyL4jl4d
zCU0TDIa6ed3vx00b6W0jIPEBBMpzMe8mUomPTOHuaP0RFUr9bLl5myfDJ445BfQG07pblBvKwGL
HxEREtAG0CuDMy0G5qBQZCqMI+XDrXNtoaO57jmjVoMWQsqhdWHYzlHpvUeUvDVWv1x1wYBtbxHv
ij/hLDgRGdak0JbrrSFLqrNR8HH0iYF0cIJRmCwBKOloHnQVE707tBDWJuVuo/OTeYqem+YeM0fu
e7/qAbWGYi7PyhzJTFg16R0Ro62KyjqjPIHqUlo5PyuURxsuF+qBgCpYsxw/YDYIGagJwOY1Kcx0
yhX5KqTsDvS7UOszJJn5ztvtTegTpEPD/0VyK1TULKiGVsYFfjmodfPFMROK6bnYELugp5FROvxs
H/MccGwiBzSM9Yq6t6iEe0c9OU5PB5axwoODiUcIPhw70lxf82gm2UKGL1UGaER77Ige88feNx+y
M4nm/yw9ihiN+QiUpVVdi9lNQbZ3evwEcmuT5CM0eq4Fzzmrksl1vowT5dfvMvsBYkj4SZDVJ7C5
TzZi4YEzpAsa/ySj3KLgKhPOaV7TThkaC0iVEmjGrQgCNcT3i0vhZHW7wA8shu1qlyntAElWRlSC
rklDRrZoGGULkfVrfGgk8wrljoxVP8wmdW5ggSCh4ZGHkp8O5477GWkiK4kHG2U9VBBcaxuqCKCS
tTMysfKQCFx4lDuHbyt0oyMnWoDVfKuCBDFub7AOplqKg+UlhcRT5L+DVdbx9G+2BSe0fmk+Z79j
eZKzNxsKyVZEfB4wa5lhuM6EW0Dex/9lVjHzFWmXy2BHiBFWT57VKsHA68wPmx6Mm3gJKoPoyfP7
Vf1hwO1m3rOWxCNu32AcQVoqj4t3ror6rEwegk9bKNKcYT+bxHciQ/wmSK7CGfNYnkyopQJx+hMP
LyRp2yEDHHR7seVePETIafHJvYv94Mo+XEPxNo9QvOJgnFmt9kW/ZfdgItDFR86N/l/GDPkBS6UE
/hTe+GScQ/QLF6RhueZGZ/2yjGu6DuoMZBK4PNAIevaUdRl92/ZPNA3q1Sw+88Frbny5KvTsdYF3
uTpSo2FnAIMR6+8+DHlsvr65bnXq1e9bwfigb2gfXulDFO+ZP2pLAT2+0ypWbK5OfnvM8KvQVAfW
4TtOxaATQtHEjPS4Ple18UF/F/OIUBhMbJ4bzbO/0w6zavJeXfO6eap8/4yCmuCIpWHxOox3iZhs
4movB7+hYsMVMqLg9xqdFa8OFWZb4MPNdOkCTTT5dJm4sZMvlnBKWa9Ytr+IfhGdpiIzWqL/9/+d
Z8EerWuNRizO2Ic5MacxMQdVxJA3QQAkEw3Mfe3EqCgXuu4P1NdpeurwWPUxj0HmKvDitnZHGSNm
jqjoVIfISUPyT5jygQaClw5Tskmbgw5ElJM0F9u90irRgwTfTUsw9rCzVJ0Ftz2A8iuRQYsLeHdp
3bwXDoAjzM9Y1tefrH5jUpSmkdwCKdBDMphr0TjF6/Ys8q2oUuRtMeaiiQltM1VUhxb5OYsDv3gh
VBqLPFYa7Dz7gepLE2c7ktF7vCcrdl1SuxYr2qTwXGsMB6p2uL1piiTVVozx6FpL4XZv4vRE6g7h
BGReB9y3zsGJygll1RDu3RMUG53GK3GdybGpedfG03ep4hQGNF9tJKchXZ/KE7zEKK1jomStMDbH
yk+oLv0/cykSkHGvw5DcXXp5U9rkenOiqELypEFGMkSizeryKEY7OvCvinTyscK2QtmSIc3dcf4N
+HOi6IdPikwONMwFNMJx7VEZIxZQikgkBa7I5Sm1ZcSUB6ohyAPrPRavttlTS3weKXQcN2BQ+6GZ
Nyk3zaynxxfHntKQa016MNTGailj542u5ZIf+js7+c8lKllKhPmJS3xtoAYFDeFgLDTCKfhi4I4v
7oE3x5yNC33SkujwaD1ZYxye1+3U8pO4Pc6CAeD+RsxSuY6eOReov3zI6uWf1h7jhG7PoyphdaCQ
A6AnYRh5dS3COsQno8x2gNIYhn+27X9Z3In9myZiqKgRH2CxLRM4rzvwLbNg8yDB8s4b6pLud0l/
iTY2Qr0HABifyOHtqJ5tg9hrfmZV4G6DLw2Jj8YyzbcDH1utXiiZLLhCa9ymhRx/puIwQnIFSrMc
lz7JymMnqpkvM1sXy8R+ziXx/TAY9J0MoJa/H1qWEatzF1+3mtkaz31cAj1kJX5SLRPce3jw8xgf
6TwQS7OCKSSD1muCm9M27xp2sbuYq5oh+hI/8nM94hMtfEYJuss9dRlFGw0q49svhQcfpuhodCOo
l9VFtNPuGQ0HLVZus+/ynR/upTgdKFPP8cjkqninScf0tWPhNNh1GecH9qhl/XNXg0aqZoHzkwDb
3pChKePRGb+VSi1oGW/e2YwYOhe+fFMBjGDW1jNKY+W1NGyJe86fi5G9oyz1VXkopcim5LE6TCSc
y3BkGLua2rPAYli4P0kkavQo6waEwIfPwZcd6FjHoTQJIpHdYoFJ1NvX/qNf7vabKf48GCz7NhDZ
FXaqFrNSZTxxvT31MSPvyv/UgJr7h3BStsHe6KiMaS568EEtHYc6tkt4EmHRBW3jE0Jj0a5i0EVC
v3bPuYBuSoMqaNWSz5hjeqmc+udnAt4wMLCU1E6BC+exKXusWetwWcNDDAyXsoHnvcutd6b1KPdl
acoFOJ2Oh8tyuR6L5cv04D5ZGkpj2bMU27PKKq6wu4X29bfIkn0ReFy5HljFhit27zEJNNCuNVlW
R8syvBeGkJ2DDY+3oYdcFPlDSoGUNJsjaxSz+0LKaDRsx9CLm+gVu1oyJNkOOe36KBa3OnALVjjx
NjnYLQsSNNsYnWFMM9yhQyi7fChGhfLkiq8qNZ2QxrHrSLHegEZ/AkcUyUQIyNRGyfK7xpeU53ta
xXZfkyGwSyNSISR309B0aQWczBwrygkavqJ9veq7Grll9XmUIZZSM9IbspsHz9gM/XOXvCI0jRsT
5aVEMXZB/2AOOtXMtIrFKSOgYjKWybFF9yMOTgKjNch+aJ1JLtzMvufRgOClWgwSYcjoWhc2USiW
eYWIKde7mAnm0yJ8hgwJAuc/18i8aUkM6z53KBYYiCoC+ecouKgKGt1C0k0z+UEx/me2JKAGdl0j
onm2zf2/fEkFPm7beJhVXkSCHqFD3FtGG/PJow9V9wbYJ1FrKe1JZ7ft7GUGJX/fZ8yV8SVYW2Rd
bNOJfgxsaDM6Yai9h+UUc6hquJ41U1+lmQ/E5XT2RgU12Jd9m7JP0Kri99q4Pj6F4eNlogfNZcb2
I+knh7GaoHD38JO/K7aCvkCLVLaWTBm7ff2zSMk0XP9oUsUvRqOZRtS3StUR7mFSZOZawpTeWe3V
81xc6QOWWMwNReBXhAGAEUkfhKOWpsy80BIwhe6C2bySkDWwMJsWlmU6S1cGnihwUVnSJnvR0hwD
KJQ+oygslkbenG666h0TrwnSHR6E42PIr+GiG2pKa9VdTF4HeVe9bWrlvKbNXcZmyzS5Rie1/e6i
cD8pR01Cfm/qZsIBrJN1AVnjQEz4H1ZZ5EdhB95I/1IN6TitLqD/2WwcCFpm9bxbgejzaFxzRP8t
bkXUTiIw4SRMKY87a1RcnYbfKcloSh7gD4ntVBPrpx9gWwfI95on85Qz4LeMf1ZI8O0wUUMZQUSj
ZgpS5uQFQ0RzIzOLDvOQIqpMDXUki2gI5OyQObtFVQzZQOheSXn6nY4bKt3ysARK9iT56/uG3Pvl
VLzvzimHnpkqNullgcCJzBahfC3a9/gbYy2jNGp62I9UFz9dXTPOwJ/PsPC1E4hx9Ugr1ETzhGZ7
IAswORqCR/o5D1azqrwBdoXb6e6hB1dAE0wQO97RNg+qSSHHV6OLNi+6qN+arEWRPUK4d88uGHqm
k3owMUY/R4ACddrDosVaXjBbSXo1NCJvsrlURAJrhi+Sv9z8HZQ1gpab3s8fMA7uIhXGoE62PUZu
wlXxTstVoxRpmOORnOoFJsj81Q3Ge6YbUNDCdOsRQPgEJ/+Fb6i0ZOnvORcg8c0s3yhaLbkWQUVT
lMEzwDe/BqxUJkW4P62ir5Fbv3JAyANMu30rJ0oUzlMXeXyoFKKbaqJfMoRMFFYfFgCkRy7lSXbq
f6bUtOto3H/Hjgk/YC1K9FLFsz2P+GOpJ6u2UUAnNy+f8LPtLRWHhM4FzDyKVVpHWwAGxPEjUYiu
LOnp46hm3TPA04zoe1TEvnVqe2chjdNp6kBLdm9RQHz5Kcq0WTA4xzFpb656sS6GxTKMC7E2d/9J
aSX72fNCM1DwaK1TE73QWtq26TLVXULeOOUZO6A4L3LY7fRYkrk49xehm33kLGGFq5yijoEO82rl
qvjEw3pstWOM6JNjkbZ/9JfT22v+fdu4IZITReXraxFdvge99dwnt67eP7VebQNBzlN4SM2lCpEN
donJNeGmER701o8BWsL3K98OKPzpE8gIJkT91qqWonZ3M78MH0OxYJA56umqv52lQb/D3e7pJykO
CsWNmsG4eAt6Bi0uTd5IbCKzz7LIVV5ASbmwurkivs6eZ7IZVb3tIvJnT4wQa/Y7LZ2PoxmQEQ5t
k0WrPI6N9ZSk+C3QS+XjOzZG7Ap3oq7WFAcw3eVHko39967vuySMPphmpXkoQWecJ9bAaUqe2FcY
wzHbJ28e77B7DfEFxPdiyyk+lIZRcu8pitE8dRzht4qRApebTeHECSdxrbIeI20d7COd0eLLTnhM
8kulLStRNrt8m2S/sv2snZYoeIlknymMpUQnznJYSlQObS1JHffOsOIHWivA4bYlm5odiLjGDQka
xl6VzngjvTMbk1P6l1jpF8097TYo8A0ev0ljNvXoWw/H7bmW0w5ngkZlEVY9ZIYQciu/jU56mYwm
zgiemCT7OI3Z/2DsCaDg5gR4n4At/E/UFDHy3KFodgSVhJVLveAUR4clRLo0+peGwnpGDLD/nI9+
9b+1noW2pNhCVN5N8ZBqLjUNzadgoNU6Wdx+c7hWJYosNdnuELYKmD5fvSWx40qQr27/ZQJpl0mh
bpu64IWSsD8wG3yNa7u5rJQWu6CwYol65b+Rk4bROkqF3+eC8b4ySSJfOEOCPOoXZ8VcsFK1xzIv
XCg34NQKpw9Tg/OFfpwgStk/c/JPjtALt1AFyJCjAWQgkNvhT+e5Up89DrerSOUvH4WNMG4HGKNn
5zgNZLIlSuu2iR7Yx9s7WLAT/Nm2/y9nRBMcXoIHF5iMX/CHMWIS5ahTx9jdYk8wlbWgXS1L7Wbm
EJZmfwcRU5ROuAJCWt4U3+jf3lPvqe7M8bEgjmLncV5DS0ShGgbgfEeyjVB21sJf6zy+IAqq3zIU
dDXeCv7w1dMz271o2+Rprn4EUidwqRZwcIO0EzaRKdzGi3xtdZk3FAwJjEkBhBggwlXt/Slr5UOL
7iuDaee1PimXdHkkTGNY4vosUojY+yBb1AZtL1c9rmfucol+sg2NyqEZ/rFeAka3G4Q94681XSvf
1QjExGFyXEH0c8l+BUg3qFups21a3SOhqBFZRqxBrCXsL63HDEj78Rzid0x5CwHHt7aOJDcLlAzi
sNjA+iu8r2ee/4njMNwoe51KdbmuYh9eGlxbX/IGnSSxTQEQYjlprFTCIRN9dfyxA2iOj0D4zo+O
48APeXCehlqZl97G2zUeEalclD2GsEADx2HwCE9zF+PD5UHjDj9OaRtZSFKSfTeVRKuQLaocecif
LwDrguckKvwteq2AR8f2ZoN54ZNvimCJLiaQuaDrhN41DjeDfe5c3ArI9Vf5C21ipKWT6hNtbahW
tXWQcx9u6gLVkgTIA1e+bjk4/D36gE4r1XlirBVn1bzn40uSIt+rUxE5/vC8lapdljTegmtLAFlq
yCP3K4igAdEAGG/XsRh/Ym09ijHpYvrnOLYoyzy2y0fvCw7xWzyoHoZ+ann9tR9jYEXop1rQJ7ed
h7JjhRv+QjKnoYAqtmkv1y2BHVWylXYvY41/x9XL2KfOmbkL6IVI08NTuJmfYcOu8nfcOe/Mr08W
Zj4sDfH0YmtIPCkYO2BWEBh0kktopi265ADjd7WsQvWWRVWr2IXxGBfMfvj+X1B3VeU+/XrE6p4w
TWm2tAZg2MYvbcO5Igt9jO3nrhrunI6F6cWEC9pe3/YfLPsnArlKW7TpISAyryBQRIrTlfUfbXOQ
xX7+/kcJ5qE5qXipQzSoKveCB1cKzSgxWdgY6udwisDtUHiZxGWCiBMR3zdoStui5NxbiNfaEgqT
dpAiSPoxy/0jl98zphyRV8PTZSkrr7aIpoEabB/AejG1oisStQh/3USAtWC475VKNGqRg0pzlA5K
PorhgBOBRiH0/0oHBoknHkSa6rK2zegOwEahPp26GpwSga8Uln6Y9zyAsW4oJywDoJVS96Gwgt01
QsjYW1v5Yyg7pKj51ywxCVW/Pi+LvOGXWYYcQBRVNWcqRUEcwHUWGKK4JMwGBCrVGhI+dxtdBi7T
kVqV2QnYk+i6xKSOx4FarEGuFkXcbK2VICfvyP3E8yVbWOSekUjRk5E7Kz27tTHhDJLRf5HElj23
tlffrrQ3AFrpmU3Hy0Hkbed+xU3TLIct5ZsjEQBKHTEzdb6vQ5vMlvg0Q8NxMZ6K4/7Ky6Nu+CtR
pSgXVfwza1EaH5B0cfJPz7CSG1zYMoqzHBMJ9suSois0+MOVWFr4keIvPMC9o9rk1YiwRP2nTJX/
UxU53lbUNSjdz3UnGlkFiIGcDDr6HGwVcrDPywbn7lmwLsDdlDLE9DhMtEqoCfNHrXALyDtcxtK4
TKRsvgd0izFzacD1A8jOY8WibbSqYnDxB3ZSHvfNigaatmK5aBtxLJi9RJz3CzEx1JUWKJKvb6d9
ROdz9kZfqK0IftzvudkodufvFw0CClK/pR38mMNKEwJxCd9neE73NHnRcfosFN+oDw3pJf8mHW0b
9+WiKIEM+KcYaduOOAZDxf2rCtEXGQUVzQHONvs+DFrs8gK2PoCjSyHNyoST17GKaeRraArGAfQp
YqwMALUh8tR/E+VT+lEXOUgDEigsb0WQz5rfuXOvnSoaSZQdRX47K4wgejO2ymzvhjnG1QKp/YsF
kvlq1BBHFmgrR+/IE+ZzsiysJb+0qzw9UPLhEpc8LvhJwDzhsAI52bug/bQ6o+Ibl9PUlw0Rrjbl
iOidIampthV8P1UTWcN8PPtdLGnm6L4+IsIFer0fOPmw5oCW9uFz1g3oOlysGnHw4j7uNpQSgWPU
2V4tcuT0TjjPzgN1YO+qbPBpvxRMn8cLnXHmU5iGb1a77I49vI8kDrtzD3iUy8kQDAY/v2fXWzhT
H/CiN99D1VKjFgggaridSqMaJiZ03KvWInWQOzxg+oxvLyH76VlLDa5qtg1EvrqUgChYmYqlFn3w
qOla2qfAkekNsHIYjaYMz1KY0y5kngSALl9gEbn7YZUk/F0UC0puwFFt6fV8LfO4Hj5JHx8po4ev
bMiGRno9MIp48KtQZXmFiWvsLGUqiFAHE0OgBrCZKWfyu7TiXu4h8bi1b0pv1U1J6PAhhz9JAx5/
jXFrvjesFUEQPppcGbB9sYKx07PjznuFtC+hNJJsGH/laUtE/YwjpnF87+APAPuwD4m6w8oCu1BH
n+fpZxgoYz7RkFzxBOYP7POaPUQzvp12AMQh0CltnOUE3pAZ996fnRK77k9vozXAEzW+0x7THqAt
FKoXVnG08oKmSrBdOlkw3imZeXdQj5r4/M702CT9NpQpp+C4Iz0KRygv4OYWmRH/4TUc47F77JpO
6mMwgLjcXRJg58jCV2ScTBd1GyMD1Td+csWG2PCi0GSRo+ImgkjbSdBg9yGkJqvtP6QK80M0jdgP
3lCwXmhbntizTxluG9K1DXG3YXolgiI2hu2pmysoVMwC1nCOVFjqiJjAGEcxNqrGdlXnlQmWETv9
EeqY9kNwiW4x9dZof0w6aV9+W08scLdFNr86zfFLV5yBWFzUaRfP6yrNi8BfVQMH2C5dvWIoOs+1
Ho3sDmeSTTV2gFqcY2kBk5ZjSZvkmOEumB6j3JelKh/QzGGITyqNkhWezP3YKN9GXD3IwhnwwORq
I5Vbqj4KDM8WEgCZOtIZATBCGm/Eyy1QHlFcb+oi5YdInSe1KuiWNiv4WmvNKOINeyQ0KScZq+OI
j5QXfbbXyus6aXs0MeA2Tulv0P57PPGV8VZmyFpMUEdkhqp+KpkgsahTWNcgZYpKTdHYaTIKvGJc
6Db5SqznoC6f8RNJUhG+RjGnhBZhrfsvNAo2WX7uY3lo1uk8qUmA0bTBtXZan+Er6Hbntp6QGEzb
Jfdzlo2KcRQuXWoPWh2Qq8I8C2tgz9Mseh1aVvHNjKcPlP8dHItbjC+aYsqWGw6GpeWIxugbtj5p
SFnLpQCOYhr+2mNdQEWqW2SAjJjEZeTVBfGD1MtT8OZO0Fj82ME0sIWdqDncG0s7At+kiuzWoI94
JS7RofugP5shecDmg+Xw5sfxJz7rS/wufRgpPGSiMyWMLaogpTvdkO8tCIBd/XK6ZCR+Qf86TbSM
Djlp+l6Zr8NRGgMBB2Gqvw3YCcqw2e+KMCVxjcot2keejxZuJfKz+GX/LdeijcnpEK/ukFGLs3fq
25H5+rkpri6oeaO0p4KwsRLf6kadLgFQbeyefYk7RTScP4MBSfcrt/mvhS9auZFz+xGwgB4zZ5PY
vA+RdxdQitjK2zAE0xtGB6p1om0SqzOVErDahtIoZlVpa0lv4FmAjlLY7M2CYvrczdYARM9DB7kf
VcbaFHvzU380hsPSBBYPbyoF+yBdn4B2EeXhjhttMbVJxkKf6T9v8K4lejXZnWzg+hjz7lIN0olP
tDkbEfpv2iR+0M5/tvH0JsZNE1UJx/EWJSovafFFUZaW3YEnbx83Fe87MDkmKbkREZ1w3Zd9Ea6p
CXyWJoYTLQiyXKU8nNrc362rvahYD/Vx0NnPm05YtDefVWYnnZAQu1kFE7foE0dfbhp3AmFiBeuj
JN7XmQdCPYwlraty1Sdcu+nqw8B93SSIjZi4WQMGC67+vzE41ClW7lKxTEESL+w76CWVG16oSlkF
KfoF0uTA/srDx3b5JyGdZwBiwwVWfI93s2C2YUijBU83gGwDtFFsMW6/ycAMqREdyIna/e3ZBoMC
2sSfuZNNsLyuxvwPPUieqsMj22nfxKkhf7ota/w9XBHkm79pEtnfL+2kXhdyG4mXg/msOiPhXktE
pMczlGOutCibGyttB5Pj8nHMRkgK68P07cPQD1LGwp+V9dvLeQhHiZlbEesLoEkC23X4nlupKO5I
8bX//oG9aFlMKdeKQlK250YDvBZWkJSM+0PfpGjYZtzRyhph5KTcFb3OefPh5e4oZD2t8Py2od+d
GRnTUlV9FiRIihAL16l+mGaWnZVDbKpmJz3Hyb11AZ5B0NfSgu2MOMfAzTyPds3XCmHtCvGCWgAd
M0H5D410onJlmJrXVxlywzLdLtAXSycbxmMtfh0ghrunz5zJaVj90m+tVIDg5lRzlPV4o+dGugxi
tnvvDzUQXSkClIQh9j1fQmH8NK3NJyJzPHQqdOKRiSgKT5Gq3Yj0GpmvxKoNo6mu5gHE0PdpQshb
DWtbX45c4YfudWnSYicHLgg6ShsQMXv7+5fGxsS89frccmSAOW6CikCDZjjqUjNs8FoYpDoUkWzI
CIZzuDNyDVQrOTYU+vRRbsTNuAyJgc0DxXX9lh9YVIAPJ6k2MDdxDdzAut05PkWZxp2O/J6YAg2m
h/YkFpIt4eeYI/zQEFAY69pWBxDQ8R44Xo2guPeDY6AAF+ic6pFDTHet7ue9PmUUd6sgqFebjEH4
/frhrE14c4vIoeQmV5wSIEr8DjRXUhmnyejHkgRvNRFKzPScOrUR2a6ExWpkpSq97/XKbFN3Cpc+
jR7Heg11EMKSCaTPmR9x1Rr+BDueUzausV0APnHF5bniIRa01Aycf7IU+CccK8LxTst1R76nI9d8
A5xJ6dMj51HHJBRds+2QCRk9pS9JGzUoK+x+LI11kG/Bo1XNMvOkbWSYiH9amwHlMRSAvNPmg25I
pSV4d1Wsu9PXyk9GJOajUtoL8Jt9aqDIb53UGyzJOhfvylqYIUNB0SeXCEcyX/S9sNFiifqPLycK
6Yjgxmia+QjmJJ8LX3XmMxxZLsDC5pGttRFHKP6XVBAIEBxL7pfJ/WOe4qKWXtTWCZRLxwYZrGK0
vHgScVslCj6IqIRbgeP0jgnT/sajaET+UPXXU0eBKH/lLunXWPcR1zdzoXXGiZRhyJB1c8tXi9C5
gnEvXHY/Gu+kCVJlj+CVR02OcpMhgDB+ckRMshXrBNsbRw/ucCbJccUMqZUk0nBiwp3mV7QNB5MG
k0+JL2StZ1idTPJGN0sIJbG7V4tJiSHYsNr9S0t+v8p9ipSal4dgpM28siFuVd+7zdoSNiwCS8If
ZORCZMAzHXUTK3EmlKMgfL2rl7ILNGN+JN8OoZfCGQHl61WHYtufo37xbHn0gMrD+2wSwaZ+q+sL
7Nl9WLwdLGIwPFuk/4s9Ar39X/oC4c4+l/Snu/ce0Srb7P6SabK+bfO92Zl/IBSEaf/ZDDNb7glR
rtAc2jKH6kh0P5UFj+DNtWvpGmqCrP37xufhA5BCg3wLiiORaxzTV4TLq9mYVtvaXkA6WcrkMvDe
n/Pne6/LdI9SsO+96lhcbca4Vrn3o+QmQkTboeabsCapLt4jpGcVixC0SdzieBK/n0XCZbiYfa2n
huArgPkSTO+yskhYO0PoueZjRU9sr/pYJzzpHEBPl+kTTIV4ZT8L+ejAP1jtUB0DQxsN2/Dz1lGs
wDzsB5pj9aS6y+kAY3fVOov44xWHWsVejA9M8FiIbah021g+znLy+HVrU4Q2U6yce6cJcroh9xLA
Arqfle/hyz0/OAdFSdZy0zVd8tamkxrWX2i5c4+NNNNC+vBpmCmqZf2cyybfR3/77GpcaVc7UgTY
KPgsoqhKv7O+Oy7X8GDx2KoStm68fkKb+E1uih2sWrVSJyyjg9iP1ialLgjriLFF5a4phRs0lssu
/ZhEFtg24GanUtPK+iZjYaEiiI2BIdarBSqMK1UupafY8FuciNHgw2+kz4oMv/k+a6eY34Gc9qNa
ozomUyuGIeuw2mJ78PtpQsxxURvA6Vzz7ZTrjtVWOT+F9vUZFdFqCR3349PerFBACPTFAe66DyT1
KVaQDCLtrbfXdGT2RGuNvPvSUFUWY7Yunzko91L7THKTBHPgaAxpiCBh9xaTO67l2Zr0dp1BHnSA
DZ8QOVDkeQjAU7PKkgheX05kU8cP5wTCaooxg3nd5Ym0VnkmJYjDZFqyhFPQn4T4fk+n8w4Q2N7X
KKw+ofehXlh2tx9rsip74eHfcC4LujOPZ+6paZN1GPfYPjIjX3uYLLHh9BpmXUOrVvZbVCh912Gm
R5xe0dzcEq4SDHKhwxCXKkdt1hvhE3on+rOaZJzf8QTjxUS3xgL0qz1tuwPgbQd+ey1fiU9EipWf
WvLHNYQixClFtk2Albfh0LDzA6IbGhjzmlQaSByaZ4Jt/+oM6saMyXRzNQ7l3Ma6JxuxM2cPxPtg
PjuGEHkCvXvV4clOYDqT/NXWCRIglEfoYX79tm6gOwzpf6Aj/8EzP769SWoCBgWnCjYxd3xY+sDs
JYcVGMzeYo5dHWuWod0eSAPe1O7TS9nldEXlhKIQpCEMbDrgP1pTDHodvBK1ftI+p3ZL1Ks5l2y6
pukqKyxqyh4iBZWHdYLVG+BLMM9LLd+yyX9FQpywPZD+fEIQVt1VT3/8oZznAKkU88DcQ267Qm1q
OU6H7unr6piGoH9I1g8vOVD4oD1CN3qpHzK5GXMKnjVRTZTSw/O/paxVVWzE/hGkNJblUd+zqZg/
CvrE4nGQGXgyxQ5JftMOGxRPTMg6kCzFRlhW3J7Xc40CXp1HqaJNARsclxT560A9toBTIsamcHjr
zlIVreNno+0jHo77JQxd8VkCovWTDviF8FR1WU1SMrnVYNQO7YxJ9yKjZiKSzlug1JvrG6bbuTXW
j4UpLX2f12rhR5xzl5BhAd9E2+RBbffDhrw+Ur3r6UvJg/sEA886dGXzL2cqMjejV231e+UDLSDN
UPTcorrF+qxb2ijxpdRGyAgRWrQCz12MwARZhXKSta3PLNe2XNrVtvIE0CMDfkcVoUOSU7VH0ucI
l0qa7kNqxXceYDfGVcRwLNIOY0gBovk26mp2WX9FDw6ZEZ0edQyeeBVu/W3dcOwrKUgA8KCXRCRC
Xt0uEgjppoph99yMmEu+DxdiyT/Xx7eTtlx5TK35m4AkZtTq5vsDkgtCcn9Pnjuuwcy79g24j+wy
UDPAsGyP4nDfNKl3WmyF04C5zzO7unoD3VIrOuSa1en9K/gz6F2KmssSoTkQaVl1G97xJZG9L02I
B/hennNpjlo5mA5geINNL/gr82Bfxcv48vMYuEgeAyn8PdmyJ2uyJPMdYb1oSC+vvA1dZcvyP9L+
potFXgzogKpgtpaUs082DYa2lDB9oGqrZipeFq6YYCD1ARK/bwGWeMDVWRgNdmfY4eZFa2lRRYFm
+clJ0r4MfTDJ4lBY54D256iKPAloEwkWcaeP17ekWbEpReufmBLVIzrqxow5WhQ52YjQFh17Ka8Q
5LT1tU/jewMy/QqAhv/xLdWqSCwjIx6pbdqGOEHm00mVK6l3dJF4p8oNgcZW1/kjb2BAflMHMM4F
8lLk+KwvDhoIzNjFV0ivqzx2uEbd13W+zDJXECr6yFIZURKeirrG1tgWFaHiX9Xv8y1zAgd2YFZX
bw11SyOXm1OjzFyLTZok9Fy9BcNkYwq3mzfv67cNQNNpZr3zvpfPoHlc3OW7VJVtBDoF6TtDtaUS
Mnqev4lL9rkvYasAl5i+v8LC003cdX+TdAZsIn7l1To9+c2KYip+POSa6vwDAvnzWlsBXt14BFkm
UMKRTnnvnjwdsOjwQFOJgMMbzuGAze8RVnFBTrcXMyXrbLkh6wp/57uZ7TqzcWpjcN1BNOW9PHiX
3FLnXgbHVxjY5wXGSz8FdPx94EDImibxx13WAj9yScOuZ2evMLMV5jnrqE/+05vyQE/o5iRzoDPS
/735TRr9HkzK5Ta4qGlkGL6bmPo0jxeGrKi5RMnH/HQW6J+ybv3UNkyEtrCvIYlpWgWuGSEw9vxk
2IP4TKWAh47eK5G0MP9t/vAq8qwE7dWLnUnjnc0ezh3wLattyrABCeNOTxGsfhLE8/rJX1LYtsMc
3LFFp/z2fpn3Ef6DqW8mFwu6w4hdr28wGpRNRb/m8mynCwE/nFlXdaMiatlOmYfJR4b9XZgn9Jce
U08QqmiNTRUdI6lPJyO5M6NYVMhRN7uH7MBmekuvn3HrQZxSbQ2g62P94JXVUbYSHgihc0Q7SRXg
jF7trcDSBeUemFxfexTqCh6RP2cNAwQ1pu6YaxwioaK4C+irfuS4ON4zaAncxy0NJYDfHe4WduGZ
kjcZCevswPfgakm6SbB7P4eP1aga7m54VRRrySLrY15Kj+34dBZuIpN3nmGox3ZLRJz9VWjXM4AO
1jyXYy2eTYRK9wptflc6g5WHyVs3JlbAvrRSGC2LAe/8HMleZtZ8fZMDEanXqVuH3EUps0TXdBXS
NiWNR6RO/MCekBKYFOzadPYnaysga4X7cIhFFw86JQbqOjVovOe5JSGahWg8+fdCTFIgekuDyb7o
zB64rhB6gqIog3qefJpgZbMSIAMr0yqJYQbvxUccafMK1E/X8wJeO7XDxSlao5Iq21F+/PIgprIO
pYwsJDtZsAzPFgllobgzR1i8VpHdhBYNfadij/wH9jhSHFyaB2u+ZF44crZ13zQyCFv6E23gkn0F
bD8zCV6zw2t8sLZsiOifflmyaR9YKT7NvPfcsg4zrviiIzQtp34L1yV5n2h74F/2mWoDb7x5Ow6w
Va50iOLX00wXMJmbX1PPuCYHuSKMUKHIqgXlj3F6RoByJCOKnFk1/C3WYMuEf+h7slPWo/Qad/xG
TfT48IO98Ndf4rWtJ87mslz2DutjoVNRiXW2zICCFDRMzBhmnidjdBj0B9Q2+z+7HDn45W2whqL9
LjQzrZY4A+K4KhG6cJqb4OD0O1IlTdRRWXYPwkDM6WmovWTqj1qq4idonZwXb8oRvhuE9AQ2DZgO
4hqgEhq22ARPTV7FmxwUnoC6WxvR85N+h/Xzxyg1Ea1Qne0mr3s8XT7nCtQtfLyDEikBM9o1Yail
b6i05OHHela2DRsciyQwEAOfSYNZ5VN50Hf7q8Tf9Vpk1Kcw+69oiGBRzyMW6lLUL+e2dshBp9ZP
e60VeHqnYrd0ZWs+B4p7ZJqICSVwdym4c4SKangCqYl1eUtctm0D9PuyawMV5YZIodpVAPUP39+J
yUhiLM10qqJwsbcyJ/H10djH/QGYl+lJlXuJAZsXIfzaE+//y21eHPtQZLpGYSsMKDH7VArVya/M
fyEd+NbxSnP/Jnm2VUdrjp8pdGmK694ndvUemCWEPCCXHZR4JIkFknubHcoGloDy7MtwBjd42uYA
0OBtSsGH2RlpVs5/MG/Y8kmHFzntbVMYUjH+25grl65fPA8saUgJtcRnXbbx37PcW3LUJDjGuNB1
CmOoEGaT5HSQk0DtlG2HWfWSsRbVAbEzbXyHE4ALeBkxgi46XCMnRmmR9nqe0BSV617c/piTHzWO
7S5XatF614p+1g2hElZmZLalx/1H/d0bF5Y003Qx6NnEy0a4flgylFHEaQuRf2suYCy31EOVIymm
Ev37eq+Moeg3IvSwJS/ukJNwX16sNydO63ihHWXn74KZ7/pMTI4ulMKczZpRru7qnI++T/BHx8dU
x4ODGk6lh3+IwFY4H23dgE2c9asbAewGm1JOhHXZ1DKfKv1RtyV6F5Y71tbKiDhXaF7e1LsTkQeP
i6YBYFNnaa+z7QVqxAixJA3wxZhOCNJHjO4m6pyFxESh8ziukxYSKlxx1cUSHZipeaSTVjj5HMin
i0kAo+FvO6sBn8V9Jvemm56GvgFlJjOTxwALkOZkt0p6Yv5ym3GXnw59nsrJWFYzWWcr9tSBPpVS
h+ZzZ5fzD4DGN7/hgAS/yRwqhzdTRkSYZ/SgsWth++9o106BVBdh3sm2f4ELpjo4kfqmvaHPSXbf
9zq71lDqJTN1z2621sRuGgP5Tm8Fu5ZzujTbHHCTj9mtfKlzz4ReB9Pqzl779xJBCWucCA5e16F9
buh6gldBpl0+FUXnHHSjPQ40IugM5AbCb2I6Kv1BDFEaEU7rtZycarpVVYFC2Me5SkWyif8K8ga+
k9Xb0eltNAhjGMa3dIoc+VkwW99rS1oaHVCfpp2ge6ndY7GTh4kc5fyvAOeaY9exeCDOxLO/6Tig
J36TrqQ+4/afx+BbFvSvqi3FxTgTihPvhcdwJc8LF2OCgxbFTwuvgCpfoHHZWQPXuTatZ2oBYLS5
VQoSzeNbdF5HxNkow4jli/BuwFegaXTdCn7Q1u7qAgcm7Kq5h8B9XpoUuqzA7khGgNUCpNq9NIb1
+lpuVDI9b1ZkefsEQGbNCpgYImjbRqxlQjDvZ24FmOCD5U0ePN/MAU1EtEFgVuEwUMynI63Elz7s
H+ncGaUQF/HyM3YzOXUlOMXi+YEo4YbeksUREvbG/ufvyxOnalRtEJL0naoPjyxunnLBIaIxMG8w
mcRyQhuM/ic/O2eNj10QwA/jo/Yj8jsNlq5pwmOXBPVMJcWuQtsOLoXkUgzE6bjWdFDk+saZN80m
hVcipRdiqHr/H77Lf8eg1y3dlrhahNa588ldP84RhIA1LPMz2+uuZgKBgiXGrpOH0fuIB+uRGsjM
j/9FvkJzoCPfXm8QNkdIYiAajPRauevcZauZwKIeZC4c4gdotakV2jUecZOQzDhNNrM9F+ghHe54
f67cNOMr4zifBjzqwBDs7whujNl2pdOkPUq20O9HUl5RxadrHKFNXaWxcbRiXEYZgr9iRe/n5v3t
TCh6XXva4fUL3LecM596nABzec9Kw90TIHrTYq9OSS+V9QMfUXM8porPOYDv6PXhrVVALdCXnkWb
iuaGxpA0igKATbUmYtQ6aIlQ4utchl5dvT8QA+yhDzKRLHE1FxxcHtmpa6x3ah2RH4L1ehlPIJ/J
k5hUozrmZrh3Yvopv1YJ1N+VjwyDO0SXDGep9eoDlizT5vWs4rW894OR73uDfDV7f4oc0nTf00qo
uEtnUj2+zmgixsdKw18+95ipzgtgiYoNTbYVs/uBkrcF0VldXFn5pCDE3I/q3cSCDm9B0si+JmTC
3KPU8Co/DvTS2kutdNJx1zY9VCZ24tY9zthx3uxTUaMekpzw1Pa0GmWCljkBFuByMwA5tHy+TAnS
/aHwDUz+INupNGDf5PTZ1bfiaq6kqLswZbuOc6CVAXfikEeyqn4EQ2YQRoTjKBkWQXwWGaDY40qR
2bQdiWryVcXonkdSdWHsEaQyRQ6gd8msXX2dJhloRxI8bKwilDITlLKXByogAn9yd/Dl0gkRx5uX
jRrjbjq4h1f5wqVKS3Ufg8xWpwUVcEAMTNuzYlqdOeJassd6G85f2tUdj+Um2iFrizC6UdgZM8wZ
zHCAz4IATSOVv30YN/+/xyJmN/8EzBI/SehrrZaua0iXyYplVe2yZprSh3WgG6CJHJiSN4ae14hz
z2T+kIvfIWrUiGc+fhFi/p1XKgk00s0fdhmWQcvfbn8vBat75ybDojdbPlmo+jd2+1k/78b2rAzL
aZqOgbVklZTgkeg3D/MtpT2RiF4dPhN2DztHxKWJzR6pfl3HwZ4hYGRp3MA/DCOBqsKNPWWpd1YR
o9dfVL/sTgj7cozQoOdN3WS5X9hu78htBF2BoEUo/8H8LrhK6vVTWKGNc4oMMHw1T7xE+9nr26uX
G+8NhSaQ5DCQp26a4k2Y/3Tql3xRgbjo5AcQNKrM7SnwZbr+onM9UlfD1GretMkuM8MWjxhQJ95w
qnmgbWV42HZcnCHRpFeEXSYZV9YilHa/z0SG/FXVlTHFOSv1RHIIJiUp/PDY83N/HF7RfqDeNvYm
RZlBzOjf3i+BCFOaxknlHYnDCWKnFtmo/swEqL51pYdzFS/08ZHRYQiR5NoZ9CfAS3+zOJmdBgF4
jPRx3DMYI1YLbUtUA8SecKf+KMtxp0mnoACQbJNsW4NI4TTwXHGQK2tNhIM7EboYgIH3XDMfHlwm
yMusO8SSKsSzU/wu0ip7J4JK8L64w2QGzWXWQ53XnMaqZw9/IqSpeclq9H8K4Adhxz5qVkzIgLPk
/Gz2gi3tnMtu1LZoyp5rsRjR7+YtutwA4tQ07lPSaJiou9H0PmyU5D11zGVEETZ3xFjgilk6FcE2
oYR8Begil5Pj8DmZ3aJBvSoT6ddAzOEFiikwH03kOhaEvBtGM+me46+hqG/LUt5xnmCs3gAdXfQ4
GmICC90lezmg7yKMxNknlxRnPh+7q+KXxfJRHvqzWGcnByC23D7wWCZL0Ms96HVW9f2kFvXDUlOP
HXE1AhNCiZReXu/dlecn4Ai0Ewfc0EYgSpqIO9DY94tgWB/xBmmO1CEgymlhJvm/BgQVQEOeQJ5B
z7NNHJ0vNgBdoIBL6MhUvM7+/mt+NQUzOPYvk4t9o4tQCx2esvN0W0iPnVcGcVB6zPt/+tr34FWN
kiU3A61slV7HOzbhYx/W908YlcG7g114qA1/STfTvEaTRMiTni6l5ypVwfpg0/wwfFeZuCq//Fcw
OKAKI5AVinqRV/l0gqzMrppyOTMD66OWB3FH9evb3WYlWZqnN8RLGFR4UnENojQ+kgtCHBGdiewJ
KYFOnbb9Ldjmz4N3nFwY+6ibwxztsCboskXs/jwTdEiGu9F+Z8xJWL9J7I1GLma+XLjbayPg43wh
avgyBjIoiKKSnqlEYn/jOWUTelYcGIBAMA7F1VtcFe3qxj9BNchgZESXYVEEUjFCjp6L+8XnEwDl
rq8Ga2icVb5dBGzZIGQsqPoi7WuiYQTRPo7lzefyeDfkFi5NhXunBrnyY9wIWPwdXiKoHruoGdAw
7+kILyfEGU2dUQRES1HjPquasNAaWqX+m/D1wFKGLJ13QWfanC362iD0iYyOWM1BPpZ2JLw44p4z
mXI3CdHkAKToF3bGuN/1Cbx06V5aEGWQcxMtGQZNLlngZ3iKrCjN01u/ioviCGpx6rIX9C8FNriW
X6KRV1OsIYhTysqA/UpgrieuHYM1oJbvLMc+/ahPnatPKcFjhKyWEeGRKSM1j/BeZZ1R/fYjuWXH
FxO+RJCfcDLryBQ8CTBNuXfIWKKrRjpuRQXyy6tybqEccjx4x27Kw8cIJlXjsOcLsG84/pnh3s/n
QZ/vsZFYrPjmtTMvlkn6wvOHrA6V6vOszQJmVwi1FVsbWtj50e746fu1JR9hqUCqHLW63vtLTjt1
4zq6gkIt5u5vpZVBDsTb3o5274kxhcWTNXmocJ0pbudtZGDllBRtXwxqIlxWtXrRR0WZhgA4gcAw
ShJqZrm1DuoNjRTGu//uYA+bayVD0+sJ8U1SXZdK0zpaUYndy+TUoaPH0LXr6G/XswxVU5xMk4wU
1hMBG9wim/+Irq13e6yYYaKnfNtqcvtUxHlV+RBh0gbe2bkkEcFEkg6FdQJAcP4WYyySAy54gxvA
C3c2dwxNW2kVl8nYyt9vNPxv3IbaP5fUq0QT/FmJfliPlhBPnyXSiAgYIS43kH2MLNCrvRoa5ZJN
DYBnvJFlKr8oOOkA/AqIQ9gthpQqgObBmPNsCSz9OQRSYXqPe19v27D50rA9Q0PTiOFBVHpLYnFd
lYClHUEzQf7CLwrs97FUEFQ6i4Tj7hOJdZyHna6HLf3xqZdHaIleHoLVNCdzP4mJ4BaDEqD/hGRq
SgOHU2lorpvI6D1ZY50L5iU1xcTM+Sr4SXsLYYmKEy9Va9jvNrEv+qlsDw0oeIm15lnCwsImVqvt
+0p2mSFNvAA8ozrmEDknMYqfVNEdbhWb0a82oqhegdwbHM69PpuGJ5Hno0ru8lGbRaUmehJ/vmFP
o7aD66iaGIePt/gL7mXaAkf7DmMn4PNI7rDAKx5rKU6uWnyjjWZq3eVpRFZeFOEzB5bPDM/NPz7w
sm6HLVtmMuHinXIP3utJWzelXFaMKIW98b8BYl9oc3KYP89sJl8SJVm1ZILZf8POUNBcUAOTheLD
kjJMBWHaPHrs081RtQ7JUba5wYjWF1sR01OYALmYYPn3U9op4ABbL1x5HkNGq9MQt2ZTiSa+VnTJ
u0OPZsjHlQfgBTYzdcN1qBbOUPTkLHzNBm2DOKoIkxykFqu0J+xMCaMBDh0PtPggeTz6dxiBN38m
LPnTi8zhEmbRyYxNsVqG35MurQSc7XR2SGJu6jbzBLXmuv39NNm7AYU0eidg8BRTU2XpXM8NTR+5
88VAdLjRuUArGm/2L98shh5/LNWu2f1WY3pT3NU9HDac3txtMjosQohTYD7Am+YWmOldHFk5RJ2E
nBTQgKGKy8g6kFEmEldySLF/hot97s4H5atOa58oSjXApZ7youx1MjA4GdcIeeuCZ/QBHyGg1T+B
MMrc0rfJBMvbf/IJhe5sQchORgSUsH7znlRZ/UrDavwMy7/4NQySRUL+GGTxF9vnsSzzZPkxg4mc
Y6O4ADARY7XIU60gv/6mS/+fDhRBAvsM4uH7ogDQo0u4s31uP1OsvEBywws5M/PAn5tmKUOenerC
IlQHQ967d5f4OlDf61upu3XfSKlX7rLryArHZgSRKyaLxCeBxFOBngNecXPDODGDLAcUoL21yCS7
rDJONnlcBCJqoK3tFNtrcV8OVVw7zZWCvl4MZgjJGeICG8uDiW8FLIU4aOH2DedDFFS3Qz7yN7Px
qNnoRSeE9NkaYGx5J79ehyk0M1sRdDHAIIIYEpmu6QMXY3sM4J8MZCb/CrYTTYbzWlQ1OE/NWfGT
sQXw4ovpKthMfaeiinpLoE42GFohU42SKTHhHNExu18Ch68T3/qCGFStTIPtka0gPDMKTBzmiF+C
SGCmNqfJ+3+9FI0pdfrjULB7NPZd1F0Uu4T0+MY8f1tlUE8UsxthF74kI7/Yjj1gfXuGtjj9bkjR
75m3cHg9x76sSlSYoOPMz09uqI2f0jghVV4q2U0OdCW/Dnitix1EwVHdsYayaKY7n7FiOvGTGyv/
tcHTTMDSvLxGcwjZMxXaw01xAOoRsdcHArfz9o5CBvED7KEcmOn8r6ivnvCQokWPPNYCBPYHeJJ/
oXvCPO5EgKP24dPcwGiBQcF/4qk2gYlcThUDVGazFIg7Z6S05x3xCZw/HEnrbB7dkE5CoXaBKx8z
P1++sOc6aBEP5XNC1GZKLlH3HQ0+soWJZB6ADzTwvzY8hWuHooxWCKOKFJPhzfffW2fqELdZgHPo
MX3gzezzvtcZpqBRXRF7mbL7ZvMeN4WOdmCGNRnVylgHl/xAMtyyHUVeD5SlK2ieZ6qzNVZAQp1+
N4/etBP0GbgKMsZarANF4LhN94YvNWuV6pQSZGyvrqIcfc7b3oYUrn0hveSBEH84K/2WCyRQogCd
m6+G08Q5J5GMR5HM9t5ElDmZLPGPgXGcqRhHj7x8/brM0R6AyCBCTkD+WKagbnXzDvQ5Ww2iywU1
15yPgt5oJI+PQw5i157P1b3sQ+qbiw0zfphMz+lqQ/FwZ1oVRgolvsyzGjbCTS168oOp65Q5SMQX
7aRg7n2Zo1vnG62sahP1i0qlRHgKOSITCWirda79AFvy24C7JULlFmsT/vd/bOnVRiOfWZNeQ5Jy
9QsC0FHA8eZgTVbM80pdrzR68uaBv67ihMa4gNpATX1lw+tRRXRa9fbUmbaT7tEDjZGTJhO7GvX2
O8XAfC1XaLOM6LlGboixgAV20CI6fAvl+gj1cjN581fLgcY9z2YZBXwTktNsiNrAEpkpvnmtAe8G
2RBJLQtqCTAsYuiWuGhFsbptLM5yz4uLeFwFy1O6g6YQ69HIZWR2gxKSYbjkpS6KMMz845ZJA3Qj
yKzcdVea59aCz7F8U1YgZJOpBskSBMnEJCaJ/TMLf5dsSx1n2gzH77dkUS0KTV60CsTx+wlE7xU1
2Gi5SV6c3lxbJI3zqw45zMQwT0gYkduzWx9LCJGWmYt+D2qVn/rt7sPA4HgXIozKejaN8A0hCkOh
xURIUexNr1dPIP6AiW2VuI1ch7M2xzOpYKbBmBwA1sZ9hQVwQb5LRbKYDD3AvbAFvnH93YRqc2OF
/LqbHK//JuEUyojyTa6tuRSb2/Nskino9v7pFszv3bhUA9u4FG5STbPwgZEnaacRbzw4XMkdb4se
1gC+wzWeksoYJTAPhpi6aPL/vxU4pSXz4fdfj5KM495sJ85ULjvGsZSKWPeSL/ojsHgoparj1rHD
w5zr4OEB8b+DA1vOzq4m2E/SYL/a9kPrFAWJgE7gL7Qu2Ou2U6kFo+Dfzw934PjfJ3OZdR3kQf8S
JA9JhFprJWbqqdLQ8g4lrbmj+cgMNWF2yuPgBdMMUSz6Kv99Kr0ZzBaoWv4SJEdctOUO80z6EfVL
yJFvByijeVtKoIrKjcpmi154tJN8/IjYMkxb7/d2IIU3JZ3Xj2M6QgzwIZ03AVqv2lPKEmAESvQj
U70LUugT3lHOrer7Pgj4FAWXKRmCNa25mt3f+ppyekZt9taUNRIqnCHLK1NjmphgSugM9Nb2Sooe
/pTpoI/R8+lWsO+R174JfOLe6f7uqB8hL+ypv4OwPRKeJKlJLl60LBpcujB7sk+X9mn7Lx8HFQU/
pCepAZba0LWPOnQultSuJ0QY/DfxQHXRlkCPTtjgX5+oTtTQ+iJXULgEXFvRSETAbDCSfL9guk/E
2E5kahKLnOT7i9UdH181hkSWMZN5ZMDDoMrtc5r481Z3KzJ0BcnvEEa34rn/WCOWRmX/JqRTnUlp
tDvJXotXnGTErVywounloujJvdgZfzEAOC7beWfoyeD1IIqLxSdGNyqKwXIeUKgdyyG/as8akXb1
5fRy60qsa7JpKDoAPxUjwthR04ZulY1gs3er6ZUimIDSb/FzR3yBMs7d0ZXTcINy3/iUPYKN+wrx
2w4LnSbMyoMsUlQmiijiXCIdHslrsBppSYi0Z8jtRYkjCqRTJKvtlxl0C8903nwQRME4qPlJLBfl
m5jbclklBYuZ4jDmeb67ttbHndMCDep5riIVaaTlhU7ZJZraDurvmuENFVsa3uI49+rDF3TNXeAd
YNGcJL1s31kwbNnqCO5Ml3eFesFPNFB0NYIj+vPNPgIoX/nXWxhr0P/oirQLUwYKoKvL5k9foC28
lQzCqyO4b2BYtk6lAotSw3sz4BPVg9Jla63Nhaalv2rIDJ2ovYqLDstg93MFPOWAFiiDRA+gPsQs
C3dlqo/LPwhJg6bbDNPmlpHVTvbM1mJUUiBxEQpp2qhohKztMOu6j74zwg6BWV2/phIKwIOj4NP4
774X6P81PPzDOYMPqyiXfPbDvIRvNgnLv3mMnrr0vYNQ3IthKagVqtFtpklgj26tptOoCDFZ+C0Y
ccn3pk9K6QFCh/nuR9E7IGSjmMajKreuMdt4QicVuQLnk38kWP0xu/mZVP8A75+QsjDbIaMrFYEk
MgcZal+m20hvGtm7lbc05RBYklUvzKU4a1Xm1oIp0atpzONhJ42RsAlcRioZTq8Y/9p9aUVqCP98
YthWAW+sDFa37vfy4T1hZ5HphmI+nK/HREwy1klmu238s3JHIOtYl9MJ7txTaW2Piq/yi4hiZ9i4
ifDq2IpVqUnMug+iciSt3sP1TdNb2Z0j4uBTiQli3CbvkUYfz8aFoF+QUuoaQnJS+My0DhpnUdUf
syKOLK18aKLNw8UOSCRA6myWOQ9onswPJ0hQqqx4NGjwDFVQw7AqIVd4eQzaVty61jsjUTANBHk1
ibxD1sa6Ym+DU1ZqwWsLx4OEqHOb76Qqj26tpJ/5bsheog734d7zOYuR6SCfVr3TA3SLdVn2kmLw
gjexvJMol+DO1e7u7h6UlrKDUYig4sqACGv80y9FKLWQ1tDi1BJuBe7XxuiJmwZLuPPASymxzOET
sj0Ngeq/DKNjt/iOzcysuahIHZ+NbME+Wq6+Y74WQ7SRSyjn4eyffRkdl4Smcg/orv95JkzSXJyA
FljxCdAr1hlxqmm/EC8YKKPDd3yV8Xgwcta7tkVLiqrGdA2E4RsLwg6/8LLQPaPAJ3Vq9UHisg6M
u9DEdMRbi5f5zO6IYVd8zozBzWzHxJ0wqnhwZXVJRj2DG54c9bMnaEdhOWtePMPOxbhh6+9e0r1/
r97kIU/23taAb+9CV3qs+Sn8U2qJSMDsl5ybzWVHD6HLJAaantJgpD+bPVCTd81QnLT0ckKuKdDB
it9/Y6iyH+0nmQzcQtDkp6xk2N63RYKsCSwna5WZzb+CkqfK1yePh4SQi+AeXADENEgImrm9ai7M
nHj1Jl0G7lMK/KXT9fao412sqa5DW5JdmsU+YU58jYQk9NYURj9S8yDloUwJp8bkNERRc9aNfvbw
tC1kGt5vSe79fm1HaCYxkcLiSOH0U+8Zu6WRUwHfuIuRzon5DMbei854SDkqf7sKtbSQTTegV7ga
kEY2zcKubXLYDLMuTt1Ti0FHCAfBEn0x6cytMp0DYKDTZ3dpYphDXhKreKU0VNaU6P++R58FZ71b
B9kq5V5nbQSVMXcZ1rpXxHHrmq/WubIBiYjiq0T/9ltvvhLpceldiW2CZSzNfbP9Ip28IoZ9LJ9P
wLWP2K0Tci/7xKY5ErVjWqd5/Toi7XmXGLdOBFd612SBaJmt586Pku6jJcscfzr/ESBZWujbfYii
WO0+YvRITJrmqie3yGGkib0wYL36zaUE+LgEgPq4eNvsWjFmm+p3LXFX++j7BAjFXpgTPcZYqjJV
g9AvHJeLK/XIM1fdSNgT5aTDh+AoW7U/g8ZsUGhxI69K9tItJL/IfMj1mB8Wv4yIZ5YVY5b5n208
uDJovPzXpsAOI0ookEUmaOCne10L7w0psj+dLXXifAam5dtWrrPnZgmn2sMd74wQi25pNtKjR0i+
ptxzm0T8MlZLabVhheFTKpwBnpbvcBgW1bPtiepsOpCSxzKjGtX4QN5vfnG+/Xci/rB7jcu4r8UH
/xWNRKTACj15p4fApyTA7bGyjErfx7Jg6qPxbeT9lJQGRQvpXuQIJVEbGMsHcfKSO++H3BhH9APw
Yv3YDhCpceG2t8hYyRpiV+R1nVR2zk0rPTSlJURFTW4xOCDy6/hU8OUWD5Ebeq/TOxLohceU2iLY
qFK0vsKXuzTjhQOVRim+8Ivwz09AP3DrlxVn2tWsJVDky6aOBYwxUMqdZgyg4Kt1wJWoJ2HOoeGK
ubGb1fDwzqTkX5N5Wo87jx2Fwlxaa/XQZbsaMDxlF9B2M76tKO2k/V2REOBttLjfoNqEdvjOlWoD
k7twCIMr/lP0FIJIORfQotqWA1bFvKDZIXo6Z6rcoU1tLnVNU9TTxW3GosmaU+O231hfd35OE4a/
E8xpsU5+iyO0klU/lv14u2rL9HZ8cjl7MjxvLuDuC6OGskRtjYXYa5bxYqNOa/QiGmPB02XY8MLr
AvBK8fYg0h6202x1HCjCKHIWR9IViz/PMiepghizkFx+N85D/+LVJQLBWsCj6OqA/CouSksTqHNk
PVQJ5kzgLIuqyTbvgaSHLjrDzc+/ae+SVMAPxYVNV86ieQ1HUTE73d6q3EYTasK8FBX6noGdKjit
CRG0oBxx2FNhQh5PsnsjPeHzVoSgEzXbmLXNjjWkDTQDSDUxL2p3GF4iq7tlFGqQ3XkLsHgr/2bC
4nePGLUg18W1/rqg1z/UxUVfF4kXuaGVAbzPCxX5E5/I95AaOh2dY815p9+nP+tE74eAFGFSPSTw
hWiMNUS58VtnyA7F4p8mDOcVasqJECs3iKupMztX9lFF6TIut9b+/yOzBTCGij/ovhRb0/yts+ny
WJjiYXhY2+1u4ADxHVVtVr6LXFiprot2ySxSaYkDe9uMjhSc7CvEr1VSPL5rG9tuzis/yunU6ku4
myeVW9ap9P8cFw6CVabPq2BYxRGs9M90bdWZ+RKX0RbxORFOFs4fxrUD9K7jeMLxJwuzdSaYAk+8
Yir0ThzJ0K3Cs4qAAaGimiu/4TcaR27FRpNRGa/LJPWbTiaBeeXNtMOHyQSW9xNzYs8p2P2skCOG
p7iLc45us5vM4sKgkT3+9tSDQYGP/4SCAids6+nO0DyLewLqcHkcLDc8dcq8muanG3U4ncEV85M+
zztPNrCKf6KLLek6cWILl/sz3VPehbeOB+KXLC0pqbWYcnDmjtjwAm9rcdDgS1bsbMvoVkVU9CAU
pp3y1a0lEQ4OqLPOYSh2qv1skT37NDNpiDryB7BdrCNxqSG5i6dUTQjWHYPmb5bw/s1LHax684So
GW1331UCpVBss8RvuwovsJuEbDBXJsb3d62aaxIev+V+RBJnG+9hIDGiM2555EickO7oDSAirPaT
/lRlYLB7BGvcYm5G7x0mxBGJpIUUoSRk56sQjSK+c36j7C4WV+TjSeQMIZt1x3ZS/TG6X7j8kiFh
dUaE3pffrYBGHWKM2ATTRXTraU25NgeIMFY+0pak4mxQl5v7xrEs2T0z62m0h+vBPG7hKKI06VIB
DPw7DC44aaee3HqJnNMWcc6IgVnl/kw5b5SpAlmV+D/B1nIfEmYFIKyBPr1KvzSA2+sHDBX8QaOd
7PVoq9kFis492CfJmnbAdgU81aHsE/kqp4gX1FAbMBe21ij/m7aAaO/AR1hdoFeRZWrEvYpcGKUz
iWH0j/bkpF/UA0U6DkbkCqhyxLsXpbwe11noxY1bHJqmIrgTfgDFFCkz7FCOkPSGXnlVqb2fcG9d
zU3zE3qGTV8lIvZS/ghBzTQogjcVohme+c2qbn0ROMlhXNSjFcmDzkY0tsqe9wxjeJkBB10jS5y0
iHBARXJqZiaXpKjG78XAe7ydZrIj/AsGTahh6TlAEfL51S0oV87YGVZ9kabgbcMeDevblw7wHCjp
dKeUw4XH5qrcBZY4vmE7OifcB0VSoISbXnLFaRDl/ZmWcXcE1F80fTBfykoWNaaN9Ubl62QUIv8m
CFWIKfCLDOhVsI4EvAOkR+KhKhGuKQ157LrVLYrA+RQt8AUK/zQipTtAUfX/wfjv22WYOOG3u8iL
FbgXtVUWDcHewFsstUYPau2T2Y3EWI8JlRkQYkN2A+kEpRs3J2DQw3NZ/HmlVpemz4vObBQn5WZs
F1JtmPtsunCidKWT5M+iIhmoonzf3xAD8kK77ziIE8fkuHnJqldkmQYO9/vPg0phw4k+FMwtlU5Q
j//oX1+cc+en0W+p89vbnnv+SGfaJLtDCNVIKIXTJfbAGoUbCjTbTY0PcUreWWbQhQOdIaBuK0wc
OGa2Eqx5vGXDi8WUnAbsycaLuVI35WOemFIChAo/xjr+U8wIk07NtlFXfThU1iPUiwqJgKVu7DpG
o5FRKGoNf3j8adfS+tImic3zy2IUmaEX+RpxRGNLuv5fXZVyryKNp0CWzSB1sqvX6mim0hHsxG4X
5ylLgEBrktiHmx23FltqoCpV8SaMpHy2inmcuxaDtFaAnCW/+Mp0rmZzRi79npWRVyTAw6af6/KH
kJ+a/kDw8/3VSmi7UeqlVLvm8jPkUyFlfVS2WlJTT+cHB5jXRoHBXUuX2jMiLfmSJxCE2j1OjXAj
FF+4QwupeEK4SMPJHJxsE0U3fWcByXMCBc00wvuotL+7O/QuGAPzTXsQrlKmVD2UU2oP1JnNBPGS
M+wUuXmFz+VgvGEfe52/NgwxRbzIngGAEFT9s9gSgXgJHpjehbHRf2jqUURIBih6L0R8c0kumsX5
oG3iUYFypmdesJtX0CA2c3ckkfEes0akh8eSPZjNQbaSW1d0/G1MTwBajE598B73SWmUntdFomYr
b0sdRR6uGCNYdYeLjRlWkBoI9PByKl1tsuFXbnjN4wR3t07Lut76DOuUbciaMHumQjTb4I8tfTOO
WqTd1Izc9C+tzLxXIzy8Hyoc0icTqRLyCOF0do5BOXk9vtVrpbquzqKYkPqcq6g7gKpA1MdVpsfR
IB9ya5GFc0Dvr2Nfc0iIZqFB3eiRnrWtXMrsUm/EHCjNFh6/Wii65PcUdZl6OU1Yzaez+Tcl4st1
rQgAc5asej3D27JdHsA+msODl9ExrUxAkONmIrFkl8Nj52KPlfbj1IcCAQLhD25IsZvxZTbepmse
K8ewxkRT55mSeKCzufv0a5Msz9JLLIxb8Ykd2msAuL2lhePfErtPskUIejLzWMZexs4hAFQU1DTx
6zVwX6dcR+E/1bQ4aMvW7xp5ZCH+rhOn2RKrhybnyq/VFLpwAwU/C5uZAEPMd1A9BbwXoGQlSxm0
/lg0Tx5PaU8mtsYoK1Y7ePMG0Qjqfr2UVLYL2Wz2Xb4KlAzrIKsBmW6ntHSAfAqRRWJ0ISHUZp+u
gHQiu8L4COfs0QE6RfNeLuLqWzGWvsVv7Zp/XB9wS9rStt3Buui9U7ufNRE0V4GNG6495EIm74Da
2XZ3KgOoT6iMGVDeb1suE0nez4YgAttc3FPrGzKby4Dy5virI4adeiLsHD6YkymzgHMlfoxvksi+
zSTeKHKl1oCNpmICBLJ8v7wui1E4W4XXjTYwMWr40PT/8NbHta+W82SngXmD3tASrAC72GoE8C+Y
KHp+trOHUYd/GxuFs9l6KO4gRIawU771QfWwRSa5nmMymF9lGcePq4kbi0kCzAJSMH5Z7DVF/ALF
pzuAUl1iBIYxCeoKSo1Nm5XKm9y99fAct4CdgwfG/yhEWQxRnkGZyIZTDVJn08bD5oxTtNDbnWZy
m6zzIrPHDyo6FU7nt0VYwG4ucJcmpN5PzBP2zmuiSZ1J9QjNnz7l/Bsh1bS2Q5u1HeVlKeOBQDkc
fIGefIF0pKpgRjwFF5Y74ROYh0UbVtf8iwk3IQx8MBUatCvt/ciobGlG35k3xINsp+6gZYk0HR1D
o2Yva0f6+tKZiCvX7sW+SVWGhLAi0NniqQt873plMjwr1Em1FkKUWW1fF5Y9cWrO7xxsgI51R4XP
slaEKko1SlzoXKCbyyv721qxuVsRd318XZzJIb+Q8ynUsFTX82bRd0gY+A4BfsGHX/P9c3rBeeHH
6jODGGYHqHkqBS2I4r3F9R8AlFAoy5NoFi03bifDCi4Nr+mYfJGetnqkHSBy40FrGmsExiC0GNrR
KZbZdLCNAJZiiYN4PMc2b0TAQ+HqMBRhfo8pdbqzyQ1SPVqTmkbJdR8t6JktVy7bKAWIGrO58e3M
wRcXvet87VW2nJ/HPX5AjwDHaNuHlpXwAa3N/54pEEIOCgwxjO5EH6m7Rc1xvWeNxTrdzqEErnKM
YSyDDqfbonkavgNp+1T03LQRymTt09ABAvUEKBa7Fq+yWHc9JQBawNXZIU5QzwHGyTDZxuHaHTnt
hH3N+qKficYe+vYXTakLB/QK+20sngMhPyEuIVVEWuTYdcXzZFDgVSDE5hxZWhxf3NCcjmbkeRWH
92JtDfwAafdUB5Nx6F9e3HF8WRXr2B4yCPyYCvVGL0uaaj7CHOHEdzUxeiGVqb/kzU0WPebQr7pD
DZyHy1gde3/W1QJ6IuNWsRq1pgEVvHtXuz3jbdVIqQmwkGVgetgeXI67qSe31eTWpylO9qASHGFN
mCPGmL05scJrpx6qoWAE0MuGRpvzlBRj2uL9v3ooF2wjByVLLiqGXg/q6Hb5FAcoDccoqKSOSsqy
YMumHgL3wblG+B67M2aGIg7SJ7oJ64q702/Pn3gbMCKo54BW+2doW6zwrhb8Pnhlj9wKrUQl4UJF
LDWIPU/h0BMkBAL9DhSF609Rhmm6oVm4EV+Dumw4CUG4AcXtplB+A/jy6tRK/NNp+Wza7ZtdyCb7
kT4yAZG8x4MCImC2ftdMWcCP+pU66BrnWs1Dt0rrGJzbIOL9HIJiM8Xql/ql9wv04/WsMmg2FGck
JiknlfM/oXNzV6P97e/nLTXab0qSe+snrTDeNE7NMWvrg8SKkVyOMCTx226J66GK/3U1nSoM9XNk
I7+B/llCzHkxMwOZG98QCayMax7TNGbujkVaB+BpUOKDc73101rN8Gn7TFnq1nTzvTgxeFcmDjRx
6PBh72YoG9CEUazjBM9gDJ/nqUAOOcIEII7f379RtbKm94sMtwnvCmsfIZW0VRL+uSkOzL17oOFS
2iiIBP8VPAL+BZOJDC+RGL2AmZND4XMfHWm5C5MBry4KbpjEZ+6HVo8iXvjF5spydAAgDq2g/3FM
US30NVV3N7qkWEUkFqYrupPbq2tcNVBPba/zfYnXYXZ7pYChaTiFLtNb/4ULNZbpTgHFZijFcI1g
95iidtrOOgnS6td3WNuX1tzHyrNvRglDPYiEpEa31tDcMunDH7KD+UBZmNZmiijrEkHSRFPxi90g
1ZFL44QiJum/1ssNhY7VqmeEmf+SvTiYNAQzdMRXwbom1txm5e1Dv4hbZRaYom8GjM1dkC4mhpmt
cAk8VJXUo9WLCsfU0jUCvnlPvdQ+qVmppqRcSm1U75HaYIX30UPG2RR5oM8yUjv37JXVBcGB1exn
barxl2QyeU3SWjmn1kXFHLfiCeC8rH7UBx0xk3i+iJ6OvOiwaHkl7vUbtCYHECNn2CpRyYILp8ot
qN01u+1DBQmXvOhGBHa/9PODpTj5gopBqxWgOAnGiOtGMJJpCUBD2nz3utyjqx+IDHS3BAV88yLX
+99qSR0ZcTloEzeAbk9sr7QGBo44ZImj/WmvK8Yk4JBorqMMrCj9wwG705wbbqJeeOBxWDkW58Z6
Hph+UQTivKN5DpXOKSl5nNYLxq65NgVtrNibNIveKCK7aoXOAcZOEZWfuPOesHzuKEdXEVkIyyls
lnI/FsMUM4nYCyvpK3kxAa8bR2Q7j7HeFSYYmlI8jWGBoscVOvkn8eYOwOkWct8VOjYr+eTJE0X/
ZViwjZ7MiIqat3iOsVm5ezX3XKlhFIJzl5iTAI4wP1ez3a/TKpvgF/y7DisD/+lh1oW2UsPo58Xz
DKxDiynj0orLEq6GYwTIpYT4HYR82iJWZolB7guFVQTW3ic2rnAz5RmvnVWRJddJYUG3YXxSgVG0
FNvr5MPfQYzf1RXyYpS55BlOePl5/ivlqQqvbiLebNqztzjT+dEMZvwl3xNdDyaUYYLpYBkpUvEW
NcEFtaZCjYSvNZukadr6TmDGF0orgqPVQa7NKH0OLx9NfAUXuDEhHU2f/pbMzockOzeH+yUDk2Gp
BA0bTp81milj51J5dqMZqzEPqiwm2vg3IqjlOe5roMpaWrEbqlEZ4yrub9gx8pqbXKIA1diRiLfW
xzwlXyfUKy+xd6muOtFmdtfI+Ew0DaoOzRCGdCX2IaWIuX5ECRSPvIjgAvunwE9rsBeBbSAVN3A/
x1cNSRr+x3X4+NH+r54dH7m3+d5ZqRVBz4xGQuH6UEzEadTQqI/xptpSVRnNSjP4ZxHROKmrO73P
6k9aYyrZgkzAB+XTutIdsg1CCW+8E55Fv9U0zeVPbapCRSOw9D3YFke+QZyJeSgxfH5+TawEmXpk
h8U3Ut9KyRmBdqasEdK30no1vlaH7XKHB5zuVJ/riPjaw4ULuGF07wGyCVZ2FgitPtCHY9hIwzQ4
B/MwOQJYqpPyrKjpb274dbASW+wAuwl+z5EWHEInSwbCnM+hdiAtlF0xso3PVZQa90N+ML+6HEJf
l9lxMFeraJjGIhdSltzxV2/PYJY7+ulPOvB3l4h924Zqb7LaSOa0SO9/AHu3xG7ib1Tf9wFtT7am
cY953I9eMVxAYvYXao68r/Kxcr8kjHpcASHtX5o85JbqwLEzJKsn3R7nozs0mGN5nctIfBvBKuhi
/ukASsZk9ce15oV7bWmVzJMVe4AQN5rd8cWyXM7wCaJEOwktjil7YK9wr4NP6LndJj4wTZF6jkDw
mSZ51tmIDAJ9Pd+51XUpD8IUtum8oBPowgqlJQD+2Q55PSh6puD94Ojnuy/lYovnP+ywLUv0E/PW
5iPrTPVzeoexzt4CyxWidl5Pm8PhIhrwGUDPPvJ4gENnw9qJaOhNKvrmxWBWnomO/THrUzsi/n1q
09hOMKsPHzXI+zW9aaEtlz2v4ARTe6B8NsNqp6VOapHUCmen0Fn9upjJ4jSWGgXwX30I3aNazXQI
m+tED3aNu7BYbeLTN6HOpix2UqsZFKSp7GzMYwnzsFLGTKQ0Gns9rFbBOGEHNSC26iCcOwYlXNWV
YPT6PVBusUl1hh7CXXyWqaDNA0KJMd3IIXUhXsc59+tjPXXV8yMxoR28+PP3xmcdsaNEkySNWKPF
ibfj+6A97FlqC8r/toLyyICB0wVfPxq4QdDMf3ZRZyIF9fbD/O5cS/ILIBD38ce2FzoCn/Eri0Vs
JRIwrlA3uvlsM1JNstWFXYIGOC+WICoENmsu6QUh8Cy2WF6dtNHMttAKRKFRgJerlftNqhj7E1U+
x0vlorA/yFRpd6hORGhRCsic49MyLduL0SACjzrB7y6/MKVRT9Q4r50tYZrcC4xKC8HfeB4OlSkp
8qK3re2WfS6DvWvQrbr6qaZKHWUZ3Icq1ihMNiaI3t2DEeuC0HrAQLYIfgv3UdPr9ViE9pb4kyOM
SpKAcl9aNT6gs3+Mzel7up+DfCJWoazdL8AYS1h37U4IqH0RYh0VryzEVIX7HXU7dMejcbDuwCOw
ekClNQYZ0DnFHSBjNm2Z8h62vin5IagyQRBl00ZlZpHpBY95ywYIpuw6qNqCJKEzGCHIAZAshKcr
IzT9aLdaw3G6C1C7zDeS53pTAm5r1NPhQMfPch8PJvJopM3TkqLm3GXv7irjS2W/F5CotiQN2Jzu
9fM6aPvZGauN/5p6PhbbZl6jzR4PrdRIdhGZMENo30xkzC4EFCZ/FkPknoJO0Ujo/bh9LV7srBei
hKdWWgmnWuQmFu2t9JVU9arqw95tI7qliD18VcGB504j3+9M2jI4wQ68w6copnZVTbGdWvsKjrFJ
LB/PRj7r5/LGbh8wwxp0HI08E+OZW5+NorIXsTpMSe8Kx9wBwcUVYnpsqAIbgzxRCk2Izfg9E2qP
7j5A/InZBTHJQP5IJ47jeGCuQhss3CJO7jkU/JCc2isGGaLVmT3Tdu0xVcEFKXF3SJZhMVG+gYei
c/hPICh0ZBVRo1u8NknW6U6/PqeU3XBXedf7uVI4sUIcM2sycFeUkp8rgs+2HCa0fI1Q1K5NUGbv
QrUNCmbPP+G1uqwbhKcYrKxUyTqu3zuo24PTSO/zb+mSUFUkXqMoD6qF0cVi6DDBKJ2xZoaVfDTX
cx6fFVJ9vIxI/5f3TofHul5Oi9tOiZHWqMWzVGbMUKhUr8MuLhBifRPpheZSTnmOJ7Kb025ULdY/
cv+Bd9+VPv5toCYlX02LK1/PJfmd/ZZSjtAsV7QWBqUhTISpfFiOSxUuxa6cJlhuL5kD/QdmB6kz
UCBVLoX6tVzIEwt10hhSWUu49C3KJg2SGhmZ3jTl4vGA7QsfC8oQ+TZxrahbAfAt42SEA4wVftFu
yNGsGoi6bH/grcMwHia/QWzMQsPBkEebCwCFEf9xLCpvEhymRIhOxTljn6gq+ZHJdmr6arr1rqOt
/1t9MAMUbnkvWs71jjLpjyfrgDRJve9QtgWvpY6IhyxogZrQkdefnDE6qhR0nraCBHRk6FrOIeSp
y6nuURMTnBTXIiQVPRdc4t4vcRBA+2fOySx9/waKskV+8A7zwZTN1EsRhVmPeUZMbap1ZlSGYjTw
gwFXQx0d/UCwYqjQ9S3FmlCvU1tHhiNAveAWLAetq+BRGWUUzHDTAnMuQaIw5TltZfV15jcNT/91
fKbJa9dm2xeuMAylhJf4HV+zgIynaqMACrRAW/BOOeb0/AeIylgiIGqsqNqBOOZhuOIPvr3vXH23
G22yPxqnMxGmdX99YcPrc6RFXbFRDGR8f5/1y2UFgP9mV+Ik8URq3HoeUBFrP5sG2pKtjgfgJ8th
Ypifos7AMuMI9pGN7KM97Un72C5AM9Bsl8s9z2tTREeC9YtbvS37R0bgdSud0BUox9/kF6Az0l3D
vPbS2aS3naPowF9sneBAeqQUqd2/4F+Aj0d3CVG49rZfwSfd2PM05VX6UggmWjXOHgA8n+IEZyIr
qh9dQtslVs+NUT2PGSECBNuWRcOxmo3bh2jh74ch3WkBbaf3ub7pvMI7EfOa0NoZbK7QnWtRKIHa
C9SILTiBOEFJVkQLSOOlYYeqz5SBgLIk1AkZp26zR/Rbl/IyXUldkyMmo8ls3aPTQlDqlupohggg
jgf3diuBf4IooimPuK8KlgBYu0cnH3jIT6DyvAjXgwj9qKNPcyluChxhBTq43ZzPuDmEpEvHSOG3
2UuNpsNdxIfL6iwQOM/iogkPBJp49vN6Q9htdIaOvL4o+AqQVRTUvShbJGxE2W8ACFBphXuBXvMS
xVy/VhlZjIgyspckWtnI3lUB0917c5gNv5z/jMa+nzfIkCitKMGtoawL9hl/QB0NCISjnYYAqJ2i
RZz6a5BmHTxkpdfnhDhZqsHNb4h53sn9wR1Nb/2C3jaoSPOaQlKO96Kp0rLvvj5yuMtFGGYpxPsn
/iNcYwcHAsLg/HLYQ6PNHGhgtgf51w2VVtdVYAtYIzivB3WFPOilr3XUqmVdcaekNN62D9WoXWI8
a9IMZ14Cj6AJnakBLJ/rnv2K4xaV9k2/CaQ+6vardwhvNlHJ2sEkd72irj1WIr9t+Hkay6gspv3m
tiIhcp4187m0fSTU4zmsqrIL6Pdl1me2K9BT95hqy97qJgyuCB0dIVEWTumkdhcltOmEdWIwdpFR
tDPyXooeal0B679iDTuCDAz5xdXynk1YXheEVTFwZfh6hV8n2Wp91OBI4rVezPMwKaKckGPwrEhi
f47oK5dkfKcuKvE89eGAWlA0j6VMntFYXSbyYTSirSXyUW0CgbtU866d4k3EPn90VMuNUr4gE8TJ
wP4y54+/fxTHioG/1oPgULZEHllLV4kVM2FyANkuRkPqtztPWe6JJhIFogBlANlCBnqD+kaAmi/w
gwxxIm8YLeXZfGpwAg+5YmiGO42B5EE2oeMQDdeAdcItJzXtDrEF9U+IUqxkMFY+OJmdWPuaUYUk
waK/mQ1by7i1Opy3Q+wz4oZIo2S4/8fexLblHlzZXQ4kD5oTr3Cx/H+qxqcbnn4LRqC5zhBOFTr8
nzztI0sDot6orR2ebiBjAXyEEf3JsUF+mQTWuRmJPn3uLRiZgs81yPrKeYot9n4vrS7A9vhztdEJ
uRh1WkNLYqgXEtYR94icdlxpzVITB7BwaDKSl/0A/QpGYXYNk31iRwAYhPNZNj8RqosBEXim+wUH
U15mY1z9Kim6AULic6RvkDjUAr3Swm8WPmhh5EgHVBWw1nIH/MbNiLEzFynJo6YWmaFb2wpUKWpi
FyvPHg1soiQR8tYSBdTfUlbK8REPvoQkQ3iOUyBT5DeHJ8aXNAfs4tdhy3i+q9EIjpyob3SIVDr6
oIcxgy6SmPNQi1PMYyTaopYbTjpmr/m1ikUWcocgtYopvnti+NLHIRNoTR02Q59FNxDMw16NVoI4
ScBrikY6yZAWOAuNIrBtLU4sVtdkWN/cCNddcXxoZ7EtEMjDXB5VVbAEWRaztNa5o1+Vd1yE0Bpb
+flHELnVoWiiNst4tIBdebRwZ52HQIxONlCGtShQuvKfmI8hh3UOQ3CWVkqRAMZA9Ka5f4hEJsqb
KFzqFdfjTYgF7G0u80LO8KCKDDIhbGzIJKedXIbfn0KQrdhashNNgh05UE1E9TbNJKSBRkYv4Yk8
1JCGdBU4G79Psyo0aq8x7NmNHdh9/Zjn7M7jAY4BxudVavmexhP/BHCNoQK0hXsKYjPVs2kqbJ+I
3gwi4KirovLuOIumSSiNlmz49JNjCAYR274Db2he3nWIQkXShhKehKLjQpJ36N+ItaFg1CpDrf5X
+fvEDnkt+vmDqJyRGCmZS7V51wI1PpyoF6w5CF+0RkFyfcmaTmuw7oTEvFfSRR6qPvNT9vkIjHuC
yRx0LqTUtuFty2tCyua8pQAaqqesAmxYBr0DXNU0yvr8u8ryTxWWxGVQoJKenYcQh5GpcDGkUsPF
gGSNdvKSRhvu1S0R22PMyghVfFRH0Mhj4eQXVpxMdc5leeIAQF0fqXB3sjX5b17n28xVkTc/+N8B
rX2Wcd5wJ/jpGw4n9XazCavZKgUwXsAs8/Hcv1IY/VYIUH5GbZ1cRJC+OQ/5cln8I0rD+FPfma8C
Tpdg+uUJ6lOPUqER7yIOCKS0FwtlXGr9wpK/3olLT5OQ7fJlpZhrRs/XAW3jBfpalmSz9cKbypUT
tndVbq2QeYlTCtgj1FlYUbpuCuFwqcQ9Vn3g3aR5LEtVoezLoYQAQSyhOQnHuAiiQWLlnK4zZSQ1
LzLtSf5qXzhMzX4LqdpwpayBqtmEUJdIvX/9cnYNnfmao8fBDHF/bcP1M2T3wtbmrDWaR1fG3/yw
9eZOFYZwlb19j6h5PrGTvAJ+xe0Nn3Y5mcQ+xfnYXYM0iP8CuJ4qatgRWikcJaJ7qIXY1j++ZmYv
MVcnfiuS+GxuUk7qYbuYgUGCWygU+kru0m/AQ17Iqe36JR6H7lwWlNS8tGZAzbj2zzmWWMCK7wpS
wGC0P2ncZN3c41mSs5Ndj/yYFkUBIyPE5Vt5fuOlgFfkDu9YrKP10GNJw+7x7W6oWXfjkkf0LI5j
0t5p8lUifP2eg5xVQXkkB0N50N7lBZKMM4hiZmZPEE8zuEPknluGBaj2l5HkaGO5LYG0srXVTfzx
DVjWafJpOij1VI6vkH6Vsrdimj0Dul/f7nPmF5K/nUxQUd9WpcIswXTd5wBwTXMln5aXA3Xf88KF
67ucU/lGZ4r18VA09CpBepoxs2gbLZftyQc7ZP/004qCOMOZEzW8+S5rVtYdJhkGwIfHtiqJC0VM
uwOC28vbKAZr2/aWzA6Do+gpX9z2T5h+BRw35PjDtGOL35bdrVixkQjWT1V+TnOgXdIGm7LIk34N
WkHCF+1MlSBS0jK/vgRTyzkzrcHPCVQl43ZVVu9UHSVZUGl4cuq/xXNhFlpFskPLTdJWQYTE/NUs
ZL3FpZAFxOby9pAe4pQ3FS8/JDikhfbQdOmXXWSTbTDvf1CGzXxMYRpKvRE48LHHPay62dqN2InG
43OrdjHgc6R/bYE+hj5SKOC+X1ZXlJafqNIB1sjT3qyC69MCid7a5GgvuLAdgoS6ejB6wb4Jl0R6
mAnbJFhplH5Z/ulfGHFVhidd7BoBxWgchphEh5/RnWQlPYGHOEyEfy8JwkUKBLgroKc/39vxY80C
YMGMtjCwsnHEAIDUgyL2t9ogcbovljFAj8z7O7pNF5lOyYtmYP08nFFxdJDUhMeOBlqt3MkqjPbw
ERtlHUf3y5x+7gwxMr/NzARRBUkFe7yy1dUhm+QCoO0UWOPwaFx/tHWvdNqqWN28z4dxdPDgZ31Z
O/ssz4FWzzbkRuXBMxH5icag/SC17feNeMuRTDoJtrY4mRPgzoSFET/8Gb9dW3FAM2oiHzC1dloR
TEXljmcvV3DKlNPQhkjOXevgksN1SOnt021K1MU5Yzc6mlxGwPXgrsycUT3CEkg5+zAJY+b6Fnxs
EmaAreVyzpG3Axsg9Vt4CqjBaBV+pE9gq/2UqdbGBjvJZns8OR2bDdf5drwIuzW8FHk6PkTRbXJW
LcDYLXhIMvMRw7bas6mzyonLZEUNm7XXYy0rg84aJvegykF3LzV3I/Kwf9FVBPMhJbOlfPhi00ZQ
16FMzjQspGWOkcStNtpZvdhfex/eSmEhKzoWtGPWZt+jOJ7bWCYuaE/9d1tJK8PKJrG5AS+sLZq8
byvc3pfH5ra7bC0XCwihbLWK3meNx0ouuU1FX4AVV8j+6FtOv4/yEJTMQlneV+SpCS8LcSkpEQy0
aGrVPdL3bUscmLpjEKF8eLZpdV0pW3d1MlHNadd11N45FwoCjCRh1WS/Xp4axqlRP6H/sR/gzHzE
mSk79kXNRjmYwprvIYCP5PntxliZFEOKa0tIET9eTdcG1T6uIbNGQvDR16vg79gWHqAPP23JDSJw
I0c3YFpr7/z3IyU0Uegj/nhzcFYjnixZFTcGn9Onqp9q6x0uorY0dSW4SpF0v0Vr1MbekIqa0qM8
hU2CTWrHLodqiscad0BwJdZbYDCccV3x8GZRWyA/ZZlkZBFoyZMb+8mSRSjrf2/cf4cT+4oxkliN
gnWJWc8BJ9os5vqCIzCFa/eQ2rzuylnUmLqKGL2u3+8nKlnyeWukjDRjsWefjtyzBi8HhtHW+xbz
vlS26d2b0RWwAdTG3Kwptr1kc7bhKKZvFi1xbPhfTZpZULiMsyWOrOog14LLK0BMQWukDczYvASg
JBGJFb7yL2IXlRCp9r7m4x8MJ0Ti39AIg9z99/8VyMNYH8+XEtYaCgayOsOADqPsOA9R1K4bb7N/
CaOdtCjM4iRO6UUpUBxyfVjb+M23vQwuCt216D/bWKfMDvxnvRAcGhiQP/iIz8tNXGEYbhaK5pjE
QedUlpVqDQJlN0WFWdhmCByjPW4e4nPRDmEA16m0cQtdNHffkTc5UUetUCuOY0FWf4uI73P8x5Q8
hLkEZXA+gJbTQM8swm0VsQkDSJk6KhIH8cu1mMgCmJLWd9CcgvzLRrF0A8GH2cA+No7eKY/e0nir
l2OCe0SGjWrQa8o+1X+OzooZGQFZpyze14lKuB6n0yD4nDZTM2+K6vBAT97GhRSX3dGmlj9VI/5y
K5DMkUrmqH+Kh+JwicSuXPIn2NfJolgKlDc8jpoQIwSKntKFllhW76dSrIhJZxq4s9X4ptM379/5
zKVzYFo5Rg9O5Q7baB46IzNFyto++5sgErTycshk3Pyc42fH1dnnGsgODCRi9YqxKDDbGWyEw0m5
i+r66um3449L/0cjuzzluX9qe+Gqt2Zh8fkMEehjZRmGxiz3L2Fbi1u2kGC2EDWYEqwqSZQYlSBw
TUwYU7EVP5fbI4EBYK7LdWS+7Cy52Du827NVZ3lSMzcgyXqIbajx17Nq0R51W9vM8S12Sv2IiyoD
2l/8DqyMedtXByk5P81CjBRPx/8LK4VbB44R79m4OE2I+U+Gt8PDiiHOHge1XiwdhiwkyBhLAjl3
KzztnaLZyqk6dKymlupAehXQ+pEcisO/FAAspVjRKcoYnC8pGfuFJ8Vrt0K99GUAHpLqQ2iSD3nQ
FzSyd8k3rVcGztJ2TP1nFnW+/4kwD5cMKVHirc9wQ/wGDCch1MO+WwiXouQDBpIALlAkOLXLS6u/
0IavucPuXXG9EWTWKFrptYkhfmI9lAJ2xgXkCh8t+o35c44hAQ+0/t+ve/69IBRDTUgBDm0IMrAy
1khgVNF3JM+5hJYnkCbfhuv3RJN1/+gYTYMj7qTGEBnqpUFNeBDOh9g5Z5ymPyz2GW5iGsUvJj33
T1LmqQSZ1wQF1+rgP+iQd8h88k39/IyvErh/rjYcDAeSRxagWcSH2hoKvIDHexKY2HM+Fyqyc9o9
BIvSxrnV/L93IAwZ1cisdQKasmnEVQF1RezhF2REcE8dXN/KhUHodxWsjhNn18vNFt1m31VBvKHm
WvVBQiUk8QWnpJwtpX3cGI0JvUPNG+t7S7sO7zVFc80aj5xbMYT9NMXGxmy+MwTkYEYHKnKhVTKm
aeL9ZE/SOyLTCMYEld02DvrmzaCp/RM1QxTqB0/bOCnu7bnd0iPYQHYvtKlD3OKJdnDRAbFAGeVE
d6iQbL7o5ox9/1KJTZst+OkAb9PiVYccpOH74s7DHURqXitrhGcWFAYjpOVx4jhrRhYkCZ8UkViF
cD9TPlz9l2YGk1BExIeCWWyCSXAHL6zxVtDB/nw42C+tS/PkUd5yJm/5uvHZt/C62YfwLbfN3s0n
fA1mYaDC3+ZKrWMQOBSDU/V4K56ERmDJXx/Th/W9wqmKGQZhPsgXxQLi9oyPbYA0PdS40JXOQ5qz
uDzIJQ/FnbfSI+DFTOmwyZJwzivhkNrHKDF2ovuL+hnJ7evgUhm8zPtrrtsM6vbdsGop3y/HdcTp
avns5RpYyUz0gJ9ZxrAl+5rD/xqKFIKSRqD7KS9S15CyPJ+hrkFR7COJD/RJ8EZkwJNIcxcACDks
2a8Uo7+af9pg9a1c9dkQIJqKA+8keiUQ1EQLkKKCTUVYxCeLLMSG+ZQcDY7UZcbbJz9W9NRNtvqU
RJWgd/omBQiFHXnRdu5RtTU6rUEq55cusv9zb+5xHUtDU0mBIv0D8+PI4tL+4KoXHDk3x9sSQKtj
10uaHDs3hp65kEmYxE/vZ0QPpdOU619B8b51lQXiX1LtPl15F09edS344Tn28/TBCcZOhzAIh8BG
6sQOCr9dK42Kc8Cx8HrYUw107+hTQW6fhUhI6N2eUAw5T+83Tr7pj+AhZsLjNKJbmrFbyfuHOshd
lY0gvLHLePtmQL2YfeC9zBK0wYFGkdrL5j8uv5SQTYLuwPfdvj2Y+XOkx9Smb6z5M4lIc+SGTpAD
/cHaA0txJKEyqwm/MRcUodTYtRYtnOHOrVK3joaCNzV3435cOmX+r1mGZKg5pEo5hERLIhLRso1z
FT2e6o5kd5vTlcgkf/5ZYpCTlRM3L5GDOROoG/7AIQUudgAwG85gf7D1UzN8OzTRtJs7Te7c4Jhv
PROhxzyDRDr0SrNtRHkeFN4H/KCmr1Rggd4o7I28RUMWUJcc9dS3V5lmp4xRjhsiH4sMrHAMrT0Y
jWb1eJHWpcMl07vY5arQR+Nd6h8gViGHsjXrM6aQxXNMpKeNawbRkyfKtrpRkMSyvvfsFwu2OPfq
KspgazP2L9OVPlfhkfyYQI46hdsvy8zDjlOAtAw3pmRFdaiW1Dn+75SWViEDpAihK53WHfEdpYDA
IhkVEFEdBJ9s7SY6s7e9iHcNyjQUQ39vBfYYwEpO/JXLaC1fF2VvVNLS940COLX/nJT9h7QalJY8
Y0gG9v3yUPjgYaugihCqYRQsYFSCgZ+MlNzdaD7NdBRInJuPl8q9vdI2EHchYacfqpp8XhWRyQ40
sbEKBXdkL7igESKXY/AXazpLfLFXvXPacUOONj2Su/O8+LSlz0xlcAD1lXXHOK4kAlrtNz3wkaLJ
wgbHWAjyvnemKS1AD5cX7KFlIS0E5yu6cwj8A9tEDuuiQO4Gf8ksU+kTYXhWkbeHW3ZylecaCkrm
MHUHCDC5nIK/+GSlmbF6uRIZ38G7CEEUgUelNaOWlDH3+7uQxXSpxiBe3V3Sc4KU9SKukIQ0pdXc
jBr/hzDU48FXit5+x1slZ3KqDWh+TYC4Y24PP3u4xSKw0nj0Eypde+m1t+DW6Ambp7/lW8WWLdx3
PHHpgS/fAJvjUY/pBsprf6YeDySqv9bLeIP8WHlahRU+Jo55jjJi3PDQyy55OAW+77ZZfHcboWiP
5uaIeSjx5vT8rFkexrzy/4VG18ucSWQ16iPgYPeanG+2GM4J+ptMSfQXO2phzZZbXwSInQDk6WCp
7lUst/cvmMRg4bzgrbhrQI68Ir1niWqKc6f2ZzSi5frGcbAmPuKu/NfSoIi4cKB4XurvIeaMkwgI
3t9MczhSpRWFu8R665wDgE7tzm5BwUdUCSpd1OZBMAywL3aDBw7meZSS9NYwdmOTmA2N5VtgA12c
IhMqhNX9kpDnKDUrmNNmzNznJ1upk9lV1bL0BphRcoUA2hMan/9cCJdQjgz++gkzCRCJmre3tIlB
ovCHrIJAbea+vmbAdn43mbMrpn8f6XJGuXI8LwR9Kp4CFNny5UKDD0NYZm/Ax1kBdv2uPoo/ziCK
aDiPI06fx9zRaMPeYL+TgJsbyV87YarVd4Rz2fcWl5KrF5qdihYXDPWaAsMDN400CKv7kISRsHrG
RHTluj1LU0dzm4f2gf4rk1obC8t2wgwQndTdREyMUYp0huCx0WM5RRXu8Lv9RBu8NMY3zXnp9QFO
ngtbrajYwjMu5uSuxAdXxhNhv6yb3bWBiQCAxLhV4gZDbDS+l3X8WD+ECS5wgCRNVQtrFGGI7IF1
hN1w1WkwwpLeD8DR+nmUDy4DX8NIBM4jDxfsAAdahug9cZBgI9OO1SezzakyNIYhwZMJwIqzG1nE
xb76MzvR5s9935dWlRM9IPgzl/6of15IDwavp0VXKmQahBL80VbmpPyul3E8drGkUeYBhohJx6sC
DFp/hCn5Qu8CjUyPTJIWf5Hf8qBLeI2YjCECz5FSewkRSaNPdTa7bTeW0A9JN7GfvJn8YEPM/Ypi
YgyDOSq7bBousLl89UkF8teTrm8X2mP2JpDKqRBPXoUuX9g3/GaayCGxlQ+FGfxXQWONtXQtqNv4
b3VkN1uh2Lb3E+fzbIiiCyBSf2lsbvm0s4u2LrHjhA94dAwby6RSJ0YiEgDPz18BYH6OXeSCvL/W
CgdSl5pB3QCJWhP3PLZtoTJ/D6HYKTcCxBmLjZjfNqvhB3lqa2+QhhrnforyyY/35Ki1nLfGwz/p
t3Zth+dZyJb98j6KnpZ/lPGmG2+wBRML3OrUuQsCH8OJg/LlxzeIXEMxAR5NWpuOSfklwgQwlK1R
cW1AJd3bSHfR91/Ccd040/Eq2jk4VGcvfm99iq9UhbjoCAGd8drDybrTmV1B0j/iPMmfFurgig3V
Xs1yirI60WYbGq1Ye+rugg8CHe7eQ4RWqgvaX+badp8FSKXOVAn8c91iN0DAMF+H9RZqH5iHpmGn
4bL2T3z0I7VWCkoml34XIb+cZj2QPvFyJ+n2KeG4cPkKoezM5z/pR2VG+DEpZrSYs4MvnP63VcYW
uziYW4QIe5tk5iDXbGw+FfcOSF+RYjH0ayV5NEIjggzlmR/7Y3MJpCfHgfQyPxEho0RAK6fFmfR+
ejE7JwFHifocI28u5iYSbXqdBmpAOp/L6Nmd1ED1jKdjAuuWgFxpa6gJwesnnKiBd7zK+f2EOGu/
DY0E5Qdbh5o2Of6Aa+3v2TPXzbzTZKIvuQsGqUAXxqt9dHwWSOUoQ35qAp7HVhmk+mNDU9LUWHzR
GoQNPHRmWImDzClULYLIS7BhmJAwHmkdo014r4ymzDuwSbPS7yGl9xl89hoxxejw5JHOBIQYCZRA
unzR6eY1K4+P9HBeOtiFyVSi7olYOyOyzP0/X7VbNkqnvLKqsyC0sFz4Jab2S9B2cicf/1WH3NOA
MB4N+3JlPBe+XyPop/Fl94VS3IR3L5c3Rzr4ogMw81oHeELChVePmaMdrSyKcOXwGtCh4OtQDSHu
ltnmJ7RKBQQt0eXdgsp9M3c/cA/6CMB7sxkyxLcojyNaNDxFJC8Lzpyzb4AmLDbsgpzBLZGCNM/9
T9zJIbM0fHPGDOcavz+q9TCTUU7ChFKMDMt1okD1y+Hk7afmL6ziL0PKqjtj6nMkJ8XSZWmgZST0
X5U4LLnDJbLKmIes9PjdhnQL7pQFCY/rmdhiNBonCSnypRp3QKm4+Btm+7XpWZoROJv0H7o1dXCt
mFkzmShzc0PPyIMBN8ijpIHAQtgxqppUI96Z5qCrlm1PSOZcfDqJLHV6CRkj5EcZxpEXSx8QU9R2
uZ+oXI+qD3LubZkLKykuyeovaXdvfb+cleBCI+QKeCKwAVzRahr8fJE3lg9tEQDVU2g2EiaFas+J
JB+kXLQ+CEScU+KD+gmzvzS+VzRv3A7VhCDrcWTd99/RylShwICY01iDGmwI2Mk2IKD8lAideiG2
qnUMJ3OjZjutFDDEO7FQjdAahZ4hFlBAhB5SI5+nHGA7xh8cpmlTsQiIr7cfZZzq/1X7rPwsfsl3
g90w4w0+6SE2Bjat82lIMBmsNA423JnVSCSCobKwS1CAZnMh03/QV0GcqklZnlMsb+EVvvLfSTYv
rUuu36c2B1noTp7+jhBOWedytcOf6I9VGG4P4yxbh3D48SO7IpPhQf9uLwDNgdZ6t0vpZnvxQNOG
njxxze381rhc7vfQhc5BUA2rA3BwacotYxsmsj1646TOAtxRiBbbk8sGC8R3aLE1+gwVWL8SjSHh
1w0ZtH4iJf9Div801yfF/9yA63Fogtpvzu2lSPDKT203BrvBbHjnLH1MIsOqMxF0hlMT0BderLNL
7E19DAwvJC7CVyo3EU97hJIGHKT9jySs91cLRw3dhFCd7Z6p+H0GUTUwgcIUebhtinDtkJ9CRdbH
V0orm2nNjxkIXtIqKxc4Qt+pmnyk55AK74FKrldWzFxLnMdh4as7FelWYrr3lg7HlBRiS3cVVGlM
yI/371l1Ozdb978lvTPOMPNbG/py1mH8LExOG0qUx+7Qj4S+2RvB5LOSbfBl63W/UdrplcK1kwRQ
Jdfg5UCF/Ud9iMqRPDdfDo2lSsuNH9TbYjLyY5+M/yYqO5kdRseJU0yHDEXcYYuCz5a4yk/ufvd4
4UDZMFy08b0sUSdi/X4t7kcTnpRmm8S9hMedw14SAN/vmrUI7WcVAMHqgzprBcNatxdmD+OreO0a
afBh+CVQMISs2L0MNhqHfqBzeFgZukGAG939Gv2m2tdQKJDHX6iA+XecbZecxmBsnO/DUnhOO1CT
r10jvGTMvQJJw7WaeXwqdR2VmjW4QPf116TU6mITG2dcwNEg1pfOm2nQye4Hr/8vMqkmWc6ps1Gy
SoDwK/qr+W8vV4qMX2dNanIaNxI+Jq8sX4jI0k8L6Qlw58j4aDNKft3SD1otA22TR3axFjdQ8ZLh
YUB/Ga4YQHcQ2Bs/U2K+wO6oEkd/YYtk+543ql9spkhCZVLc87Ye+PqyAGIae3M/KmbdJp320gSJ
4pvkuiOXifJCsIa4tdhXOv6SlVJ64GlfPf4bPS63FM8LVOfyDP4yP8yoW/uffWy70UEMbc0zKH3l
GdEGzeuWf4qmTShDDkPa/Lnf/H+HUK96LSlCyvRMY72JeZv3W4VD0xL3YVKFMlUqKbOWswsr6uwn
fobJqun8uZ739e6e0z1aI1jgIb447NulbnRSGumk2hU0Q/qSzSUVwPkCOzUFEP42cAvcZ2vMd20F
FptCS5CRtMQjkWrKKSjFhlgQqmBjbXTsy67gqyiZh2fckHrAoOIjXO2ZzF4z2GhlDS+3pnBBha9K
DZtKc2dXBiyq65rP3qIinfZUnrC6uAbOltyvhWg/UoXXBmhvi5023vnbQMV0skriOJltWM26A6Nw
0b8fxE0O71NzQ+PFSexw7bBsLUS+KyeIGXN0ZYqQdCeQuUSJPNxac3TTw+wZmZa13l8jQQUOaXFJ
anObr+CuHkoEe0MdM44MbyTUC0ca/OmmSpQV5ErvVIyIuD3A7b90kFnOpjeJZ798deku2XBZi8Bg
4egrmbqaRvF8AfrwE2aSC/ncGLPE92ZZxg5U/4A3jBB21WTfayEG9bn1WPUDLEJ7UB2xqMEVx9/A
gZeX3YI8hRUqTkXvNRNIGSCs7d5iDCLfcdtPQAwlg0O1WGG2ztFeqUR3mf5Ef5RvYW0y9PilVqzB
KnaS7ruKUHAmx9fVF6+i/b8qtVjHHR3HqoXcqfPLe1TOoPYjngIGoFfxjwDAgydKr6h3JaMlr4Jt
uJ6A6mvdJX2RwTbu7ZQZ6e+Xj0AWzJRKiU1Gdoy1pCfXoTzlw8f4Mr3bFXgJvvIips6sViHmnd2e
6yDg1MbJV72aynJFKYk1nroNQmOP/SXP50hGTX3yc2atWaYyuO/DHIhKXyGWt6/ie0e/LE/PERXd
5hsoeJsqzeyRaJZU4nR4HnC20lSZvtT48Cb6WsnDwCA6yG+hiKUDVMXK4/vqoQ1q2vRI8uBUv4mc
SUW7pmvSbyYKPWjuYNTx43WRqmijlUq0f3eLrezrGTLqHSDQ/v+Xan9bSHdzL2Hx1mMisuvynE4D
BS/QtxzDBh9nMNkyXSpkcD2yZjH7mhxJlnqUX4u2tZKEn36z6z3uTuj957VE1a/txJq73cUR9cwT
DEPM57LlOdCbTwa/T50NMayIpICkmQzmDf6bq5lr47HFq3D/PwV8363VE1VPzc2gfPWIoihN5zBo
qXPuD6G+agdybKNGlJbOuK8MRIzVMBH+IEqzF4vnaMggv0isssegbPS/e0r1u9eddlfLL7+72sqx
zvQYwmrIqYDts3VU295YQwRZ568mTKzmljyH7FIhEwiyoeAWX2XrfmhqKnpyvUHIF/EIhFJD4BmA
0/WDsB4SIH8aMX+9xiGDB7lYY4oqZhlowz1e6alpKQ+7oDfMll8SXx1Ct+hVQ5LmQmaAn3CqgYbs
9dRrWhASMV1vjGbniSvpE2ZMm7dfyFlA+g3Pjahs8gIY1M8za/Np2gc8+qiW9cST5Jmr51nMZTT3
1LXswm1r0Hy19sgKWKMeaMPaADpQHKrtU5es4EdSzbS3bCTnL7EtLdRX1CjijKkHS9mnzmbAy1QI
C++zolKK+N8PtRHVeUMcxcV6opwhOBxbseG1s0pXddZu2pXdvfdZRArvR6KFOLE41QnfbL6ry8E0
S21DWybySSXWpg1xaUJOWqt7QCECUXB0JBAOhxnTUWZ0h+RaoKk5tT3u7gQyn7cCfIM4bDT7yd1e
Cvs2EP5mGRwnJE5KWDwKAMrhClOO0Hf9I65eGcrMWRoK+iOvyj1QMkYTLS+ZtDz6xh40RCSIxGRm
WB/ER1HdYdIZZiw/u8MpWk9Cn++BDxKtpFt5vDp8icUy+kgJm9WLRTy5PPLgLrVDeI34WkLMGeph
AI6dGkrV6x31E46cR1D6ClMsIRSNVQ3Bozsanf9ORyXHwr2aO62WsB8RsVWXgjE9vek3qG6lekLZ
0jevRWpzmSD2qoGnjnokB01GbZFbWihaGus57Zd738d56K+UnOk/E1aL9+LaGcMqz5Yx9D3KDo7v
5/CKa4v2m5e7WguyGbYOcCA9++Y+u2UZ1yVqOwIxRXb/Esp1bIfVqoAeWbhb1ZR/3EOKemGvDWIo
DnDGNy9D7QJgIH62nlED4VLFXa9fz4Skydrpqw4S3HPNM8lKswq+v1jbLideikg3k7Fm+7nDQr1d
3vFjPxM0F3py3yfr1tsF5IOJ7W1GDTLtkIPOq4AD12CHIcRpV/M3b8xmn2o5sU/OdLvOR3WzQfZZ
SP2xurwM6VJECOPTgLe/fd/MdgJoVA/whPmAxabjSlI+tHM6u0MuBIYYvK+QJoMuKndlcI5vPA4G
GlOixYkseqWyJ/QXjJcDYQclcM2sqgbuzqINsJmc0n2nxdANeqdWuKKmzdveP8ag66F4LeKjdWTS
VeSfhVq+GHYzuoiRRGyBnK+b9Tei7bcJsmmvJOEXEgDDeMmpodhn5/kIb3k95F/Mkrl1lCUbn0MS
pMJafGxHvVTM0yQhiyO6RRc+4gSXpXg232fXrKyvBmFvwbbfpQXVHLktTJ5yZBseeLsvaKspBHT0
SVxp2vu7TsNXHkAQrNqjFrL7ojigyOixYfcDXeB1jLjJq5C1pCM24NvmWobpPELY/Vaz5QLekY7R
vylfsr1on5TCSkUn9q1zoQ/8yntP9pKffJdMdF45iQbLsyZUKv4wqMPPRkTPOY28iw4p9VPjhgc+
B1BOhzEz+yp/qzb2VjoctUFqRCPISmJ3WWAEpv6YQgNZGrMo3z1sKXJHuY920/hoPW+6UC+FUWxP
io3KxOAol+LpQVg+ywCDrgaH5KUqp3xISF39Jr6/hKsjbRaZOtLmDma0MboLzAQ5BEHGDBmUea0X
jTXqx0FK1bi5O2+YAyfP9IeO+8E+HbyJuUgMdUEVyUMmvkOb9f5A4TBjKSyEp5fXPehtjyzVEbtb
qSiL2Mn8k3X1+jhzWu/mctWERx9XUocJ34oPIeOddmVbtj3/6E17+9acDA5DX2jv558Z9U7PbaOw
DibbCXo51uQ6g7RG9SCI4kMAFMd/FvazZBwqDvfCZBtpn3UEf8EV4gskjGmuEFC5NR8ISWjGuBw+
h3LVo2vYDep2XwSGlGbt2gaMyfjmyNU1lNLlCkCdRcvVa/dAzjJC6DpoA974CTbipFQyEecT6YWj
qvC054LkGtKlJ+P7Fx/XLO+XfhClcmuP3V5Shz3tpA7JT+uH2ftNPJV1VmWuowuyYSJSLIJNHdVa
0szW7Z696779o6qu6saYQ1B5nVEFc6WV4nZXEd0k0xs+9IRsxAfxhb1+f/Kjkm4cMDLzv8Rk0KfP
KYxtoshbuoWkaCX2lLs792RMV1IgzfEodXyMKPdDhuPI/mx5/f+ns2ywQvaU5MvKY7s+EgiBUmPx
TzvneqjKuTLPqGsXIQbvSX4kUEISeV/G6BCmlzV6F1kvib4XzPBwGzdj3F797Y5iD4eRzAOZinBl
Kb3maG6G+Kmyq0HVGhWeTaTfA8ExuILB0G4p5sbE6A4G0pgqIlsXz/i+GnH+Y60Be9tL2eaKn614
TVKugoymo8l4NbTLwq4P66d+VJm1OG07lgMzIDu2hrUBJ9h9KNTVaaITu+kDkTgCFbZVGt9cALIn
fmowE3TqdyoQkHz3Poz3+NoC6xBLPmuP7FbTvK6w0AAtxfswyF5AtuRtL7Qgv43+E7nw1o+x/8Bu
Co0BPVehKfaOF/pj8GOX7P8ZcJwbL0Cn3DSp7pwdy4O3eQ2PnayJjSDo96b2swzKAw9VkEHVEYSf
2OyrykQnHvYvS2/WMmpcwkOf1tZbt9qynT5CJk7jPe/s4Y/O2cNL7S3zEfNObSo65SoNT00YE4by
yGEcA6ghtZxVOuk058NmMK5MzN7t0MWmpir9Ggzf/EsUJnsJ7pIGYMiJRqlS66nlbTorFbMu/68i
GVGGhlDsO6CYOq76D1zLTxOksn8hQ0z58hirOLTFEhOq8XeTZ3kKE4jig23hdAO2j66rN4GjNjjG
XS7Uh1a+cUjrlEpJ0ksaAY+E8vwMEJQOHqIPW/vUFbwY+BF11/FnAaWaQ/dVbSqO1JHs/1fuZCz/
X1xDxvfDHbTZghbALNm33jmmJTxmobBaeQRFL0qSa1RKjzjPGl93iFbZbzO3CSKZXgkva4agCRRa
/bQost1Kd6IHFm5NM98TkY7M932z9edvRqU+6vac6IwADVrVni7Rac8f4NpncEnUx9DGlWQef6so
GIOzmeHnzNNOY8X+uhC87d24Z5rZtKwv0OfJ+L+AGOYS9rbudGa18Jyz1e4etQ1HJVXdZ9lW+zzt
h9lIZIyZolMqtOZRG2aEWRWX9tg5Tf6yLAcMAedEmeIv045dtoZbMx29ID5uHzjP2gIae2woPZY8
hcfknIheWxSRSrJLkGD+XEZlk2ni8GXWa2tgp/EQv8OwYKluZQx6KWLCA3iJHFn20PogNINScslz
hi04I3TAlyqKqEpkZVc7m5+HF0WIDe4VIm40a/S/q+mAZnWjcf841mfkhSF5A4kPdzlsp8YtEnqD
A76SP1EpNwdUtMATGndm0/ER4N8haHZ4XpdogMgir8/NX2HieShJact4tlORHHyecmPTlYNZ7DIL
mPXlzjUjT55CGkY8sWokL5n1el9kt90R9O3WISqBPrGTQbFxtlT4R6aOSaMsAjppmVNFueuiAHRJ
6v/Imrst9VTmZ9RA3sD7jc0LTReoh1ekwNd3IS0SbPCO4hxzls94uZvxXO/i5WBrukF/Zo0MTBo5
wQjlVzZjzuxvhfJ/z7SgMRbdUtmCGMPKGgWTxKsFbQKRtvfPNgCW+9ZQp9JkVrMicack6UvvX3rv
Hgy8DDPG8y0C/5rCJdEBEXP3eUwT2GwiGkevkbzRC3KhLvtNef1TAPboY/EegZQdfh+CdwhQna6P
M12oH3BKbQWOMIedhGhb8oeOQINypfzWvZwCl/S+VZWBwV7l6TLsY0p8wOslogqTSJNkX8vMmaBG
BJA3x20ulGbBDyP/E0JvyAkKvUc9bOcKmQxWgoNkeyfzlAed2FJvUgZqD7GwMd6XiHCW0DPSBFSf
cs8OpT/OUoDDNnfJ0ms+FG0TbT78x4lU6kJf6hkNoRizxyAbca2HcEp3D4ikDtLXXIIlnyPAQXVG
qly4raFgOGGuFygxFts+ThsRJvUNx0yVIIYuLvGAyJMoGXkDj617+XNvA4NKA9QD6YcvGLmSx1N8
pBiThO0cfhAymJcj7vN+4Il4S3qpCKDd+N3VWMh3171AA8LnnvxzA32oui1biM1kpc5TJPfZtyKr
CQjlLh0szZNLWYbWl1jFWMkFhy/VP/tJYOmZvEgQ5E0jhb6TulAERoVMwOO5q1pVlXUptqzW3EWp
j3uzh1YgBeAhrun+nwJZXivPsDqFf/floYqEXb3LJp8MjEgjRWK/4kZmIjVl8vqXOfXpaoGPSpiF
jiQ8m0x1mspbK1+CYmgV6YFXPuCKbXnE0f5p1pqWZ5gd7/HRRt2eiktUKc+xnktAQSf3kUD7CmjI
n7kDjVrdHs9yItnxGZlkwxUooCysDm4XPi1ihnncwVYdZGqgZkkJZ6b/35PLGI/fS1cNgpfLgzvi
H3S7z/8nMVte7M+9yS60dtA10Y1ysPTKH1Ckq2Jev7z++0jevbMTVuwOfVN4PZfPxjv8UsRUACBF
/EEfhPOj+radkIGNIwvfkkh25Y6swoM1w6stRJawP4O53hPoyFhLWhiER1r3Oc717p5y+SeoxuqV
WiCimqE57QV6LNaKvcEF10PgkUKbxKqm+7ONj7eGbi41DpCI2hJeLHWFrvaIKFUcLekEWEssZzN5
QmRkdVD7lhkO/nnG9AaOAG3Z/yH7m4fNxii+VioDrsilXclKlyg5yD3SL/sMg+JQSGivz4PcZozc
myahGHd62+pCi6OL54I0glkzDo/GkX9IdBXs2J/XcypiwV0a/Dgwcxkp7O4wiQ2LC27ocPCeO1X8
yRdWpK7VG5BFuZBlA8CVUvYLVypkvlimbdmPhlqpI+w8fXuaP/wv1X7c9ehow3GCFMZMKHkTwsoe
cOtljUXubko8QQyYTgOzKTXbNmngI0EQKB4I7V64pU/X7C9FbesEdHDBJjM2okDm5U1hEy1Y0Rgz
pn4Lhdecg8SPzLQ3FKCLvE2qKMdcKnMiqEcNteZTELZ1utyL7Kj1F2VbE9H7taWgYBVUABe8QQfQ
HseQu5XXnwZw4qhRjfcjP6afowd3o+Ek7KYi5iXauELBLQ/oaZGWg9cjvhZpfkf2cewRLja9h+lZ
OF16q4uE49RXpO7h1mUPJWVo4tcncCPDX4F+7Sz2/irQq2gLhPYGT0izUoHms5Xj36CBWBl1oFyz
XJeaze5RGPwR/tq/MJxeZ3KPnWGG6oXt6bahpX+miL+J98LQ+/QiD2bbdwhn4gpiqeBqVxGLt7Dj
+AcBG7SNlr2lYLP7k8pJKUZrhts5mJjhVbZ3Uu7N2vk4IVgjGsLQB2OjBuc/fwYI8znCRuwwZZNy
P9OjvXF3NEUkD4XOX2xJ8CzPpaA8+Sad6+IZl0tncSsr7r15YdENQWVnG7ox/NyJqQc2cWc5QoLB
+kEjfNsq0ICSmb1msfYrKOAfqOxPuwpkXs0XQwBIfZplDrCdDAAY5o3ANex/oBvLtLfUkPchxKVW
LYqGZFRSTXWrjjhf0QBoz0qT2/6F7+/sbCGWrO0UA9hTFUNGxkg/EztWLa2kOQm3iWh5X0JivO/A
UPyH35oY0HVjdemkmdXkrg85/3ZEElJIj+mbsQVT1a/mmyfOdWVxBfXyqfu9IG3KZ21WEUJDvBoy
8qc/wILCx6/RE4U/UtzWd2KI7CvkswMdsd+pDyGAI0qzTz1U9K2KtHq6PvHZgzd2MusrRRuoNtQ6
BfvpGQjujVDWk9zQ6mRpjE0DpJagZMLb4maASTnfZ9z9f44YRWJKsOOvlW+ucrAqc8iAAWwp4Ccn
79Yc82oNXfa6i22+p4tGW446Tn3iea/Xqik6R1m70p1RT7nBOONA20GPQavhT2UUsKA8GjrseBKg
dX7KekPsOV7oCkpzySHhdK+TrroMZo5RkgZLeYngobTpY0kGUEb1XGbLX2sEpXlwh1x9+yOXmTJT
C8Z/9dFMNn2bFrBxIVNffYvsb+aJ//56XdCIDb0z5/vUiyW2ZlZv5onwRRZFjYcpcaSN6pG+wWIC
9WkGtxR9JvYyrkkaR2O5WYLVJdB35aTWu4TYgX0OYe+jNIVqX2Jzbql5YHbjsUEszhnU1KrkzdeS
+TYHokH7IkgQ2EEbS3cBMPMfYLtlpF3ESXPv8HZ9XR6vt80mgkYIveeM/0wdZHkJUjMqXCKiF5J7
ULkJPA40+edqrEGpOF6K5O3xwmbknQbF/pqEW9NrEz6UhmxA6CNviCsaKO9JbSQD47Yvoo3hs9Mt
iyailfDsukmLjLdAGWH5MORjtjlpOGm0WZcY+P0GGKy6RyDuMFVs62hWS19kyJsmXmU9Zf3TR/p7
CmKabcHeWTB8kIFQIi+TQqjIcqqc7ySJoLak5o6QbhPtk2ES0ihlti4Rp9c76ZWDjSZUQbMN/+DP
RSkDsKT/w2tgD6s+Cu/6DsoVjiYnlnrZbHjGe+cBmrOWbyhqQDx9JrLJcEHh94ZcvBigta2jtQ2p
eoPQEB3EvS0hmTLS6zxO5TRHvYuRA0/e1WFALeL0YrhGwWSIsDzrGG5gp1/Isr73JkoN6DdzFuNs
s0PQ9UpqrWqnPDPGpIVsljYHl6sggDnc6MSHgkK+b+XmViPhZnqHHoCvaFWekfD3IDR8lnAElNw1
u2HFfd+FCH45dZZAQ8mVhQIG9MkpCyu6xARHIx+WpSsjwlT37Awm+JocRvwPRN6RPkWRGQjxDpLe
aZ7OG25Hnh/ro1jpZx8oIk5dAPMJ9bjfu1VHxQ4VO8eZgruR9b7EWHV6a4GTfOggEcFwXCBFOoix
JJWu8/HcHDxhCpL9aLdb6QP8TDE/QPFJeAM5fLCm0eHu8KhbHQJFOB6DMwM7fGoSiWG4eJMkHluw
3qkyQjQMnBsCZkuaBZ6I2DNkI++J8XlEfde2/VoObrGSn6egdn9WqY+00gtnHzCWBqGUClswgJPS
56/853ioWzh+NSuma1tGwVWNp0xFjlkDAaxANT6algQfMMs1WOInFrXLcFu1jFkoVRVE2E+aCnNJ
XlBHSIEDrfWt+OApTyvTtzHzE7IsXQh7h29/2NS2LSmrZhl6k87OCA9DCRCHk/oRhY+EB+5AeceG
Y9dJB5Uk3Vdg5W7gyx2OpUkB29JedZhvvjIflxY5Qo9EbaHBoDikfM4Fj9v4qAAD82CDO6w4hR+d
GMMVgMMtltpLBC46PzBhjS+Fn3Nua6rzD9gOK4sLGUowYv+EVt5i3yiaXIakUzP4TRp+RxL5i1c4
isxsmuLVGvc3H7WR3uH2IjJbnrBJ1mRcjG6DoDiN9vjoxdyrwAJsbP0Dad/QdMi4IWYTKRk/V0na
mA2QIibJrWWW2PHofTgdKQXkxyv9kbrUtAXXfWzKvc/vEbD4uurX99eqJELHRcnlaMOhwyoPi+8T
0skcCbab04NPyLqXyw1HXwMrh88C9raxGxAATNtXLxSEo3UIXkdS8kQucKn00oWP/NP/sO6dJNFD
QkfMUTw7GSh0beSU/0EPLzUwJkMCappdHxfFw7XZBR/LtzCTDYfhK7OLI189w2/XeTKPQ+KB/bGm
yywXo/OfWgdAqmXljv2PEZCpGz2wfLzLqmrvOtHgSmgp4QF9MpywSp9tTxlL6aZGEC5Ikx7OYKhQ
QEFHUq1n5bT6J5VWPww3bnjrgk2HgSqv616lsNE3oO9LN3IN/shUB85GmTgUNAYWwEjUeJQTsAeT
c+300gJQJmjKaemOleeH/sV2B/Yk3v5W34rfB+u6FCvqmvKJlJNdbzXpY05RKV4Lbw5nfcQxmMIj
DthU0SFW0d6TWG8rszVtEmIdKEOSm73N4p/WqheNNX/DdKBO60DWCnev9D+gfK+mS9wh3hZu4Ofz
/M8lEcErv+E1BPXl97fhee9Qz9/SMcUueq9UL2/nxu0L3WJ7M2y7JC+oqW8qpfaFixorZPjPz388
RWYBuvckwVr0j0g94oQJC9v0Fpn+EI3eRTQNfUaNVS9k4ZjDmcXSCfSipr8AgLXtTafNdColcdiX
HvBveZ6/s6A2UtFTzwleW/rL/cGEVTIDwspNus81uuyQCRai/3cehmhhZUeU2YsFfCSLBnjXhj3N
igxuHf1uC3NlTV2eeR8sSHzIrfuJ5BxJcd2+uee8D6LbG64W6sBquaKR/KsqH8dlZJUCY9OFPRmb
GHrOW3O0axu/Be4K/EtKyjbnitCPMwYuRdxeOdk1QvSGYh0UZ2cbN2dSPyg51k76Tbzvj8iOkCBc
rz/RSdBl7A0e4+QzNMCzDm2GavfBy19R60grh35RCdst6cmH9hNbhyFiC6PEhzRVyddPBNGan5o9
BiVau2NraIetE9yqB91sw449AQHQvfO2nsZwZN9ZGfnPO3BgGHReZZYHdAfLUyBIK6CykacGvTb9
kGdafRg20mUh53rXRuPGGstz0TAnsI8EWLaBLzfpfMK3vE12rLmHksL3BIp0//U5efzkZmLzCXOK
pXPsv0HCGrnZY5v6wCOC0ggqYkGFdRaRrx1gZ9Tfvb/u1fOSdgHfeKM5iM1fWoCaGov3F7fLniXj
ivbdIGStfQb9utijg4d7nCUYRhj15tU6+bUo05rzKBLktPHMZ5UHXMHUmfbRxFDCOkhqLfLH4d+X
6/Se65xnT6A9U46+P8IOIBA0WQPuBRtj7yNSVkJNVMacDJv6bRp2VJ222TIq9KwsMRanyVGOEFHR
1JuhKD2RBjmKDhh1D36LrELmDMxC/SK4Vj9e30xeKOWuhHEITEk9kkltofMtlOhtXBGMxZ7yJ5EA
pyNA/st4VLAxc0FJCfxNdCBnOuRQIeCLMVM3sIVcISqizT9IGLSPq+43uwPSdRGbV/alcGkUdm1X
zt3PL79WEErZ5v2iii6XtHrFCoaGxuRwlr4QbHCpA16+3RvzFHhWz6/eT2cCVt28L0kRlykvudZT
X9ODeTZELSfvHUndDyY7kh7+1pKHIeZGIXhfeYGX27vkFaM3n0HoOvNwasEeqh4DK+5WyR0UF1LR
dXs5ls0jI2KimreBd8VRKEtdjfncAHUBBXr7X6VwvgBLP8Cy3qpYld2USX/7GgfG3WE1R2n2LnSp
C1VOJmW3IQF5dJ3SNFq01vWUjVmlkNeN6+N0zeFSFthLJDuSM8+ISwpyxIpfSaQb9I0C4La0QdQj
xNbBi5Kv5aWSPP7uFi9us3LxLPMv2VQoW5JEBGQypR3npQssL6YA6bkxIGMsUoG38GpUuV/gXIvI
/MBYddVwuK2BSrkoZPVrLOJAfYmdJzvmM7tVgIFrBEDRVz6M6+B+u3GE7unHDKtiW3MFAjKat/Qi
hybBgMLU4tOJ+vfwX0Q9ORHYSGis+4nROpDEpbFNSGBrnkBXexIezoNz9eYUPbtUV+qdv7nhC9ad
DS7a1SBRU4DLpb/0DgvsgIU+715MmSLibl6MuHLUTOLVrMEqrA8eEh3yPMmFgcL5upj9JAVIRBVH
nF/6OXSJCTd+ZLwThl8EBxTwK1xZ6A9PtupqoXzzElEXZQJn5/SESnnXClE+iFTiGIfoZRPAG1VO
DbORaGvAdqjt0osisa1REbUdr7qRajAJPwUmXRPu+JdLpuKlC7r/vTYY2TuqqTyuSGhEO6+WJVTV
Q6kUhwZkaeSwQXEebB2EkLAlRlcb7WuMPODkyJJvohNczthUeR2YZAafY324X/AeHy442TGPJVgD
9xmID6FW2Ug42zYJH6R9n8KiVRPn25YggpMVMxVZdjppeT1Kfn6a5SnX1B46ysgmpAEJnJldpp2x
GUgutZjIp1vXw7eMu2padWdzTm6I8C6MANSw6ikhmuTYnYUrMoBtCMpGS3NWSkI5ajMpS7i5L/E2
6nVgv2U+qpzImmQa8zLrxbta6uGspX2pwfUHmYjKG78Y/t3N7cq3aDFf68qVU50DRl4rX1je0OE8
UeZEuC/a+Bz9SIJhSzztXPeu2fvCA5ttWIwuHk1LpLAheAMdeJSpXaX5dB0Up7fBhPwYqjj3W/UK
zzWF4zxL7m9ObnQDK/vmOXT0eWUiOPy56bG2EWmKzQ1hx1/7RqQdL6Cg2/91wj8MalJf4UQ0M9hW
J29GcpZXs/sN3aGFbYMB/fVWGxH7XP7sHrch0gsfcykdlEiwY/O3BmXdrwOHup/moQjwTA5TdQy8
fvcZeL711YMYDBwWBOPhCEmiLiXVzz0bHjdn0w2ylqaEAeuezlrDmI9Sw4jQFslPvx0I34/IxPob
25vsAEBI7bfF7AC1KbxyWCnwvhDRpulK0o1oS+7lF8d+SAam8IuLh3JlRQo1/XuTO5MV40Gol0jP
Ee0i1csVtX84wGUaSFyZ3RV+svHFmGobEYUTv4BFs5pwLQiY2nPopVfxOjjpnS57c5c+d2z4Skhm
GqLnOQ57TL+v6CzqwdK/cnlibSLpGeYnfm/NrZKGGFHmDC5ZBIz5m8ZdFzx3Ar9jsYrlAnqUVz0k
/c5UvlRBcw71JhlZ8TprCLDb5pPXsdz/EKCBA5KhR3Qm7t7GAtMZeEyVIeOe1KsgoCFHsx8VDc2O
QLujBDl0HEUDyVFh6OaQQAbrqZcYUZUD1s429quLvODcE5PQJ7hddhz1MjOkVIC3sBe2tiqsxyav
yMGbI+5HMxckFF7KXCbAMTjSbtE1YAd0l/Q6mXpPtQEYHC9qradJC9V0wVRiymRuGcL/JK1S+7a5
QfKCIbTYkuYJDD37c2b4EAcqAlIxr8cvk9+Niml8oYqAnlw1ClSvUgSrlRoAstQkpZ8Aj5/cEsc7
awwqXqiLl5EreALZjSMAYjeuLZCUmCrSm8PpX3kzzOr/QaRFEjYN2atbFnR6KztVYF+kpviUhtGd
FzG2P1vC3OSCV3v5JXYuRcBu3DDZIejLXzyRzfO+sC2TUbmd/1GcgmfzLJVfLV2KJwZEZz6BQo2z
P5QjSUNG0mBZDEQ/qCI5REkiSG1rvKRDvmn8GZuD8QTOdKOOoHcE31XeU7CgK/1dfLUBWcPXaL/+
K8LYlGcugM+vW+gGMR6+iKG5exWbxDIIMIc+4r+oXKyxMQAJvV9mxe63yHcKHUJFYtng/tvGYEk2
fdjFZpKJJaOMO8mXT2tbJMieZrNKcB8VKAm2naFhZKTXXlByuTHq3O7DZjvc4mEMyFwzieo54SaM
9GOCaW0r2Xn7Ny9+gYIaUQOd11HlJF9Sw1j0gcXhcAW0Am2Pt5u4WXK65b/NuJgNwFpeYfo0cHve
wkM03ce7kkkLUC+mqJEBhvcd/aTZ/dchZCSqjKLsH1AJu+sYR3pvYTdyCpf4XYF+NunDkiTFqSwY
5In0Oseq2uUeJ0XphTqjZHi7SrW75NNdQ6l+i8iGoOuNc06Gx3mTBF8q5r9qvl1bGqjBORaLcU4N
G794hH+B9HpEvCsvXomLJjWWhqVyhhmitlJabM1ibtSRieSZpAHj0f7HlTDfJcbi2DYmYJr2sCAY
RhKhIDXoy/2/rpSY6lBblOuAo4DXutJr94jOotZcitENc4vpMPkwA3OrI29fBmMKMrsZbwihxAsI
Fu4/4+UqAEUKeE8GpPGtjsnW+5o7J5bvesBIiyH/FrddgBC8jAMkw7K4ApuQMfRU2n2fbbFsppXI
IeOwD1jDscGsedIZKifiY+GWA9M+OvTIhVMRQDGvYsVJ/30KvXpY4dURHIeufK0gUXneHpbUaxQ4
vUZOxLUCRwX06ludSglmItZOo1oxioEdxbckvO7l+fUPpvEqjlZ/q9vrGjb3TiHgawpS8tD40+wK
MkEbcyKSB8x7aOY5XRM0uNc6TencDTWXHKTrTOSygGDo6Hw14ArHBwOA7HKDpwWojTJ8KWuuGvG5
Xf1BO4yjiKj6OMkGUU+ksSpkSBK8xF1zqJzLb2RTl4dE2mylO73Z2Z6Q9MCDkf1Wtf+Gb8v/SNMX
c7ZBv5uUsVHcP/+4xXU/AzSlFW3sXp8lYSRfeNl6h3lOa+469psDUAk31ZkVoEWT948nKQjfuYg9
5WKM473WVr2SXKYqHyjatcmuZOW3nOFzq0VXcF+P9Ry9pKT7o7A+wAZy59Q1EV9q+JGmNMMoFnM1
JzXSJ5NRCe0N9QjJHrCLn2R3a/tF+LuXaRGhHzyDxI1YA3cpYlur7Sx+fGWZCByILrCxk053F4XE
iTRlKiEmRPn2b3x7Z07y1qH6qFHFq2UhGtP9gKIOo+wUjAjv3ugiE2QZyCt/ws3H/sfg81mS8zZz
mcoajq2jRAvjx0NaTT3EyKlh5eL/qrHNexQe5ETL3FdEo8h1njn/mjcmc8j66/TFLtx/Cm6/qsGC
6WVotWhZv/8o0GtS75Dn532edfoLum17gGJOy8D7cvbvRcKUjNSgo9miyRH5MrB9DLOsBCVXmHrg
nfLcWtxfo8YhlDy4eiP8YEUCLtuuwu8s0fOqBBQcMWCvEShRSHo2/Q470yK+SYND3e+3+ADQG2EX
wwKq8gidrxWIfdau0nv1t2wruZmqPszQr0UYx6KFWt3oRArQCSyQ9kjFSoEBLQ6ABoC5hw5eEqwm
k+oyxBV+rvZxNHzSBz5/ZXQItjGRWa6AQfI9WuvtE22kaCflS/0QDTtCxfXjHVxX0AN8H2A3LTEl
5zfA+xSfdlYpfjFIZ7jvheVAHlWzrhouDocTkrW7ZbpdgPkiLlbvBtlXOPQBWazSDGF+qD74sPD9
Zanf2lSKFnc3dNDOnfqoA0Ib1KUtNJN5+gPRZXyf94Ld23HOKaLB+sFhYyWtjEqaMo5+aEpwkUd1
NLklZsFy/rXg1BYhhhKNms6wk0IKVayjuVBUP+BDeBbckdyAzQHAo7RTIBy7bCuGeTUcBqMyqGcw
iJDFr3EXOVUBLyEj8UzG2DuINxJivTfakg1zgKyuvjTggQN5rlrr6CRCyFGI4yLzZnA7BfngJyn4
bk7dkOYIOaMExfjvKqV+ktUoqiqlwq905YEnLJm0hHarhbIfON0cCff/7X41+n/6w+FXDsLzVABg
Z8WmRSL2dJuS+mR6OLV/1Jx4ta02rUXy1NqRU/o7560LDtplmPcEksKYk4/jDdJrnFcEf652NoOl
oeyuqAbv4MPxqGmcGqZbgKum03S6cyIxeAaol2utn9oFD+9kZ2OzC3hEb3xKIokbwXsvvLWM8fyV
HB3DtiTvW70WH45bP+jgIQoDa5VI9VnCMRUjdoTYg5W/ALDMzyjD/IC8hmoW9j/6DdwVWKK4s7X2
wWvkBusSbDg4nTq9uaY5Rk+RLVVRRaepGj95a3URMPu2XLWe4aFGi9OYRPOgONG3z25eoAcqfTgG
ZBpgB0V6P5ZcsNT3+KzP2qIuKcjeu314w/5kWHEwi2hAf11dBqY/k50/x4ggZ4Jr06ECcCKBBSCL
GIBLS7yJ/6/KwDTw/yi3W1CO5zjUnYRRXQPl+Lf7z7KSQnrV38G4P3hQdDXU3YwxbcTDL8vroq2X
Im0Oj6LXLFjEebunpnrdmWqQDnD6fVbgFjAA/FXOh3US0YmPc4+YS3AOpSNtpPn7Cp3l6Bw71FDe
cYbdfXaQOzmdQ/4r+gvBHg7KBs0gkR/Nk0QMoWFhlNE61fJ5oirzpqMCzCGG2V6KbHY2K17bxBvi
+DLDqpFNsuvUpuGjVc8RXTFNb0TJ1MdYResuzla8JaYyQ1mjqD6hMzJ1SIy+JI4ICDVzRpQ3w27H
zHMA7gQpzEAsdWDVBrUYckz/jONTgRIZFkUyvxVpmYnxeHPpmP4ggTh7Ssmzb3pnKWRMq8gTTP17
Q4MWE3irZmy4mAdJVBR1ufrR/DG/ItneKkWUK03HH9Xk0JzWVSfkdRXJFGfaG3Vb2N+d/+UrI4/z
oMTj2yLWIQo89a7iqS45AFVTC2wM8Yfi0fxEdhPpjwGdZcx+WXVZ4fwpBh4ELWTICSMMyeJAMTzQ
Q/0W51siaWKtWNBUIUREhPwY9Q+ck0W+dacd6kBwYxFa0rwGLKUWHxtseYB8+kNOTIv2L0pvCfCI
/eJgJFWvSDf0A6YTTLMjKJwYbNZSTKzIecm3y/MqS8CJJjzRr4cOZyaeVXVBCRhaESbBCh+prFm2
MZZXsFV9U2ib7uAfa5VKWjLFIyoDOlRygGOrGMGWV7dWl4kSulNbJphWQsXKUkQ/ZAlp2hO2/pac
zLM1Dnw/gKCszyv3Rf+Tu9lB20dc8Nr/x5KuHjj98zchjJecvv1n8ys3jvPNiXTuZUmhoPP63ccu
oGjse82zon/0HgT/3rsyAx0D1sco/W89ACJOMRIbT85/Dnj4+l4YpclhbG0uHD0Xgxm8X7s0BLZt
HSDuPoy534cTH2czNcwCwYl7ra8SmTEENaKsHAMFAFescYVIlD4VzRP4LdN8eg4xMSzowMIGbi8d
yWT/ET69Nl+mS0ama8HtT+qxaVT8fWqxTij3zRMYLnThTOQDJUtiVGtEUvDDxSYraW3WHpjFMm/D
eyPRf+5K6is22Fqh2kxUS/lovIBvV+CEuu4g1hVy0b6bb1jVcPQ20x9FL9iDUHxLz3OO9TGOsJuc
D5HNxsRYxYtGIDPzLWWp4HXLfvPY/B+6YJjKXIwm0qmyU3GiZVnAnfU1Z9jBtDnTf0+KT+acCwyX
+cXB7RtDkZpWR42sXqF7odicxrRDnK+IsnXGQ5+2PAXnd/Vowk00U+1PTPVani41A0kOA+J5sxNX
8KR3Q5OKkWJnY18ZmCOIAhIqhF+LefaF4vDxevZoHuSaajBRnT1icv20ztTgM1fSoauqMuJPZCKb
cvCJRxlGY4FVHGmx6S73j63Emlyjwp4+euWeXY8YyAIsDZvBobm+B/cCvk3Qe1cZiIE+8VZ9Yfgj
bpdEi6uu9Te/rXpYMwOH7q5/ii9Dt1wrS6Y8kWq+87r2Wn5d0Cr1uVUgsO3qww+Z/HPmEDmyi9SV
XBiHLrMqzzA/0mB6dbK5ZS0F5fsdqPCaIRLz91AxF5WgLxv7ewqVYBr4K9lwwRdT0xuJaFbfpgdk
fZGR+lZSCN+pHItgCdj+NKFN56i2hNXHqCGXf8EheQ/iy9LhhrKR3WRwHNdMkec5QSkuHfoVSa4V
+YYz1IAqQA2UDB4cXJvqThKJ5lzjCqTyGSBYiEDVELIecAO9AfBsfSYI/JKuLSdeV3wTUWx6YreS
dFq0Ft6fpo7o90NYLQAR+R2VYz7oQ3ONnTB1UK0KZW1ahce5hT1oHlGoMIZ/eJGgB4YaDNbA53CX
CduIO2n8AZNo/YMwPNLOUDzjOh0g41xjrpHJMZcvPVLZH3DxQ8+BPwQEtQYMq9x0ffEGWoqKnHJN
nhRHHl6lx1P54BcErNHG66ZAdfG2TVVS9Mhf1tkass5BJ2Pi2x+jbRcEUCD3jHswjUQCsMvmsqdP
iAlz4zW70FBzR4DmfZBd99dpwHxoLGBkXoTKll4Yg7N0k3tELeI82SrkJgRiY0LewsXjfzttkWEE
6DTzYJluuHk0Q62OEm/c08UCh5ky47hWIyItF54p7ud/h3XmCuEJ0u7iDSve5itkbzP7pIGmWGDP
jnob1gydHPW5/GDUBfwH8PBkXT5C5EYl61Xr1imeqSRlNB0js0Y/VgTEka8mTTq2GP1WPwvi7+pm
EEaia3uLDBhMuumLlkrHdkzGUnucYqrSh1T5BwG3fCU87he24tqKRwRmTyJ3jKT0At7vVQxkWp6D
qeJBwcN5lLGJbVttlC8EcPMJsUFbjMuMzD8GVw3b7z3Adf2YLYiBJfOMayevuH4ptGl7zDSASSPr
l6FvK09nnqCQnGEF/xtt7UsRBg8UVgmKrUZYLEnhpVbCk6+E58Nh1qpWdGe+ITTSjc/jCFN529w4
QBxsi2v8SzT90ha19ve0qoOPK508EHAIBGnj2unPKliZH7aSqpHxgF7PbqbBSbFBLON2ksbDe6hQ
MGBMCS0eLMURZ9lU3OxrcRqDW6nGeeFvWJ+hlS41V91WsiR39fXOsBaAVWbRdEP94kreqse9F+kk
wQUqgUyFeCkmGQjvHgSYpUky3rzwIgHm1Qj+bwgK0Z3wOpeepUaEa4yugSpXk9KhHXCuiyon4eRx
LkdylC/Tu1Hf+uE1FrRYN5RTlEc57r9xSVZTTFCP2jLROp9TQmECaPol5FXrkVaKlccc0FOAVTvu
grautzW/1zoii7N5IHP954xML2Sdp56342PxXaJsiKDgEniwJVJy/d7JSSkDxib1bwbCVOMsNKog
ytbhq777JDPPPLZYYyuh7PDXdYTyY1fNf5KbEXXQYBxTUVbYjBDfVn/F+XOSVPb92XcnVdqgfAlB
rPednsIKvTfX8K9DrjqXsp1Dh7wiFZd5gnx5FHodE1x7k0AUrHuIPjBA+MMOSNlZbKmnAQRCZJYD
ohIHMqPq2o701lepWlSfbMEn7gALZRwnLx0TuYFmoyShkod7hrBNGiRAO51NP6Rq4fRUKA4Ds8En
PPyNyFy6oMN3Bfpf8G4K70KL1i3c01/AUxC+41mNi4g2b3nsF4qfLzmZTY+pbGkS3obna5jRTnow
BVOAFO5pV2yXVqsoQsJLkdd4dmlg9/7E77rz8xjpCqLDEyXjuBJWEPglDwjyHLdImhTXHCFCaP5w
bXFRrxoZrHbPrOfaOgXVmkaXBWOQEyhBWgIkTDeFZKQNN1Uo8rzmBU6w8mz7Lm9KHlkqSPqi6Ygq
jadfqdsYLZVtvZ1iNcMJ5jPgscytnQCRS+HNLo8vhTcoHQadRTJQJVLz8+kczCvOzSGSiwRK8HvQ
tA7X89/9+eaAEl3HYwr6AwPwqkcDG7RTPTpWW0aPGQAfCY5zRGHmj6SeRO3YCf/iomBwtSbAdAAL
DmvY0YJtrlcmwuQHtO2eiHdlQaIYpBEX84Wt6g8A+pM+3UEhoXQG9wpBQiTgVjUZbBbn2GheiuCi
T8GKUpf8vCD96wm6WKj2Ol/yNlgAN0tsc9V/zBeJ3FZ7GfkNasakcfXi6tH3fRCPW7wV923+y2GL
rlkJGc2VB5Scvhx+vCHz3E0lDew/UYau0Zj1gjHIH6uKJFPHmabzZFfRZkJ35xh/WSV6FGPox6i8
IWucamZoHc62SfC4ED2YU3wnyTYZaoRO4pVNzqf3M2BgfwZLxBmix/ZRF2r4vO4kAbrFv7vjIzQ4
McX5H6i4UQlwH1Kuk9h9ODdSP8xf8qQwntG4PfM9KNi/aD9gmTmQGh2O5bMPYp7BxuMqZOmZAQ56
sPWqB4jBdeYPE1jyQZyfv/vUCgAhCVy+3jKIznvhprYZu/uc52kVzVR1hhjcx36Bpn4N/zmEQM7w
DhOzNO4FJAs8Ga2HsSbP9T9ikwNB/mcqSxcYmKQbGGRQQdotZh7ys0PXUhP1zebe7LwfPURIo25G
vyx35xq2FDExzHJ+E2fP7QCG/AGvMh4NUDcl1ak3VTjUg2IxjnpZGOHyl9itBfOsp8XIUrOCHGcq
7sLt13/WNBw6qP2LEJ2awnZmffVaCtpZFUeby5Sx7+TwSD3iYWKFCAu8F5Kik2u9U7FvuZIt4OIO
IchuNHaj29pyjb+xnl1QiReOjMTvb2Ol8uDehizEGfj8m6MwyjmE1y0r6kYJmWVJWp0jVbL0j74g
dT2u2SRvQ4EwlX4NoPpm4/VedJ3/50iVhSLT7FqzTA11Qyw2Ja8MjKrH/BZXXSQWVa/1QQKN95Pd
EUfhiU2XjR/lrLQ6v8RrYhNo128SwUOqAA8W9Un3CJ+QzWedr8y/sAKCXr8Xg0cdo+8p2dQxZbrE
vXAdRudPvoGvWVKS+WMdT9N+ETWIpzGEMRPjkZKX+JqGwDSFPdq7cqSQEEc6jf06jY8fwjXOXme+
bb4HL/kQMn8el1t59Fk8In4IGcLEMLfrxi+wSQpqDCpjceQo3nViOWQfckihHDStWL+3gc72c9Dn
H601tUb2LDo/QpKRoeT2R07aLwZOakv08AGeleAyEjiCZ/KefQPMOy+ZHx9e44k6XTmssTjJoMAP
XzMj029tdThG4IwIc3RTqrW4mntPG/BpdFwAQuwqc1Pd4HN9zqTTGW5ocfkhVI/ja7n9IzRPZ2n8
cGGa4+BoSK0tWGnzXjUfmQqcsUIIXV8A9bnKUUcgdneKPRaua7ZhGndEFArJYwxHmHDCCjt3OLWj
XCWp1RK4T7gpF/HEeg0syz2VQkkC1OkJnCCRh8/Tz4dAJ7WKwBPlgtKNygaYJXlf+irMzS02ZJ0v
G7y5OnYLR7CuYgv1P6Wr+ePgRLIB+UnvehOkija6fbKnK7ESDZOd7UkhG2Vo5iXxkH08WhD6urw3
/k/M5MOXbK7oRMIr0LWs6JVMENxSoA+wfUxydX5KKOaAJI6bzMtZihHxMSVEB/hbVO7hbbVMELLo
HkaytLOWNwJ5ayJfPOCRwLaH+ST01Axepf2PKQ0ji79HEwR4MA4AH/lvUEUhaH1fSN/EDydipWVT
HTLt6TkMk8ghuBhtRTBdYuCA0ozs2jOH/2vcIf2aT9F4m+0DkeFqnGD3ecUI/GhAivjmoSgC8amn
4EuftLklHNtPlg3jrG4/BXSEbdV2QVrTFTb39RugyQA2eGYsEC5DZS00W2ajGQhpCKwT/z2+thss
+d1Ntybi8X5cmqSELQJv0r9LiKvB6o7BgOk0OHOcp5UTxiYdyHtIhpS6/MpmY4EcElc5IHWL4ezS
T4sS3FOehP0mvUfpA/5kCJlea3ucHanh3XjjORRd/PuaZTQrILPa94hSAEO6SvWwEbCuBv5OiAyy
gxpg/7uIRvie4awwdKJIe9YXDPhBzDn0sIAAEEEAUT0e9VaehC4o4f2fE2JLiCMr7+zWidAzLvAJ
ExAiBERoo9EawGp7DZ4pmmgyqQmDyxhdfVJ9rfsqJRpTMFc5mk3zLoKB8oZf4IOKDhjXPkK+KOaQ
IDNG+qZ8ZpzLPpEFBXsuJmXqMlMkWv50S7hHpNTSRb96j3JgaQZ7/saYGS9KslDw1dYVlBs/giD1
YdeEHuE01Sq8xhruzL39B+hLvqeGeZtWt70+FxsvOLaskQc/Sevxkp4vz71pyL+5xiAE2+PPuBNi
uVP7Be/qbpfFcW2aOKQCuigvN6kmOQ3WppKC9tZOWS1jZFV34cC8PrNffzv9uBDh+1e2pLCWGmEd
cAXaucrvjEi5GSkCgNSusxX5K5M/8jx4i055FTWDREt1VWJj40Ga7emCa0vRgs8AwXm4hx0OH+D+
IxIj1NwEU6CWwrecvde2A/is9ADIwxXyQQQnk0XUihYnOjKv3DJ5mNoCdZLa/hIQGvsjhDcz/Yax
7g8mN+bVM9IAnsNrAOm5kahSQZrvMSGV6cwReJdzgCvUbb5eCF5q8mVxRBBzdAHUX5sSc8TIf/Z0
hD+eiIoFLCqERFXoEoVxKqtjU3A1IHkBakRJlwdi+3rYSzUJtbuya3NOGeSKqyaF+BXKy/mrGvNn
08utgxRUSyAhbzeflXs3fVNwuOjA/wJx82uZNYckDJ7aqfa05omYtej/AeA85iIXzyJXk3PcGCs7
t4bH0apAZ7Kz7hSDAqsK7xK1vQ4DeCwwEu/POp2Ij4dZjUcrJ6ugfTVN5TF25scCFb6xFst8lsjv
lzDHs8l5r/48pils5B14IXOZf5uifz42AQ/ECnt9HPkIVGxP6d446Dhjl+/AhuTfWhAjnhmFISWO
6az3syEt8kslM8fe+XbtgezUneMHyRecqho0TCRNZgRUEK+P8Qj6tPUOVTzWrnA5ROtdc47lRMQO
lUIMoZkceHnONKWGjFoAkFt4ZoALLwe8246arbdB5+SnPW/ybdbetYSjqp0k/EJSBEr9ZLhwv1F0
Gj11yZaWekESqPOuKhEaP3p5hG4R2EK1KuZ4cQMU9b0fQh2HwDph1bKM2ILVG0DI1lIZ5M0HG/48
RV++/Cg5ozFQASPfVFVeKY8oWnCpxv7M43xZfxo/waMcIGLLDxSfBSvT39i7pFL2hIl8X5j4jY1u
f8DN0IS0x7E5oHKd6a86nGszbujJxq/LDjOmYt4sRIcUnApbcihQ7B9w8DUrQsvSISpi9TrsQm4O
tLH+PSGbxrrRDRu15PCBG+fWb48MZzo46qmXoNZdz+6jDPUhkYTwvG2rY3PmXIdFV9mmg/ZCtokp
8Q0CYNpQhZZyhr8cdQg8Ney1sI7/EUUvTAyMfF2UBJU+8yUG4eGcR26nDNAQGVfLafA181pTd/+k
DMss0OhbHvOp/4P/utJrYZ7A2t+kOzZ61fyROk/OJqV0VgA4xfC2dfzwbCzTwz2OPLVrr5b0BE4o
wO0KDUaYvvyHakx12fahxA+Rc40+c84FZ7vEsgP7XcFnhpJCOsUYrE+vLWxTbTumvs240TcAGBDb
gJMliZi0uaHuZ6f1BNsPP88xQvWAqvwdQxkJCjvpp4xPB050ZHX4keFhBVrOiVVxUzK4DePtzNC8
Dcdry/q9NwqSJeRhRH3YjFOzoUNFQsXv/c4JYQeAOloUIsBXHcIYLE68BioIvZ0Sy5ZjiWIQKycH
mQpG80edEJ9/xxQNqXj2bOTdXs7AfMJJ+eTxr5p1Cc7rn1lsR+ctjeoyuTq9HmwYA1ttlU5KjKfx
czJxWlkWVj4Gs5AjWaPR62Si8HhiPWvJwuQCmXWYZ6PCuNnAQkMiSzOnZBz8nx9SHshDxcniEuH/
T/OaoOuk9wFlJQVyppPItQi9vJfrjr9V9vA4O44IUHvsiqycM87udI+AX4aCDRRgodoQMDPtwTNf
6NXAuiTF7OEVFYLKow+XX5CbOX6KzNeCGiYakM20hgmLwu56Tcc91j11DJtfkdZ09UAUiQID8L3L
7h6jn41BKMec5JOZenQ7vmgwOTAmfFeS6TOpFOe2inO27zeDps2oO/CUeDiGyK2/PGQI+ouRWvU2
N12zzjA4x8EdpEfx+peb5cbhxnELAcGoLzWIJgra75gq3hhKvLRVbXLSL4cPDD8bwRR6vqcznuk9
k0HO6iZiYTy7jNlbDwfjM5Ddu3q7/PpQTIy3FuPJ+OoBfC3hTy9iL3QJ5Wv6z6ourSLi+DUs8vVN
7nqYWhTX4j+A2xWXaB0g6liGL83vNdbbkaqTJor2M/60xvGDoXwB3G9D+hxgQ1fq40YA7OFtI4c/
mkcmBc4FG5aT9qtcpe4rxyzjt9F7yuRBqp2szuq6tFYci7/FGlDGNKcSosHvBOzjWGd3KisYpDs5
RrSp5Ytn47EyK7VvW+iQGnbpQQhsOXHeHuPvgYzHIIM2ihKoqfwdZJ5dgjZjhOtC/jQRDO278mFE
1tcsvLO7tzY7vFuy0CY74ltrrJpq8gaBgpopY+Or623IvGREyfVYltFp+ug/+eAOgrm8q0nkLpBG
8SD8ZX7jdYIMMq3lPMg+zjMkXllZOuAHhxjrgzu4PLVVsUYUWcCuB30M5QiYXlrEU/CnPOHRtpiL
xpYoj8FJto/E4gxEBl//qZXTzG/S4hmiB9YWPmt9BseG2Zck+69GiMU3nKLN0VjwYSflMF2yMZX0
kvFw/4ZXZ6tvW8vLobbMcQCdGqNzAfm2uPTTd4C9+nsm1YkL7Bhqi3Jo2juqcaKTHuXtx80Xpava
gu7U8UC0FEc38Faa14OEDqUPogl0Ipun1+yBK9tkMBEwVtPvUEOXwNgRdrcof2CTHSlMrgaMTHOH
5jeKf+UEreT9Yzd3KA5+gRGvXE0ukX2fkc1JKqa8YENV4YbbOy6Y9ZXyC3/LJmfS1gPy4zU7+4H/
NuJ1L1SQdGgUfgcqXY76yx43PPITyUBOOA2QdLtc4qxbW8v9+1N6wy7VbWVNRyWM66V74cLUZg9j
6v05PT5vDz6SEFkQB3X/KXYrOE1qUxRiETMCLsmQKnRWafvFapO6ENs30EkDzQhh8wxFRB/r3Zpv
1h2x3qSujUyY3fLI/Na+5vdF/NQMMYb4N31YzNaY4XP4Ti5EsxxP0n3/Zk6zvKvmWJMbTTjJDDiX
zIiwUPyLtig+aPnvJFY2yKjWjtLRLI+KLvz1mG3iIaMwddHuoKtGSHcg7mBwI8a3dh7SXOig3C9Y
HDsP2yzuPuEY2/WaDU4oNON2AHEkjrId4MdJA7O0mZlpFseczi2tfJxwaQKupz8GRITeBLCBQUNX
ragLa2pqAZs9Xo6elzTVFNsJlGzMsVKOjgqwOhUCf1sJrPH5Z/mJ0jzXOjjvIeNdbAtq6aZ0VUvM
WRNTG1q8ztn7frsgVqCOHjWAKTrhv8J58IZ1qp1kpuS4LmjVQXEyX04FRwzRqm8j5Dv6bD71mh4m
mZMRRmYHbP8nqSedxKX+ux5lJol6bPoWdXZ6Huchc7iE7hsZQxc40vhG++6LwzV4GAzgDL4K1Zbm
e6NdWFL/hqVOeA6X49qPEdFNgCUIPJW3i7Uol86+7Evg+eu8/DOMuKvHXXN2AAZNOFyYgz8Bnv4H
oh3zZ4fQSTCtFpjMCJKL2tCQAyWXITMtsmVefuLaKnY9Cf4r/62SYxJeqasGeanWmpeeLz+FhdFB
4T6uVAvFh7aiZchplNVyzHfyROBSb/obxAvIyAwhpiF2BLr6hSFPUvjSKmZ1rTXeiGdw5+HiphF6
K4mTgUcPjY8uWf2xSW2fhi6iIHf5qUpky7lRLrLiPZxfges546vA1gpeHvv0KVS2T2xkJZxR5LtG
nFddNa6FVK7EVh7C9Ha+LJt2a6oseyfs7LTZVh+mokZk4CWJCVHVoDtSWWWX8877jKpnUnr7xGKd
KDq3pXMmdVYe0vDcs2DnP7AQfl6vIK81WjI3op+BThf3I1RH/qjuTqgdGvPP6CA8zNAdJIw/nkon
LIprQe4eSA//i54EKt7nW+KHzCiaOQcKfN/UfqORCfXI37YDtyqG1YvTUmq6xwD8PR4joXdOjmqE
FGLR2xGOXfVbNJjKeFqTyemj7lMGN7hPv8OVLYsMRjwN/RYWJlVfkhyVwTwHoL4+Xv2DXhn6M8E5
ybTEcD2yoqixc5QdjzRH56O5t6Xd3nmdsW2meyUN3lMttiFAusCELyvisdQ37mbBQZDkdjs+HdBI
2cRKly3XbR9sxDym4YG9XJCAvZagGbGlc09UJ4CPeBJhZn1dH9eURTaC6/0aRAWEeVV0r7yVfpJ8
N2hHtdJvMy+X8NgSore+E7IMAu+6dKktUAzv6FuStwV/hDQbRG4v0/mgJXqJN7E4TDfYBqooGRZ6
3qVYBnVM/ckiiqi2mjZ1pM9JIwRwl4Jl3I/PS1xuQqlpgC6HSB7PJwXPyApJEIQwJ+/WGNNeW9Cy
1Y/xkWZkHn0IE2Gu4CufjobyOjsdk/EVloGd1+VMe6DsQ5wwmTpA+p7+0qeQc6wMdiruDxNNlPby
W8S2o+kYpO2CpwIOCeyt+lFci5XjrcsohH060sAmHqOVJ/oW20prVxbHKyL3cvuNWEzZfQ8+/Civ
YvWeajSotvN7Qi4tX4qq8k5O8g6hGZgC2AyQvrcv++gezhy/+WQfddtXwoORAWFV7s29WZbAfNKD
8atXj5ttNsx+LCQjSilHD0uUkikUqyWMKUzyxQM6alKi7hhif6CH61dzZi19w0aSwIcF/ZCVa6zx
idtJ0KEbeG0uNjbbPFE7Y5oi9Tjd09v3BHX/04oNj++zaf/LsLwBuwQOfC78jiYhXd1refQAkib5
axq4lO2icjKBTaSlxdjNnkA4EeIBaUSE+13H9pkFMAEzCm2pP4RPMi2awF1aoSbeG3I0oITReKyb
ELCUAS/VZbg7/ZDZBW2cI5VIYXCzwYYluR9FAP+HXfPkBvS1GTkqVz8kInuBXkxklm4mZYZUWdmu
mnzpHwPlENkenpnhLDHnQQCwq6KqBsJrMx6ed2Ub5tNzw6KB80QhEKjArT5ig5jm534/c8wUYkAt
hyz8XQXznaeRbwD+pJKio9GntSMMH1ql1gS/r6qe4XEazaSilcL5CMDxkAo/TgfonJ44CvF1qdN7
aVZZe43skSt2oQsmcikLhc6eRpfPNg7V8efJEbJBGr1Wb3uUEa3DM9yJrrU9UU12sRrXH9iriNPr
zh4Prm+voSRxxpBIdB6wgBvDChvYRs7O1Ge3w8CLpSmfnEuHJ1/cSzpuyj4tbrpP4SQjuejkBjKJ
jKqbE2IPHGKd+nspuQDq7yBGXyjMIMK48Rsl1V0lHCTiUI5WHrwBv0O9rNke9cjTfobh+F8+U3Sk
CoBbF80oF2cEKveULMNTSvR/P7ENuwCn5nOSU+9mWEntB/Z49NS+pGOrVxgt82GytweyLOEiWmjl
z5lsvEubj3j4q+JxbC6ncNgVQj7ETRCvHc9vREp0j/oYSTthTBHZgov/3MPMoQ2ohA+C+oHI7ojp
1uKCryaKsXUD3PSSayIgRXhlkCti7y9ph/LZesXp9Z7VyH3kjRIEM6rNgt1Yjtfxm1LrpOu9lz2S
khOvm3rrtuWXiUgofTp2WaL4dFN0sBKkwxs4GjdLOKFvX+F1dJghdwoIV2gCvQuU/P129xXG42NV
a4ACfDnw2uZXYlHZpmaDnJUz84Iq+afkJZ880d34YSP16amWOh1dlhfpYEU09/gH43LsJ91R8eSk
ydVNDZignQmE3SWz1vbrcCM6Uua+M54Iy12+VEtIjrw0nmIECE9W9Y/U+g23dHSV4COOtSnIdzDZ
0gA882vCR3BJYhZUBRjxl6mUshbtkBO/TSPTOcyjlfbhBW6E+5qnAP4PHrZGpW/u+owq7j2rsyEo
1K7xOZIR6mcSPPWST602Rx7/EXM832WWa73lfpeX2I9M0sGDUOljLgZvpqwT/6MJOxqXVJRIOEUE
uI8ZxEcKGJjAj0xe/xOjIM5WOHkflN8wWNJpswjwcIi477qBmHiZroAZTFSPPexdP3hul1ZpM4Gy
axXCNmmomli6Vf9QK745a4IbFcGlCd+V70fDNLAAdArp7YK/UY3LoH0YLTzAsTX470VtVmkAENQB
hO/algYdnATFKTbIiimsjJncQ5+ec9RbrwcfdqXPHKTd+Ynu6NXQOjzDqOq2nnO1fMbKtWvUHcOO
p8xwuS6YVaOoCZj3rRcX3soeWLUI2NWQq7jJ+1wpDnm45H3XFJ2wSRpoL7PiRb3u9N+NiKEzfsHs
iNYIaPE1ggjnQH4GG0J6N9Oj/ss6in4QP6oQTC24lGSD/qfyV3UhETT3Jq1OqfkHgLFI1vtjbEBN
LU66/a22z3Ir13YGly4QzvLwJpCTQfaezTlGsMfXX1nESne4z/xlhwoxacHo14u10QXqrEqBq6kN
2c0jB58PVisSaGC87eupUsZSLL7JjKPm1frZ4+AdpOfWvalZIY7AQRixpJvoDTpL51yUCZnqmbFU
HAgXokYTj7ZMHD6X6soOg+xWMC2rl+Yd/K3pluzxtwl4RnV4XCax/43ugrQThlc2n8MzjyKZv1aU
Sio2/krBkdxUzrCmFirZm9B+OF4eHvQq4LFaEe8VX9H39Gc3R0bQT3VPJisJmyklfxbEeZOv1dQg
PpZ5ZUhTmg2r+xTKvvjPX3MmtgV6GclF79mWmq/TD7aJePZFd2XhguSIP/OkO89QfT1V1fbWr1aV
MUOrKmBIlUSb2wVTaTBzVqczV1vn8ykgkNOaXAr//uECGzj9/ZT4yCrvfoVkcJ/z6NhH8tqrF7/x
oieDgzGKErUNpc6mhKBT5syn9bqgxgqMYxkFrLLMxTJD7flEI8VodYSVXIos1FVmR4PuRJwOztVl
tSMBhHdWeC/PSUnW344lAg3uEjuD9oDNbo50v17PJBadJEvif8jYAcHRP+vteREbxAzex2PMYNmw
pR7wTGzz7bRaJFOUTMnlcBro8lKeo1c2qP+ANTJ9321UOLRxfRcRVcXGWlxaPPOE+akrzkJTb761
NzVpBELKUcfQpNXTFjbQoFTst9KLVQxGbUhkfJg/GsFiEntjn77X2WZZl7w/5knJil8jzwgUXE69
W3VxOmRhlEti4KrU19KTdsW8oMuYeES+5jAgyJL0LT7N9SEKaURU/i8+AyuY3Z35R1mlMO/JBz0a
Z6FtE4sYLuEonzrSupDuIaJe6poIcoScIsm4cU6g/oAFKXAueb6DS9RtIx8w0RR/Mgq86Qg7Um5s
FjNVHpf7CH305moWpRJBfDF3xABiQu8YzZNx8gLOhTy8CFc+3APLqtn89iLcpDRg/VZCwP4ri64E
b7km8OO6zTJCkeMDU1JxOtbmh6Xxam7dTSmm7iyEkmB8oSQMCHCfaCtR5Hs4CplhkWrglBQJytCp
QwqA/Tsny3s+1yIwQPYCeRZEQKKdgFJl23yYv4y24/EbDACcp2Tv6m1YhLP9Xk8JGa6wjUOp3y+z
KcZs5sj6Gu7sEnYQufbHdwXwSsDFjGqQzxwkZGWVagTnlxW8AnhBBHW0oU6OyqZ05sJi1QozFI38
4RBygdf5gzI2lFXGngkxl2oLhKr0MEk1CiP09YSr+F+15oWFI5fc4S5egGopinRW0vqOzNt+1HFT
ZcRc9HGzOcx3Tsr7zOj0me12HKs4/hDWZaxI6kGLWg5eV0o+prXukUicunCRhqaOtZqTTBbOdcuL
FWwFlqIqx7Zd+qOyCiDzxBhQ4G8ZxQd5BOG7eTn9dGEXYJGOIqv5flBSH6rejq1t2/yK7h0Gzo+e
MAOFTEzLG4exSAEkvVlEoB2HdCC7ynuk0jD60MFSA3VD9A0TCCgvM6BOmbplgYVM/FoDd3yHUen6
VxImD2kyCe+5ZQkbl4f7A8MEjQuZr33fUmAvubRvGWcZ93u9CGLZQnj7yvO8ljjZyco3XZ5DZeVu
2SoZz19Mzq/kxt6mLCjBAvoOoSDR8rxyOKaIdkR0yC0y+J8o6LnedCrSHrEKPPmE01VTrWR9fdkC
kLmIiXZZ3eXj6pSmKx4pzcq1tvadRleH35+bmh5BeWjxO04xdRhEX6CkYY8Rk6FuRSyOJQGljKTi
jUWdtAMxwAgHkqcxR5NwUc+gKQyC8fX6t4E50SJ0XMpiF6gywlA/tElgUigdx0ialxxySUMZmGmW
L2KsEtDHh0NOLP+uT7F0ULqXKVea8LHZ9XzuvBPiIKU0xxbE3GS6R0TEflz9Z7fvqtUl8guqajLi
Y5xCLwK4gip0oDH1i/BwrDMez5FahLNPf3iQmJt7y0dNPJ3nJc3zWGqnoqsgA0SubpiM1tBnkl9k
bqPt/gGff7dn7/p6A4Bm6F2o8IBaW+ZAfTIl2O944oOrUhmnpSqk6+Wv3gjS5Hz1ddeAEIioLNqm
cT1TKPNY6OHqPye3i2gv1XDtjU4EuhOfXS32vpbp+XJrOJBVqi3W1FCz5PZe5W1Z1cAyYdAKtFsh
0fFCS2iUiLpom+B62kw7/9b3jo6Mtc5/RlmynYsArU3xuWWaVd+aMjZYcK+OJFSM7kbd4XvTgiiq
vVUJaTSNbSRf1rV3C+c6aW9rzkhGyVHQUixYjobWXd/qyniOOq8/6Im+C9f0/HZDMPH0tXeKAFow
j5RdELX61LVi6idgiLY+XicDt78/XLeRvPyR+0zCJH2hK9kzO+aatqFqFpyD8ycSrCXG5BUD6qm+
EP6dMa0NKPU3pvkr0os8/11PiSxkXw7hLg+AFGYBiWWUrsGow1TKpMpyg5Wnw/BhnuJ02cD5B5q1
KpXyaMU301A4YhLh7sZc5MffARtilnOi2D/E6IRPOO8YhknaRUB+/SkAP3CQBkjs89JZ/bGeuUnN
prh3z6HOVRdwCPgMQHCU3dc0yL74tT83gV+gMYV60lZmjqpOirfaeWx0HRct2yqkwlKTMlFF+0ug
K0DMnyiyTZMWoDjB9ct6syBL5UGyLWDUwYKgCoCLBd8P9WbJaFeN5AlhBSFVDXpBWcu9jYU6W4/+
QI7Fbxz/lnPqfSnqpVMLcXC1tC/lj/RpR1j4EvVTW5I1a56deotL8cpVxzzyGc4IqNM6FYx+mGRu
BnpuYUqOsSea8o+JrAKCS5ygk8jse4namIYW3/7gRkJHMQ+2H9G0yBeQB7Jh7EwmDXmIDqeomDPu
Q4vpgZZ1LWrFml4tQaJVlVlXscuXI2YjpYsgecLNxhWdekKCd7aktl1tSNnnd2+MfJPM0KXQ9RoU
URIX3fgXF+umI5IWJYADPehb5EPQpGi9mIn+/UmCqoaXToB0VZXJ+oaXEp3cbbSOyG4I99bgpivI
FMWRXdAEV+aMb4Hvxf8W8N4dPUCRk7oShlhUFKHk9ZKYt23HGeBBkNdwbUu63/vRO1CDQQXYgMr2
fSjg110IClbOY6/VO/BGMXrYmUwAhGR4mtv/kscLbmXAYDbC+0MCcl8gIatQtjQLo7cCTpPDoDol
LTUN/s91c9HLiDZsmmRFdCdYtYvFaoBE/XOHxonUYRdHDYQcC1i78bef8juueAs+Mdts6622T9cf
oUC/p9akO7u8hL2CtSmHw+5XTUuxlR6+hL+4BM5ACVekgQqVNrzVZQpWU6xbTkMkiPo6KCZ9dcLk
QTrcGoLpMGO+W6Pg/gUVdWIr1kV0tDH8GRl/d3WeoHI/gGloByPazepUSyg933czYRORPNECLHBY
XyNgc9leJW+DB2YrvtN1DzlYxizQcpkg6NgjftHsY8Cel9j5OLAki5XaM+bWDVqL8arhTNvl50rX
GbX439eQjTOtixqgR/t41sqsUNj/zRu5vSq5gZR2gucMpHYDEihmUkAXuvy5tzj3CF+enyuWINat
UXAfJAEnhX1OglSvj8ilB9Cve6to/+aWKelFghE6yEmHfWiqZr6+pDtNrUk/zA9HDcR77jZauldr
dxXRsAieDk5EQ6Qz7orIWNFSHmttKj0wveh/UocrDTWV8cV9ia007Vr+Xd0kgPStqh6im+6Zrt3s
B254BuKekJXb+plhfWKa52mDIzPPm/4tnEybRb498lX9l4/Cws73YLpbXjShgoDoNXQAb3iUUc3A
bkAxCvF6WHFp5TU0xrEOTjTpH7SHbhV66RkbA1d1HOaiIWhu/6y58nDrxy0IzRQUF0RaTrhMlnXf
Ut5qrwVTZa/IUlAikckfJFq4SGhHY11Sn3H9sbgp/6bPG8kfnzztbWm5hkuhDUVEXZbKyUQtwwr8
GZup2eqJ2f3PlsMSFUg8Cw3zUfdpO4ilDriZ2NAAam1ZRGUZVbnsz1VHXx2/MjVKBIjn04z5k3b7
lYp2w4IY2buZjO4QGy7FS/8B/tz8I6NYnWCTmKeSrXj9lsAO+Nksa8lRV3HUnzbNhhyWzqtawt+g
Gowv+asJC+AH+txuj/ngReQKDjk28wIyPTwrvnnrRG0n6Zy062s+YDNmtKC4tI3gjd6ta4mKhjXW
x/rsc1DWafUga1HImcv1wRv9rE6xTXMGe7fgPnotofZLbAmcYwxKNZIUJHfmxGKPWafmRzEST6UW
IwDNT/1STgt8t7LUEQOtyFCcmHD5k0gYIQTM+gN/GS8ejGU6Esosh4JGCaFC0mz++BP4TXxfICSb
/rnZJsFcLjlvib6RySCPDWElqCHm6lulqyjq6KbERg7CbckQnNY7rt6fovrffVDrK/a46MGP0N7W
LrE8/CHapQoq25WeiL30hmdPsFcImhbZCw8ktJjwhUqYUQwaghn9RFE7mWA+PhaKAHCfy6tX5HJC
OccWQHE5AkeKlGfdDQD0uO8RkouYBPgcgAqqv2cBGeWs0Vsxyda5wTI/YEuK+k+FqVYhlHROVViW
MpcWazCe52N96fQxS9FOz+eIyIL4lR7YT8y9AUhcsGxh7MdicEk5Yopk9bZVNriAkGhoc3SZGjVP
sbGKhv3IK/1UP+Umly0iYC7fUzJCog1LlenZXPs9Dut+xr+kAi8vTJEwJZ4FTRf3f2lRhDX/eLcv
2IGU6w/ffj8JbdxFOx1ZzfFVoy4NOkUZa1xme5jtW7l6bwtA3cKrnzynfnmG/JoWhBkt2F1jAAxh
GRbG8BM8PBkA3nx0PMmhLs2aYL6PTvY4SXyeX1bW11EFnleQYUixgCRr2SEHAIvCdUTk5LngLc1v
Af5g78fnPCWV5JBBXzec3TYwjm3nxG/fEIT9KkFlphIPIikh3kqpt2yv58EEf+zUm/udlaRsGG8Q
34+JVcu8i5AHAyIjBMqQMx7Ru78d0ZVkofxjUovE/yidQjB+//dRbxDSva+Dd25WKkUKwAcT4Q9g
+zQ4oUZzFXwnqa4gz8QnKWTPzw6Sx0gXT4tGwOxxHytpOsLyOjl8KEBmolnePIlK0/UaMl8Owh15
tYtr5L5doxHj/gQFdbXlyfJE6sNrs5MwGjlYDs74dBPohJ2JOo7yAZty/FJEFQuBT2pscIgYmFmd
ReaBdK8FXzhIgjsNQMp5A+SDjm4Hj9oZOEl65jopD47WJgMCku336cUfaIpTVkGA6eiSWipToeNF
w387pZlpuEfc9UUFVx4M3ziCTOdxipMZABPPCFnefLUtvaJ9RUGuOpZ2OK0ekgLJYvw6ljLc8QOP
G4dZ3mIEaUpFVULsRqYmD1s4jlg82OD5dtwOebNvg1ULjqkvxHjPCthXQV1Vxtqmae4lhJHKsvj+
2IG/vlku2WvCF3qNrVAGpycAaH/tM5nV/qIVL5LfudtDtKJgrFkMk6XerST5LT7TeYRlVKMzmtYx
CwzJfU3hLKqGtiPV+XPM8npJlXwx4vlvOrioTAu7VXwDx+3tT5QewQdUjf/RKx/RYvfNiarQwrjG
Y1ug6p2RAUPjQJd41M0oo8XIeJ6giO4igasehtQ0KhocmuU5HRxpP1vUzcc6et/hvXa/QvLY4kFf
lo+6w39hk21fVOjb1AiUoJMw5nVoC9y8MRrVH4wfFIzARPuUMh3RjZXzYfzoZ9nrmM0EkefvyGsA
9q7LQqbWJBfWrrGyjKjSCp8f2qmKvMcba7/et/8tArgwGxKHbPJsZ3A3I9KvfWzM1E6yUo0Npu2f
Q42AaBXaMtbXlu5O+8r+BW78ujBWOXRygfhMgcOgtaSZ7uD/2fTyInq+K9Nup4oPfso9wZ0iTmI5
8ANvXeD5mCMASo8fn8DYC/Z8J5gEUlasI79QYMS4V8rLnIsbR4EElyV9RFjDaUJqqzdHOYxEL5Xw
5YZYuixcSs4VpcAjQczMWoHZRdC/waskCuEyGypeEtwzyHOMp2FRc6BhcT1NtVNDWaZDcy9KN1hF
hlV8DWI9QgpKzf0jE7m9nqVfXZDAwFThiEpifaxLjL64N0Cn5gXpdpTgRF5zEIt11OUU4DzizveF
GBc/wA2HIVR5hpDhr58bUnWLAl7doxAUcgYW8IDiOoCi/67ZqUAgmnIM69UnBaQk7C1C2WfWKILW
FGSJA9uvgNHU3ZSDHzyGPrOIj3UhpwPR5AcPwDFMR0eSi6M82Qc0U8/Yj2OCSPjHInBp/TWuGRCE
V7m9y1Im7ekJL6Yo9W+3JXRejnkocubUWMQu9VimHNpQMO9ifZ6d14PO1Q1zIKSU5XYSvUcNcfu2
9ea4jZ/WB749qmCuOPUxjPdb8llmgIlmpioOjy7oLgwKGfUk62821Z31r4L/76b8EHv36F+6nkmd
7hq+Ivs9x6MIKLr6IHMGkkSsQ9lrUjQPKEDQ8//P7Qnv3AJUX/0425mnJkvUQZdjBcXsrntZWds0
CHeeWMJvsleFWZWWZgBsTqrWMTTrwBoQbpHmvWmCp9JUA73ZWl25eB1jHHJZf2LhEhQ5MuCNWdS+
yo3oaW8Ce/Ri5EJtTsGoON5OkPvgWC4VbeevgajBCgPtDRccvY1thDG+3FNLGpuzEExDBEQB+qL9
VkpqQr5+q9QS0W3p35t08n8XzGR+rW75BxqHpvPOKeBOdfiJ9URMgfXfAGgfxNTxiRMhKBdwMFUo
FpHppTP3Iusm2SVVoxpwEakfAXYITqhPG0ZKqcLNIpf8npV8tEKxcl84jCgFZDyE2pv+Y9gm6+u8
6qs+sj81cCk/eFSCvqJBBNOaCip1s2wdOPFGTwto2U/u+FM3OxIyTeEmA8E15oVtfv3Fxcq3RmA0
iBUB3LzzNpzl/HpVBoswNP1YIsJRGIg24NFp+MfOGNZfCTQMYX18GQpgW+kGcd5zqYMh7woXRgH0
tDp27UIXMoxXluYzOdnto4y55mi6o/qw6bDKprhvrhv68Tk82wKKD11noYtjLYBExCoyXnF0b3vz
GntrVh/VcPOZGIPNhbcSw9jCJMjsATprzY5dJ4rvWqj59G+8ZFeE06qkkXK6GOF3Gea/fCG14OcU
5SDLYpIRaBHm7kTVXUN2SOkzk2et7IK+cOESOhHRoLDeNiknJ1LU3Q3W+v1i1hehdYgDNnRMA1oO
09pyAKdXWmm45Llt+qwXqpee9nuk46QNPivmB6eKYJXIAyD7K1p6ZgwberdEEyde8idAWKg/s9aH
UOiLBIr8O9du5zfebS2zaW/Dq5vX3M1rzPv1qlSZeKaqyWLDEJKokCPk2g2aHWoKU+QJfKoW7uUG
p5zXonvj5VlWr0yjt5lO+TLHskbftCj6Fm0QtO2ZRyNJUK9qErxD1wHlXFXhDnzb2mbd+qJscCQs
3g8Gsfvsxd5Qxrklhv+shV0tra2uSLF+BzPL3sbZQTVfmMPXCN3WfaL+xfwhT5MFC6fjy3BHuVbD
i34tdmzWueyvFlSgfQ1eglnnfKPrXtcy1hnqvsCL4Ds/JMGmy1k+S7g/L4tDQgeldeJenLesdlPd
KwM0JIAwyt1BkONkDJXOiyCz/dfv+OZAQ9MO8PFMnxK7rkzDPxV3r5nx98hkrV8N1jSBBcxf+peo
UfQNtZ81ASIRbXJiraAN7/rpwjKW6ScLomCuw/P9C44tkG3PEXbKO1VrD5yL3leUk/3D3UXyHHXb
AlOwHn33l+oaFWyMRsd8k4+bWYY3TS9pSDB/gnGL71q2bov6w+fO67U83Ae/F1Dq0wOkzRyETBrE
HF02SLxvTyujaO7ZGk9+U9hMu+4293FBO5fuJBkWoy4jPPvKFRo2VPNjIt3bkdNtHt+QGCQvmi/J
UjIM/X/atkeR9hknoFZMdAL893M5uAwdXkZKoPcUUPUL7vGulz8Ib/sRKBRxL2JSZAZsdQ5GeMOf
Why1dbhELMOvYlWJI1cEcnu4xZU3+7NCuT/JDL4AbIhxgRGOuFD7MDA9eTntnTG/4uUjChzWPEV+
OqrTB18NS96tLQ0QsW/30OUI8FxNQ5unhEL/4fLvFrhMEH8cmJMoD0ORWkMFw6Cw1QdL6+KVlwJu
xVsLp8dBQlzVSfUkQ+1Osge2YPdwhABw3puyRdYoIpHgTpgeYJLAYXGeWv8JOdsum+s5pGK1sPsU
NLHiWZFqEEOCY/oRkLsfrllrbOEKhlK3weLPuLp6VYkhMe/AtXqTHEY2DdgKosovAnaCfx4N2cXG
bLiKfzT93LPrGwlWq2gv5NFQAob67pQc4t0sLkPxNz72JIw54E+4ffAJAgR32IVNmYuXpASkMF39
m4BSdfjaNAlWY/FKURo0ZGKkMO8IkHsChuOvwr9ViUj317x8X5OlVN9RSmw6TppqrvUthEJnzsjG
G6szqONpL64asR6ada5XhxiJZxMs2cPnJi8VfjuC1JyhE8/oybZBWKO7UAN0icp5yh233r6Y6UcZ
Witz0M5U8U2HT+Os+O9oc3wdrI47bQ8aNjEjGOp1RCKvs1rZWVvm9LNPCM7AgiWXNrk5dAe5vElR
a69hWJUyxOv6SIAbC1s0HEgnDoCaPvA7l+suqHyiIpwM5jHopHQbeb/ghEKoVlquoxxiQUf1LV+x
Yv/rkzrG89ZR/fuCM++PxQ6aqa2ksjN6+31S27afSabXEyTlesEPWLylkp2AzHCkBmX9Zf57cgxk
MmLkupeJ/ksPTN2vHEDj7e26hb7TcFs9aHGCQqGZ1Sya/qO/w11aN+gCyhi7BdusaV+ijDASZcCT
6v/6Px69Mw/N5tCaX0R79hyu65pwqg6QCan8U8mkHdNr2h0VpGyPwShztWvFmyEVN/RWvEvFS4Ob
Vi1NEqEDMkEWX8laOPE1v1fPhLtj220bxJggiyO4Jezr59wBfD1e/W4JiEUpkdxEvihkSdPrThos
5mN7w2uFCoZWTUG3Rb/izCNkGnlfi80P4esnbZ4AV6nQ4SIPwl3iue1yWmUjRnnMhygg4Bg8tzFT
+yQo94FN56FOEy8hSViJB0CjL/oWUQ8WPfBpnhCCX8sjbK3agSlvlG11Szic0V5NmvBva0mwwqHZ
MsC7kKYy3pOL6IqrHEC5M4IUdBnCdgNcQlbpQm9iXo5LDTos3D6EmI9YMvg+y5VLuzCzGFcvypZl
c1/YFBDynI/HhM5gxtgNztIjpdfkBTov2YnnC9uxeMN99QjEv6NiYMKVx2Yn01PdH5kO4eJ3wgR7
LPh74Fqk/zjcumdG90DZZbHOs+UlObyWBx0wFoPl0GnlWg8zrEqVqt69BD2bBS7MD8uS3Bts9Wqu
lx/276YAys6LOm1UaiozY1tWm/+jBiUMKLxq0KV/raUax1EuvZzyWRd1kzS+X61Iykk5sBnYudtV
UkU3HJuGvXF3jOq3C6goGTY/o2rFJhkxSANK+Ta1OmVQyTlQ8MyFCtW6/h6widUbfqJmmpZY9y6Z
muFWOkYo09nTpF/m++BV2bSB1A6qp4G2FB6iT0ACYM/tVekbltODuOh61u5tOo0TR5IX16A0Yv3b
DuVoJbtjelLSIqrsakFhj2lC/RpB8QQx6USSNQn7dZvsIyD2ArazCEJzfov6KrMyJsYE9yTo1Cgf
17VytN3xHrehAj6ws7hQrtSemZsC8Rm3B563JHjeyegjs6pEqGABuVAylRqIHPcYXcbwmH9UIiFZ
G+UxpbtxvU0gYWTCUlxrnPQKYfSPY/JjZWFREXCe5GBYOWEt69FEQKt++TqvPO1c7hleOtfRUYmB
Ed5srFQuOfjl4DTR4VMvaRy+OSR108vJIXxL776Vfl8pj6zv6E4jNb1HaPCjnKuhc+0Cp/gm6Ycs
QsgwehZ4mIYf7gfKEHmq1wQguF4cX5YFjl/wbtsVHp9P7f7vAQfyGJFwnvfh7paNgr7NQvIeeSNA
uagg1UFT9aWx+1O1H8uFiWOubDJyI8CZIdBHFCp6P7qBAICP1uNBFwjjUmJkKMy5mWiuBHXpfguB
5YzrCew3tziCE6LW1HI9oQuQjZ7za5UcIQ/7W1epgs7AVekcakmJ08VRa0Yfz0le68vQkq6RDz7P
vkaQ6P5DXotLP/CXDtS40rwdaG4o5wTWeAMzf7CucFfDzTnf1nmcn+OMpIteLiCjF1PdZ5CrBgzR
bRGaBdhsAOzY1zipCGp61VH2oUn+M7TB495O+8wysc2QqcvHGhGyG854cxX7Erg7t+Ya61bBjBRg
znzNnz9TIdqAVxLM7VZRSJ1Ip74GDVaCCvm6126NXNiSPDGhtohhYuoP8o2TPVuhuaTI+mXVcEIM
hMRH6KMEm0dCfJOEGOSXJ630tJaEUjmFbT61mpSquWQ/6gGJlrzdbxEJWyJImpsirl0O98ZqtzUo
Or5z5Cm8NyQt4APfIA9SYzXVCF6ChIXlnZ4c++2xqVRyFqI+h23J1RxCDKpoybrfEAAk3+eTwH2/
ZWYGOK09QsjImzgk9ryAO7pH2dt+5MKYlSrQj+KEptq6Gdwg83gyW+Re0Yil5MUbdUkLZp4zNax8
swpmIuWl1O8hhVHrMphdgpbTNy3KeIyKWYbR3zYsnfopNYRZ3hY0YSbziMUCkV7YdxONX13Y/M1k
AyPnFzZGqiu8k+1ELO6N+w+k3ACunlcrNB1EWqagfno2YLMmp9VV5Mdaoary+YQduQq+bHMS7iLv
L1X3YyISwFfMqPTHC/NaIRPwDz0u2lvLrlsodgHtpKUSoTgAZZK0e4KkkRNgpOoORpBCrjeUYKyn
HUz9TvqOYFNH7gYG3WYtiXfLpDX3dwQ0oLFtcI6I20abURR1t2Es4h/hm0lqMhVHVwQUhThylOa7
5QVNXOukSbiP7wQfD9dyMX6hIE5yvuCyKRF5tJLh47hC3H6PkZtHQ40EZtTx+wBB8fesvtf6SsZe
21S03w9TrUEFBc4jzcBnV0wgNlwCXddSMvUoco+xPkB9DCMv0uV5R+aZFWe4UcfH4FWowd0bFw1C
WIeLX3z51NGQtX8kbh/gyA9weCfVJWOmwWc3OoCdS92jrjAHlnkjuGFko43vc40bOmVzWysE7449
nr/b2cIhf1UTvAFPz/3pA0sP8w4sxkWvusTim8tlOWWbBuLUnp3dLzwDKdGmyGMuusRoNgnp7zFc
ddM7b6GXxO+HzHylhYKUS4TDN+JS028eLxiRjL/zT+sPs7/FMR7uO2/sopxTDRvGsjp3O1z6nfv+
YtX8yyToYlg0icintq5ecmOKROsA+jKkrey8BbwrhDt9omcww1JLyeozHzyu3BvslsT70VcBYep7
O1uwk0HYa09CBPs4L50EyuYH5Xr+eHaFBgc6VUZT4y91eiry5YedfSbnG3SPCE70ffyePhabotya
/euf0RbrdpDFS2GhN5nW6Y40/JdL3kZhObiekpJXHD+V0WBS+b2ebbPnZrPBw/yF7iICI4ZHto5W
4Jx3an1pS3R6OzJ2kIl+Z66flewaJm99nVIc7Hsnvjt6q+NfWR2BkXJT3uMb0X04gEeP8nYyr4/+
X29kYf5kdNKe2c41ZJXGNCX49SRNCUSqX3xjixi63GZFLoiNFD03XXvqTBRCE1jQKd+KkaXzvzvP
N7E/vupfrthpaLFygqWpjo1xo3cef9GyTbvLtDGD1pBtYv/bm3dSyxuSqaP7g0d+e3Bx4rFRiQuQ
f1pkMRke2ftIK2C0hIQwEhTGfZOCPkDFqm5u2KvM3fmAk9C3P/hqGVA+zacPyKTgSmqILaKr57no
TeBB+JBjH1451mnxjLnOFL0jVjGBXYu1fc64VA3zL2OK495Ihik2Bc/8OjpoKU7JypomnB3zMA1X
0atkcoNmUfdDFjcpygGhY4nP79SNPznzDjIuj6i1jXKsGmd6LfIES1HhgJ8Uh5Yu0/MnxF1lB4Fq
/GcsbqOu6AhqdYQ6Qyhvj3U7G1s3TP3c8cQCmHoHv5u86hLwb9c90g06kl1QN5sJ5VgaCn3vwkXG
m+FuQrbq63MVouVtsGg0bebX02GTZSeoDvLod0EPGB2k3EBoQGD2n9EnoxcR2b12Vnjzhpm0rkpJ
7URL6uLP3pBlHyAQIevSK+W2mow5+gRwejeZ6Fd5r5FiOPr06xBO5oi5W1lv1ulJxZLGBX+jyy2e
fPivNt9gYrCjuPApbX00jPZEGOtr9j2QN2To9VCVEmsU+OSLHYWbIgB+PBI2W34ApRMiZeTHHGxs
QKdajzrjpq5v5KpVym64UgrDbrF+h2XzaVTvFCO7Gr0XdpkcX8ySY1auBTmZZ/joPf+qowdM9PqH
yT8ZaRH67Sc4Hh08tXUYKsL3WPygLNMSRIP21fzYZR8wz6ZZw3oG0T7tJtJYwJDHhFDVtM8zzLZ8
NK+N6gEj5RBo7hrIk4zN2eDzWmz/+4lEhFCr0isUzj7Brc9g84g2zOfCVLyI18vakot5cnv1toEB
RZ7sPmYAy6w2GeBU0BHcHMFK0E1kYXumMxtkQX1/B+vLVWo+R7lNmiWLGKvegzMfrv0srTCJxPPB
y5gW2h3Bbt3/QSjeavNJjrlSZn3DLJrhX1Zhkgn+uA/NpcLkmcjDxOF/b6ehCMXrSDgdYKKAmDhp
YropWn/15mm3klOj9W/yTHG8rRXiX85S1VEmshOQOnCjcF5sUhsrBwz7BGioaX+67HjVpr1q9yoz
0tLlGkMUXQX5SKfAHyt+dsDPTbeoRE4yeXg1hY2ZlTvh9ZCiauaAGJzRjnZDmU91iWfDemcywrmf
0Wwg9ktAvbqCwjkW6Tk/EnSLryod5a5s1WFgYWLciEg/4w2x+goGIKfJmfQm0wV6mUqszUAYsQQk
buhRtybnq9KG2VBKFunsIY80xs3QbZZbAwGFEHxP4D+CcP73LZp/iAx6XYiTO+jVhowFaliuIoaG
HjjZwNbd+dRwtDaoukfsGhrL+UIeTjRxKBsub47DcxCiiSZIqBOSgPASbLR8KtRXLb8Jc93qJ77g
K6Bgh3Z9ZyH/72arjOqZF5VFsTows8oJPr3uVmfhwELgUCUV/kkvtwBJY6Ns9gP5yNI/Jd01ZFJo
QZWWksisohHmsH+T47AbUBBWXxvdYz+r6bINQTaMdukkVv+K8tggVNqZzmgmPGGtvohml2vWUubv
v747w32omzHXRHWTTaUp2sXVKUUEzdpT7sMT1yZ7S8eK27CC3cxFCkPhUrDYGkmcc1H9coWcHlMA
Si6aScb99xmiptoNHbqIdAF2MOANOzJPp124+WPPE7lnUgtIRFROXmlyNVp8jg6rYOAlYiu7OK9K
8OGRQzGrWBkCc4tJk+ItYeINHxzzKXZZmQ5qMqaxVBOWizXEmmkH1sxnpLtgw6UmRBFHsN8mS7TF
plo5wk7ahM/ZH2KGaPtWw/gYtRuLG8yRo2WpUhO8Wv+jP/a1WXjPHAV6/kGTwfJtEtp3M2YTEc27
0s9kYR9mNppnoVaweT9rTJ6JKSV8OHn5bdpDL5yFXZCABJR/MSpSsnNEYmE8K16FysEJhYdWwkth
bMMMzcW/meEXNXfRHprREvJltr/tpkqrfoJfCMIoSLLDRvyy5jxtAdupA2zYiHe83IKNJazXJsHn
RXdE/ToKWSUPqy7IB7ACwnzddEpUYtWHGnvZSK9WNpbPL2M8yUUYjlhujtkl+r/oVMo+N1/ECEwn
uC0iNTcSAeE4QzQCN0Q1D5VYNlIkfe6yQj3vZhKGyxAMar34WiD2v1p9Q/XDlFYjXWoJWr9rHYum
49nGiDCbeOVJY67pTxcSJ08RyKatvggXdAEDeYbxchVRmrqo07NJnyjmXBpwXU7onNxWWuDIv460
b3YDlwylfyz3jZp8/mU/WMbel1EBjJ3SR0xbFpk4aRXb/dPcgIe/QWZ1k+cC9uqMSFLJMD1WZZak
AK8Q+6b4VZKF1qJ9+pCeGXtp8j76U9WvMzPksbLu+tX9k6mNHb+dOC27yzdzikMqyF4yxx7a27uK
jo5aBgXsd+PmJNXNzwC27TVVKQOouy9TCNNk0fRalPIi4WV9JhVWv/QKkJchDYaZ8EOdNoGn/el1
G5PhVfBoutAaBhVL863K1NbZlgR/TzgStJVZOSjPPKG9NPTV7Bw5/LP5uiPTqXCZkSDZ959QJ0pL
57dirs91eS+Qro63n0QWnMwLSCZZRPY9rEbnjjP/kZkDoyZLC3CXOcozVh2QtarV4yF1EM1QlonB
cQRl3jwQblR7Wm6GH54hXLauxPkY4ylGvRjvDLquYYIr9AroxJJ1fFBvY+kp72Y1Ku2NoXHm1JIP
fvTWMqrVFH5L1kVzIiVhK6JGZ8ywTUdVmWDzCuqTIrWLNsT//A3Z2noGGOUe0cJKsK+MWJCItRrG
9sSxDgOutuhcSX3GkTGPcMMeYVqPuSCfLF5pB39stcQFWY5QgDpIX5HqiRa35lPoi5tyMR7X+sKu
7hXMnOMleZbmSD/yHWYICuKboql+qOoi9qJtz12X9QQiNRtAOkFbI8MLfe0HDy4t97fToOnp3vUN
7tYiBK/g0imOADiEV6DpL4O+xTI31X2MjceEc9TVE0SHuyOUZzHaya2acULTps7qpIvcqpL9wpsy
XXylzR0q12YB9Yt2DWVsW6hFhgy0V24p99OV7tE0e370MnToXcpnKnQPbF0SdLZhyfXrtotb/nPj
F6ydFxwZIjCXQJE/mIovehBPXDjvizCXY4RJr0WveznGyqnJm1qgxQZHpUEKCFZEIRRzES0ACUt2
gqduNW7IOOxTCKcohrXx2sS4tkNKnn/lj+ha+XzAcUdWCV2nifm2SOGhhpMLiJQKPlyNx+Y5SDkK
/eOO+YbnN5bg3sdxgEb73olTlwqCj4Ra1MiKn60ZBOjvHa+l2151IXOPpFY1GnpPzlIfYhQ+mhP4
843B1uhrtx0Anvaupbdq4/wT3cKSElbnBz1Hh8M0DOkrR0OEPE9yja4wxBxwnIXkQKngv8KP/LpK
VOyEwcQAmaqnyskLw8WN6EXcDKl0Z5UqcX7dcBwmcA8emJTtrVHh1UhclCkznilzAF/KDe3yBRJG
P6hVaSbW+51YRPfg9OI3AWGThWWQHVl0pfpi4YxNH4t6JGHqQZLBpuR01BJ150FNPtATOQDZZMt6
GOfL9m2p0RJzP7wgVziQndzdYWomTQXrDtDhdu1CdRPhSLEFq/tkmBZiqRqUYIH09XxcgmzxrkdD
RCL0SXI+SiToD3Fwa37G9QGXKDlsMjn8WcQqux2txpt3eWXVjxcZj+xCGK5AhtGsIj7UxNd1rS4F
6tLuwswd1n/Kl7SgITbF2qtPeWbAkLxq1Sm9xKYD30bgfM3lhiIZ907PE6CRwNPmrRKMIHUhrXdK
W7vn3ag2RHl6Jb4I1/eH88lH9TC/nHdHJ77IHmGCSBP4oU/9K+0yVR5CjmPI6i9LbPNMwdB1mqFQ
F7AFjsJEG9VAWUvciCT4bM5F21vingiJcfr2HgLcc9/Uu7pkFd/Dyk7CZdptsswdtwt1isAqjQJI
epLR92BNsBrj6IXF5jGFANSt5vi+OfGXU538TWiPiBzNj7Ov18lINIjTWwhno2JbbMbTjTKZnCps
FhaUVXogwITk48GhzPOrMsGsjdkQct7FyAkkUHeDroPBXdCVQNEIDe13P3i3HQ/r8Xh7GWf7UgqD
XYi+AEUXhcqYjkr+noziWkQKhVfa7QK1A18lH3hqubikqEBUzjWjwcTJfOObVzd+X243tdaX6A5p
HJ71YBPQGg0BNsZ35OKYKq7fOrCI4737aMSao977S7niaaYiiA/XFMv293OrnbI2+y5l/KW+Vqzc
SrrkKCzoT+c5+G73qIkOE7Vz/lpdAs2HFk6aPFt8AiTXfu7E6CTKXpyC5mtFjcish4hxG/kmIXOn
0CxyJtwBpwR9LiHLu3McSFXHFjG/8Oo9YZfdEJY4tNZtmbWEhI3O9weIm6SD4rDc6F3/VYW4Si+w
fhkBenIAzSM0zlmsrbVvA/BJb749T0LoFLhHgHXLIGKmmnhGvScf5eixF8KYDBMvvS+S53TVRlgC
eHWo5QrKQp9laKK99N34v2jIHFdb2LnoyqlYhPlC+3YQUaRlGOK14R6fkekgiBPzD477mSjRy2y8
8BaLpJ07oTy2MJsa4GoFIBH1ZkSYTUo7H9uuprfck0elp4v3vwLRG9FKiz1rAWtUwemqjHe6NCWg
tkxwLJ74XPFuGYAfuZHa+sgJZcYMMqOnE22uxbuxPd+dsX7ib9lFBpDqtiazmN5q5A0qErKHtkRX
fs6hFMhzylykYxI5/FCzH0/XCG2WUlulbycOSDj785zW4jkwBeubpV8Y6dvBzONp8ZrrBqJhChYL
5u7nUt0MVdJxnbquuv5LAVpNzh9EWQLRSCFOMUHDNHGOSqV7ReTo2OoBST7VsC16EVVI7fmZfztc
Qf5vbtKZj18HLlhqrAT7bcqlXpjzgaRj1PDML63Wju2vHUuT7QRi5zo+CBdkaDTZ5WyZBFYWSnoQ
phebBukxTX/T3BWwsCHp7EsO3s0M2ZHXMFC/QTuhqD/lbgCIbsygSIQmJZvGESTmlCKNwSTLhn2d
+cD07dO5MnATnmxxOR1nCkbM580sb0g8G/s2f5Td1UdlqhqQxyG0RS/CNowpywU9nWbjyCiIfih5
XXf9U+wz3WI7pv9Q+yMyQx8OUj5X3bVvZ4E5qNkjBdqD5ztwJbNS37LqOcXm0pRvaa63dWQ12R/+
+WQXmP5qfXeW4vrIKKYF0OyaGn5B2g6rytxtppbHgizOGl+hNU8txLfDFykhVMFxgWJpB5jpZ2GS
bA/QBEKxHavfpzUiuLW52RLOiNk49Y5Dsk8ZH5OpSAW3BiMAty10Af1G954z/2VTtAQtTZul5PBw
5WhGuQekdlcNFouC9iQlbRBhyOp0D8j83quVIMp0rlcsFRW6TrEfjX7Z9q4gco27mC/KzKvrtkR5
Q2gCi7p/CBTYKL1MOopIbM6qs6gZlEd5KitJXz8bwSKmUhoT80OeSCNOeukWHhdfZvIhdUUkBIZK
1uqLABMTje3dcLY28ZWncS9tWX8k+7PYaylfSLe+HR3O1G2FF/hIIOVub6ZgDo7JzQ0Pj1Nrrxna
0icFn+rLrUEM87UA+0fYFl4SA9gl3rr8QYyCeMDCQgzJcN4Rsp9ZEgSekH0308GJc+D13oNHl+Fp
YlEBdAlJXEcNP0iFvKg4QPZXyLAFOjPNG9pvu98FZIs5vRGGw4UVwUsmAZMgQIT3o5hEzWSKJy9D
MobCinq+VJHS3XwPz78gSXauybX1FTo0fW7h41gIgaGO7uOeGdVdwR11yzxeYfs2FYtvl07dYgvx
nQVm3O7DGJf+D9Q2lCA6UhAEk72QKdbnepTtaYvMwJmJbp7bATKl8+hZuMHzHfiZKnc/T6ADnxJd
IUUWNSU3UfQJQm2uQ64oGJBmZi1Jlx3YbKgQNoj3wYLBe94cFDazBfuEfu3mjTsoUtv2VwFGWt+B
o8/OwF9i8DV5LagcLwmONYmnjfmipZoiq2/0i1sUaaKxvd5syWqWm/B0g4V4q+XtqqTf/2FlrHDy
UWTTDG3Ngxl1CIA1q7aV80gWwmBzi3mIGZ9RdIGGfhSc8F5hAzRE+Mk1BdJyQVamGB9bYB0po206
yoxF9pM8E3kn9Y/Z/RMGEcz5rhkCt5+UdSxsn3yu+t+xDjc7txG3FMCBCrPBpBMJpTrsXbvIeWma
AvDI12IQ8nF4jn9HQYx1VF3PT3BHUBpvNFCOQF5AVXqYwjKajMfmazrodqAQ7ynZLwKjb+G3wxMY
JGb0JyLdLRZw6U12QUoY5UYjKX0nUqooew+IAahKU4K2MHIsyUQMupw2wPpsWdTEkmlgZpHFnA4D
w6cKgt8ImMbkYCLbuRESk+x8aslJfu5Se3UKeBNhZPj5gQCT/bim598VBIB2V541ijCJnr3mTdT0
8UHlZ4ulfapNwIzRI0tUv69GZpSoa5MQtwi5HaIfWKimHNxH2622paeYkeqKgDPd38fw7w+WSAWW
lfuICHm2uHx40EeuBZ8YazqgKjjM9GdG689GJcWS73BrRdtEEZp35Sc+6s/ZSeGqC5Em7aPSkIWG
3Uf6SBrwAzKKo5HQ6H8r+H1FSzUIjYkrpRTpVuTyTXqQofSSiDooHgDzQAj4/HPrvoqO1+O4vjO2
qcrKCEOgBb78jQaA/y0zjSwYu+CF1tUc2slGGFtd7FvujWh2oO1xXxv5D2v1jcyW9WbaDufm39IU
adHCoV+crp9Dl99RQlhdy/LjyQuXOjuazBHzq6sLZad+RqiDViIlPxpXU1c/QYXurL1v65/Uo8qT
AjLoXYOc86BHm+0nZF2m3FLV3y9+A6TRRcT0xV563ESQQZ+snMlIW6Mv/8QHe5ULQtnGfr21T08f
qqIIfFZblsqOAiM3EqO/2dO4zzCzpuUdWIYxv/h69CyKftST6pijC/e0eKozyFVF/iWw9yYlL++Z
5Jx2UmIzov7/2Cix8Nwk7CxDx4kWJCRropXNb5PPxfn4G7vsd8YSTB95Cq8bNo1sfsmoqyrcDvp8
bm+0RF7ytZYGEb3Jf4U+lcI8kuguV9Hh4cDDXp0azlm9YoPObvzDbfs5UW9SRKLUagwoONTOlDot
cjeBTD1cuCMntwZdUAKkBLDFfYZar3FAJ9HTdHbZC3ajZXG2sntTWbXDs3opPDR6XhPjfhXUn/Q2
zBq9niALlWlmwv8SQdlqPi8+qveh/2zdB+tCmYBivryq9xlSz+JfKv62xr3nfW+VpAfwc/arr7OI
ZIxrtQVPlS53KGwPrhCas7DRDFpEy6mrKAB5Cpg4sVePKzmR0BAiTjxxMtWb8vSuMsE/3bxVjv7T
yE/T0o6mHWRMko/E2v7JFvWXfiZW4CRCQo+zkyPKtY5eVdW6XsruRlHyC3KWVZn1CigSn+fQ898Y
qytkvVj3pbXdG3XFT6pfRdW3N0bnGOQL+7J1AQfwL3EqzYM7Vmws6no4AxT/EEG22lLd83lS0ZKv
yO/xuiw5mD4IFAEI5hGwEY1PA0o4oFvcSn+2EqPIY9u9ir7z9AJT5dPE476m9fWNU1zJGijFx1zV
kXVgU8RkLal7oguf83f0DCas4EAQuQL+FmnP2F5rzJraMeErrDe9Qqz90ySKcj3WG5EAcCx2avPg
qBKXxrzYjjk6ZxY//deftPdMwLa8kinbtbR+HlV5drxvHBoWI7pBfWWKKmJcoUJTJoSyFESfZyJp
fr38oTKE1mokAeEk931GWmDNLpFEfoO1XioEKnUPtT/QeZbliIVQsH4lLbDST2bsT7hq2ohBsBIO
DrCbY60C2Y9UkGDAB4CllxbPNlZNjLQ3GFT8UXoAo6fENqf4wmroTWQdn/KdWs7z+zc6jm+vi12a
K7Fb6GFsCEoJZ0svjEgu9vzXzT8rZRxSPKVas3ohIXHFZKGMXsSIbno7HLmQtfwTRgHyOCCWfcjG
ZxqI+gNsTK1+Iue0hedM70DXzSqFSTS8kCR3JGSCrl2OSUqkp4zbU2QiVDfTDb6vklfklQTsCKgH
Cm36ubooJRp35YeAY9T3QFLDgusPrEzm+7GYxY0bhx+Q6Vcg4RjIpHLQ45Z8L6+vtLV1ehH8+PBw
G8V+MbupP+T4KV0IxnQfAHYEyC6gieVigVfZjeRlSG2ZPNyjHwWs6MID8XuDvO+QXvvrVxyYJdbU
iYcFBUm3U/U8Tbo4oXOvkMAPYAwYS/99CFIWRWcoZaeVpyw2lVToGss4wZkNgU6uBg8qAmSzomui
EAcb4pQsX9eI7m3lZriNpcNj29EkeQPegKbQa6aqUX1mhJ3cenft/Gxy5oZ9aSs6HlvLNWQebpet
JlKzqtGBiXLsbkNX8z1R+vfORIX7yE6racjL6iC/tQq+lJmpAC+5JlWrxaslMxxatF5zKDTkLTjK
c7F8Iogb7XHmB+aCisVj59JGytesI2ZxZNSMFlC3W9H4dfMYOe42FUehFvs8GpE0Lej0b6AouB7R
Qmx/URR8Kr7b7S1hl/oim9A10gDqdm0nArwFCnnzB3LmpE6EQXe+pn/vziFY/GxMpflj0jQpAClR
3JR2E2zLq+jbFhs+sAKmMWCLChyZ3cqJFJMyRx503tCcAGZWD4oFsyd1i7DMO1z7h7Grg2VElEAf
U8gc8upXefyKk8hp9FsfN9MstXVf8gFUuz3ClTh8qkvAL6UufEjxdR/+Y03opWCbyTg1wmuxT8Az
lhaLe5eSMCfPudTFFpwwQ7loVnx6yQsZCLmiTTfefALD+3/6Ad7d9X/KUdOM3rHUSgmvdj4Xn/4A
zibyvRMcGtGHoR7qurJf63hvno9qbVjmLoIMHKYeBVx3/NdVYj4luhEsC27wZyhLq3Zk8JFxhx5w
tycLIM3PY1phWQdrjZ7uRodzkmiQlAZe5fzi0I9fPunqpYxA2jGq7CF+ufyU1lkTlWgZvmtHXA8z
rfjGV943vDKLCk2lexXBmTSxzBEF1qYcY1ONL0yYFFyVw3UU+1w7+ku+OSEilBgZSS6TOBDXNrbp
K5y21DACMbJ1xPYpeyVYvtwMzcTJI3jneZMpPk9efcjbnyRftSZxFDI3p1f5nFAymngzkt/DK2S+
W/txzOBb6k7K3vlIOP2A/lb3tGrynNQa5t5JL0z/eNjF1PvwMHpz+BILViAF6ch2V55tNMYLt2PR
6LFQM4HD8I/4uDN9+Mvfdw7KCiIBGV+OiXxX9hjiVnTap1o9sCi8tnuLYz8l8S7oeS1MnPREImzd
He3HF+5WrFZInrUUNMRra8PnJanM9Ytje5vIXqnUcwB1rJu0nXqiw1JPgDqFqtCJGE9y91wfenDS
/0sYMSxspQGiRcqHurzkxv1Xc/+YXjSbxPkkEEJq7K+KzRSSAVchX75GRFCB7XNn1oATritcpM3i
6B5LDin7FfxWVO4olkZvleJtCEcli/F21ptNScJCwpLFRG5RpyG00/1FPuCMyO0okAhwRIOD+wIk
snfszuRg4HptAVnrc/Qnf5OnWz1DRM+gqjHzTYjBhVJa1905c9Nz6TSnXH53blSJb7hH43lfMjtX
Qdp9Tf9eq9L+xi7wSvq/3vHHfjCRTqJ+6mK84pFWlxzynGuiLtNvEA+z/0PM3uiW1xqkNv8VVpOl
gNwUp+cfdnZzljsNV/tc0fc6cJ5ztjpuGH1XqD4CJiItMvy8c33mKMye60ida1gp2+zzAZFRIVNZ
ECy2U5Cc6q5V7et4PFnJF8EUm/q9pQY1I7+SL9F8fjNfDfKCjx7uFNay774jqdgSoWSLyN7UzVzm
kVtTMhkFE9AknXLYu9LDyHNBmymZDWuU+dqBln1oHnIVjnojVoKqSC2V5j+l7Y6iZ+CXaJPaHOwd
9zSk+tB0oTfSDXSVrzUUOSx9wRFK49z8RGB2toft7HKV0jwAv3cybBCW4qSdnft82kup7QhcOyo9
Oj/sBRiiLknVGc9NQK0CfnGecllc+VPxWOGjb/rIalGLvlrNV8hAEm8xuW8XNjhYcIUwskb2TBru
IIjnjYUUSSdz65XomDp9nax/z2Li9QyKvVfXuuoms/IunWlvw6DL8pUh1DP9a8ls4b5BhVVA31Aa
4ndJzNT+jGQTLUpmkLZR9Y3kc5+3SB+DnKOhXTdtHzGrJ2yzuVbhhkycGggWrYlK4qkca2MOJ+Rr
keBYaoHbb5nXu2Dw7UmvUwuwJudpf2KiwGGGLtPn3Bi6VfCVyzZ3rPD9ojKzzOa4zutiuhUash7S
rsx69432c8Z4WoxwVYzKZy46f3P07bNUBi2Swgd+lTBh3Wd8Lc/dCeGhaknxqSEcmtF14/tdKLK0
0j+aAoXXH63JhU3djlyfyitxI/VWGw6kNuP7/Q3hp5PNMaIU9JaLDoufbUP3TDnhs5HpAv+RZth4
1u2gHV/YyDtkQJBcUw8790R5HayF+/MANPJ3g29Dwho2vUdXGqQIwWKuRSXVTaNf+1J0JuIgOhFq
NPIlvgMJc81Q+0SvL49K05W3pThKX0Lu+WBs/68tAhMkvWSs02mbXCuVF2//qbbbg1+IfsZvlgw4
st4zuKkwlgsC4DgIbEeipm/UZ7FupR25k7J5RstokAL7Sn/tYoGI3vpilAXfzFueJEFI7Evg4UpQ
+qYmQYNpMG4ZaRY7KQo+OuF+JA/UN2D1vE9VUJYqtxF4wq+kLVWxxAun0OamDe5EIFofob0gDpsu
Peb5aD/E8Kp2/lnltJ8+xoM3HrVLnUbsFVVSmkaXgGX742H9LbnprRq/McCZ6FvTImkGL4elJbza
pGKci6NtdbLvyLXAdcZiBmbo1eULKorAikrsYZppinzj9sr54T7mDWcnx6yoM3UYwJWdJVvpSdkt
I8YkL5jn8GRMAORnY28WDqVwlwlkyR9RV1Tnz3u4HBEJZpGoGRlnl2YZmxC/6gsbJUev6yKUJsak
QRg2Csj6HxaTXGd/l1ywtGgPbxJNManvFz2vU1eYgZj8EsKlzqof/uFrzcjBss0JgZc7bOidpRVu
nt4DOE/IaZ9RY8vPP38aNuqvEHeC0V6VIXGIYbyaj/gFP2HjvG5XBIVmpysCobWRGDY9y9rE9TXn
lH7+J/+T9Cu1632bk9qvKcA9QDJKxhijNxJjWJ5Mhy5Su9Uq7IUm0tSfR2mpIk7JmZTXRZ09/1B9
73hRgSSMT7h6zIlXf87twIBFElt5Atx3AwB2Y8WsQDYVymgPv0Hm5ycJtcaLnWA8lgOCjxS3pWV4
j0iSzVcLyimQBnyBz5IEkO7bqWPui9uBJwj13dUOFKeflgJza0Yw9aI1jsNaPCzbTWOg96L3muF1
7j8A79H75xnCoSnznrKVPKkcnwvEncKxQaVOWDpDRQkBckTK3CDPoij+fS6+Uh4pWap+D98UdylG
ZHxQt/2GIsxVKBCAx9s6WY+MJ92Pwvo/dzL6nV/uZQm8Ws6LCTSjPpoXQERwurWynMvrlDJNml5d
EtEPbCloG32ISIl/rQnNEyTIbsoIuacO+y252WC7zJuR0DswMJJf0uXhUiF0Xj729tw3rmmbBoGI
D8xlZybTsdBh4Y5UMvdzsljv+d87dR92gb5b1KJKGhkrk9yuZtC8zVUaFlNu/H4lbbxSR9q1ZHhY
yktUb58FDppw5Ji7NUZmZs06izuFf9WplwCGqqF5jmUH/bzZBWw1//h8uktEHMOoFenjvqCPDP9A
mrPFbQRSdfhagc0Q/bV2C/USUQKyCmMJCQMQ/MawDevTcccgY8NqFZRwcIc2uscjnNIWujKQL3p4
xRoxfLhTv72OWOS9GR2lngEAqOy0wHsR2M+Ek1lGU8G6jV7MlzlV/JZmJN4ybbyKxkf2Ea5eG/a5
h2yVWCuZePMXlsfNNAt4jSQa6AxbwmF1ezJpSdssG4DrK4oytBXAhntL2+aK3jhERLZBK66TmOG1
TCe1cVaH0f2jF4NY+5UQ47jzP39CleM0QxdkZF0QUG0+5JtU3okU33jZB6EbSh1enrR4U76lH/Ra
OcMXNon4xu/ckqG1Cj110GzzBIkMCDglPRT4DBxgWzhU20ym2JBynSgMC/5XamtklaoB/Rlw3Cfk
18gC9mJMUBEJnx0CLyAvRC8QBiBKidiCNZhi38rSm5BOve4EgNiuTndeGJ/AiOdjg+JDCTSKRRuA
vrCqx2/RtzBAo/7mUxwdBeL66TM2JJe33cJpKspKQfsbCIYxerfaLzZO4ZbONDUTa2KcOFRXemmF
yIyMc8G2YmilpyaKrYsjT8sdQxujeXNpLgnAxE5LVdECxCimUdomkhLv9inBWzhrXGvieq1Q4Ysn
vEztBohntGl4wfzel9cB7dFpTq9ZPv+/qVlsE/Nul36XjL26KMqcQkLuclir+ZwFSR2/B9NBSeZQ
M5eqOOZNuG1GrjJT388ienzIIlBCC5E7Ux/RTSgixQUuy2kAQB+Y4/vrDD0sO3nBDv90Ou0K1ald
nWsxJVISilwjGFpWf5fxx9uAqY99cRcylAbW65fkMF2Wbr5oaYwZCOgT/U/7YjZHUCaPRkENj1zx
HiLggqfNzfczfg3PNQABFaQqAe+1tl1cG+Udrx0HWYB3HHr4gjceYdNMjm/kyb6OkF8vqxWzxTV0
lD6dlpDTl+taOj7Iqrj2YqlSMyITzqSKZICvjt5dsHvegb5r5YVPU82yUoicO1MPU5yI01uCeZIE
vcfsqgH74ioTT/RBIgzbcY8nTXLr0WI2x5yK5fdQvojwLVKVD4wPFtwPlT3fMnBeuvdzQ/Qv8UUH
jsPyjlNYUKuU4Bq91tkZdKnTFpQG/Cb8GRlay3Jgg94LwbOZOqPcrA9OUQnx/ZLY1xvAgmJ/yOLh
yeu+NvARFsJFE0ERgWRhJkqtzDpg2MctkrQFxmT2BGRL8/sbeNlmYWpqiczswntM3QEYWyhTMnjv
3tIxtaMVvhT7dnHTbHG82ylfMFLu9pkJTFOR4ORlCgT22E3jvp9d1toEpnggDe07TH6KKWrOhw9t
S7e9U8m/WkyEiNdyHUwV1zJ2H/mWMrXFSsUgz2/EicNlq2l5udxg0FbHbFNVgHaIinMj3mawhipg
3yEOoFL770a88uZiQ8V2TOcdFBcTgY2snuoCJX9tj09TmV1tW4koFYAzfw+K0mh9DiPpW/Y9ECym
gHaSxK4J+ayQ2Tbtcj3bDq334uBVqeXfurkmhRSWQwBK7Vx8Zb73FDjMscV89Hl/ZGNpyJqTrgUV
cJ8Ej3RTWDShk9kQgtdtBnLQ5r+sQbrkC1hQDgYzmhe+gi/uJBorphRR3q/Uopub1WdfvHdBg7yz
hWx/5NJG+rDun7varfc/27uMeUb8eLH+j9mZ2LCvULRWsVQA7C2273PaKwCHtAfzduWbONK9m0ia
gb9BeDMqqvCfHQUmKlqy+NeZLm+AgMBz/Ot4iIymN5gscPjgkBcEh4S87KBL7qkwDokpbHijd2uD
VMY4+s1zjjiPMWIw2VeWOLlTjJuMDyO+tfOi8k4vvv4eDoasIWJIQJ+CpyLDGvql2QbLnmb4EVCX
4cCTzrBKE9DZ6Y0nTjrAgQpBhSmBd25tMzJzGplY2AkP8muUD0UPsu+Atk+HtlYjCWna0sWuGxGL
ID2vOcmvneIzL5EeTyH04PqFXQKP8MIRo46fAFx2QeQZAIpfiJQ+hyPOZ/ZsOwJMGQxme/B4DwHa
j2CAqrYYnhBK7mVrzEnEywnXnT7noFHLEiOH8RXsaPFV/7S7j5pn7A4SATYXkebVLCeNINAuKKa8
MNF8EwhKpoLo++wS/IdwHpEaB8NzK7HvGKGjUMGRwhg8+I5ktnsd51IgB2iFZFbDaH5D5mwPaeUA
65jr1MQuIs8yD4zXJzdq3aGd5YPN8NE6DsHIepDybnxsfl2Q0UsI5mYmSv37HTDuNaYUT/OcrVzb
mmqY/GaYfw5loswVa3piwJB0gkOwfS6mEwfQpIikxTNjU4dgrI7HNHWyV3UKpnBv+fyfmaLPog1j
fg4wz5hHiCKLUuyV1gvv6GW5ek3Q/Kr0mnhslhpd3Jw/9rbSB6AuQFmd8YT5OIIMEm2erRSgfY53
+s14mKPyzXMv5Cj2ZLkW14a2ID7BEey3aexKN6tqhiD6LfJ5EXbawK3Rg3bO9+CbXt7R71yMIpNa
5jDeX6HJb/MOLf7qvFrLAmimzcGZWULoKtTx3Qb3fejG4s8nkesduHLGZN/AhJAY87XUn82EFCZ/
IQC3BhoXGDqCgsIz0I3VnKVds2QNrBoEMHDqVocHOAg8vgfv6nBxax51QRWU0RueH0VhFmh2uH1Y
Ay6yZgb7ApyDOghrRDFKi6Pb4hvtzVBxZr4U9fe9TLx3j102/qbs5lw6D2ZJCrfW/MtQQa3swe/5
GCwmaQffCbomyGF4UuHrY+tOknthP3ydguQUJjIzd2Hh0MbBb/y/Zi1sIe60ygpR/7OYnhJfdRGW
SIN1x/8vsWLWZwCW/+UTtT1vNbLNRkFillZzgcZHde7gYiHXA+eOxQxFUPPhONrWB2erVF7y18D+
kL5oopcncAjVq+25Q1yE2uWPFc/sv8wXXlnWPfYdmeyHx5CGFlac2IUEBuaLK3EZimZMeCZqPNk8
BJUzZZLOB+G8b4Zxo05vMvfkZdObgwpRfxiugH/j30YJvrlWyYVkWkL7nmBPqk8l1h2DDbaiTGop
PKOFzGqzGaG1onkyg+J40o4/DIN7gWOvQuct7kQWZXm8hOuXSUfAy2sgrPPw/S/Tn8l0VPE1nLIQ
nnQ5896vqcfzgmPr3i91rHDSp0KN/5EmpG6PgcAee8zvUIIO7XIOUcCYqSbh3uzR/GEYqR2/sF8F
s/GqsJD9GhPdndmmEwAIsnTTCqzVUpBj+UTf4tkL8SGoCSfv36ZIXgU+1h2604nAfVXc5BwKM3xi
55qcWpRNMS+4hq5uLpSHgVkO1xoPRTETqjxqTlSJbOzbr1qbKeZ1/55pw8YxVBa+oqZkopPM7zUV
8y5P5rjPn0AJ/QBnGes1XTCmgiHR9opauJUFtZi8h8t0fN1wt0kYByXSL1z8czP5Z6j29v9yr3Yt
eUFetyiVBGnJUHfI9j/vAvl2BddM8l3W1CYVKvPus1lE9q8lpz4q6A+X9Mky/DhM18SiXrCA5kG9
QrW+T+ImJx7cSPuXSnu7KZFQQ7nuvNfOqMduuMKt9eCFZN8lEl9v3sHTpAUMd3p3YLHA0YKZYet7
nBl58c0FkzHqDxYv+eWVEujtxWrs3X5L8RotGIoYktv4IHtU12r2A/ubHMyVawP1ZXHNqhsoHDCn
LtMuPQhRIRtSnHy0pAJOUJuadix0ocAc31xqZdONpDai+HhxRdJgvjjy8k0xal8uTJ/DNxZKJJBX
yEdZroAwF13hB4MDbDZDRPt3nqvsLgLOjWraMMBC8FvaM5gOOGf93whSxPhcnUHzseyqLaI/u+wt
H1n1ewsn+ZN0yFVwQ+2/vYH4s9YjnpJ1cf1Se8FOPp1F0PihjnJPQTnS50D2p4qDjhYbjnnda4Bq
zOtBqD4IPUdgJOK2gL9aneq5LhmzkF/gvjZntaS78Yi1hD4O2UBlba8RgNFDftoEBjpg3UnhowpY
mxy25ZnO9TyeWnjY58MYEEAnlwLuSCJIzHNDsYtYK3UGTOsXhZOK0RHvGVFEsIV5Q/YynnDiHIUA
Z8KoH2QvqUtYC8dtWPlBAM4zB4wkmB47UXrf38lYHwtC01h4GLL9kQavc5EklBk/96rLsumLYbhD
VyXY2rfRBI615ym8Za7Ji5SF+BWxJycb1SivhTnlAnvcsNrFrNI4eWizBLavFms4DflcITnDOL30
c15u5+FF7p+iKzv/ELAt0FZHB39wl83va/D6DzbxVGdjerSKuMpTv2ZyAdLbgLwV5CXPD4CPs6Aw
BWQextjear4HgQdG1Gm2xoUxkE3FvumBrCiTxVlNV/dQXLRlGHt1srdzanmzD35oosjaLmsaYdQB
4Nkil3NRAfXKyTmnXwV9q8NnXAbLTYcrm1twcf/42ZZgfRgMg1kGfh0+c4k1vKoRmks0VV/w4tGf
P5cwrf7/+YtfZjJpBz5yAaLw9iETHhpKFUB5qOj0JXhKwOLFAzp6hhB3rWFSoEXMupBT/9uoWKTk
hBUakm2jr5MgosXZS19VJ9ra+Nn9dHz2Wer0m3OXZl6tkHCCJCwQyStrt5TVMeAw63BlYLFAZ475
s1q3CDkfg3adPyOHa/pypVpGgkK86j8rc6pBZXto7JtwFV0JDAdN1qDdmZUS7npYLGhw2zAoYc/O
lt7muQyYyBEep0/rAI3jAeGb0YQ9e78a230SCwAhSlD3DvSNJ7pUXveWsIx6J6d8gdsCY5zGDXwT
Gb9rY48uc9LH9nsoq4cS+nqIwNpWvb0GfWdWy1a9P7mpr1qKAvAPOvM8PJPuLUTMXolPduZLFWKx
7YXRJZlBFunlxM7igx98ktJ6P/yclAZmJtZ+ZxLb2E+z3VvkoZ4sWnyZARE/xaMOd1OfyqWfS9UV
wqnt4YpRSs3rCMIrcjQHaXP6KkdRgJO4weqB8p2cmwc3Bc4ha7UjZ8cWj/GPsZC40eqy2R3zIAyU
X6X6eVOvVKLr+PFAb2Ckrn6gF7SLjwYftJiglY52f6LJRLUVhe+h0547BQE8Aeki9eJkReux75+7
Hd4uyfIDFYv82Q55tA8qqZoslsnch79cwC3SeJJ7KMDSN9ouAS11V4jNviuoGAmlatEiKcPiZmQk
46RyDZli211ituCS0dkOxOlRFMJb76ErM1l7LVyGnco0k0qjuocf+yLYYBFGA02+v+86n/eN2yp8
02kLafx8LHul3hNVD9n3Odsh7kttTMNz/5qDeLpnb/sDVKljbIrFOmc/O1eEvgL5PIri0HyVTXyu
h/KmgA8Xb/RaMXkGkEdqXnqMnBq/61yuD9OlbXakADltxBRbOE3A0cPHGwdZBLy4CHl8tmd6f6Ok
hrOC45L5PdAdbCSDHymbXUzUM+/Tks9u5ERp2uUw76j6BtR+8jCLrNfmTGCroYjnFOpZm1wNBWpZ
0NuDUnQ9b300WeBKMI+DHPRuLexEnCK8tq25WXjBO3YCqvu1vi8T3IOHygRa8WDt1lH2F7e8D+Jq
ubngJsu3m4LQusZBCKo9cxA71iOpeJyu12GihjxSvQbAKwLgULLADJbKdgnPmBi1UPYQQ5nDE+w3
NGummtdtm5PQBm46foxDQDoQNcXAqYljIkvso87P18X8B703baaoubF7p+J38XbAT4qAdtiK/7Ya
p5XNgrTzqYnuOr1P4sdG8/wRo4kMvHU+nXXUxn4SB4fjPv9vBn2YXQ+3S8pSdhqBcILZ2/I9PTYa
uU1xCxW2Qu07Jd78aw/kkRjykrS5er133LOEk6F2KFOo3Ct/y2h62x1/zErPe3gfcY2vtolmDMrC
G89tNXw7dEt8I5nGL3bjibKJK4/Oe2oLmnmpP7+E+nkNJEUTigEFbPRObglkg7gY4SlTYstvXyLa
tJ3wanCq809yFzIvfwfHR/0gut/D7JpHC0xehmpB2gPaNE6W7qXkT20AroLiZixOuV2wKL1WJ1v6
yJR14UsY6g9thv331o21jkghdV6ef374fuEoU1JNR2EZRWkQa9ks5h1NbncFUW3pfts6p6o+B8vX
Dc3WobuCWi9yJ4kx/dhCjYkRaRV5xqrxtNynBhMi4YWiu15vo2IqlNBs2e4PLvtwzRZSXA7a2MDi
QEvWETkomwl76Py1E8iyjWixNVOUpwDN5o2BNe5wpM2qUEl2dbZjdXRKcqXq5OfVQGMitP+HMMHO
K5qKjmPZDSr+aEAEzqVcpUQYJvwbiKqUe6a3V9rPrTaBM8TBNN+SR+00tbux0pyoBjYOgutAVe27
OTGOLJz+inxViot9i7zs6vQydLFyU9pTEDlVvT+TxfKWD/pRJVvIYBc97HzYaAzv3X4grk1jVN72
x6oCycgROR0FJ+45PAWN54dv4EfJ1KjrEXXp2VQ9MN3HSATKQH+8KxSU8XvZ2wDUhMZL1TvhMfpw
nvhiV5klVNdLgdFcXkfSiM8bhYqShb1pspzAImObvDwobrtg6bHHmH14DGr9HVFnuau/ymg3+PWW
rjHki2yxdzykx3DYOq2akVVuV9KDYhjsn7FAcVc7P1VJUZQ9VjnZEP9JUkNGgjwBp1dPpkdfmaGT
4N1ghrkirCY5w5m27Wro9jxBy1NpKAhdAPY0FtPWHB3X7emLGGS0Oa9bhRDvU5Yft1gXOepMuEzG
F/a+S3UkVmTzpEzs3QIZ7O6pZ1Je0XkG6Pi4su0qw+USgcQPuxvUEk167kx5jmW3fKU7xmA8ltd0
v39NCttWqnPiULe2ssH9yjRxZpCeAG+ZvH8/kLOEZYoRTvk93jKFjp+50zYLCSTirs0SypA4Su9S
W3WJHJQc1qqSlJWjaXE/idSz/It6OKUgw56yl5r5FRVpe8Gi/wL2Xv3SPWWxE0a/a2lg18lTlbxf
Eh264k4EIEWYpwc7w7ZeOv3niO4Aa7WPbL2tFtiFiZ4N+U7TIWFzrc6ua0MbzB/5/IDMsHfBApmf
9hbg777p1q3d/IOTgHxei1hd1W1zdH7z16Okewt+HgcRUmKXj7F/6zqwOje7Puy321ZNE5VWvoVR
R+pTCHUMXqqCtDpmHUSqd55jh2HuW1aue6EOnDYrR5QHeXAwMU0cN4P7XvACxNYPwd1XodKtYXx3
UxY3rKPJBixB1X1BtTcTSi6k1uv8IK6u0pLrdWyehbkRCWfuXbHGEoEc6Zp3UC5k4hVHFafBLaQx
IcMsjbPamAsaK6RiUwXslQwQ+a8kfRQAKKRBXA+gtUi0gzAaRUbWYMLwzBZys0ckmt1oFiJpbXyN
9xpOAM7gxWrzN7X/irENY9XALwcHnbNFYNVevV/qjmHIbYAAjcDuufaeA4vzxZ3E0XJUouKHv9vC
VyBWoPxWHI0kLuIoc+V6HKxmNq0C1YWEIzjZtIAvu/1FZTfaSAQElBi6axL4OkWEfHujPWROKiMD
IIadMFTX7lPKDY1gqMnjahopZFNNE80e1Q/oKLWmygejP5GonAGA6/xwWjDKzpAHsN76dCGn3yyV
QriZrWUAMG8ViPsIy378xh09izwhpRNPsL3b3oNry7PK+ulvQxOmwQgdG8NFYa12XqDehpwYOc4h
G15yCRd6iXy69lERg36Eowu0IAN2F2F3p4xxg+p71ntjnIGUzb6KyWZzPgCCsXr9OSFrRZvRur7b
EIXzXJACCncs9x3hnuAKEtSd+CHBTei76oFPWMsI9OsVetIkx0dIl72dSj05o3xbcSGsaRteFjCp
Zi4o+VMdr4Ih/cVHNfYWpYaqX8FjqlcTe/P3BrfD+WtOdTcqGgI/5lQZKJ+2+R2dd8Nt0x6yxk+O
UGj1CH7GcM6hR0OXx2Ey17JoJ9ZsRtxLX71JyJOslMw41cqrng3VWrkEdHoy0sMpRnc4pUWL976j
kvkNFEP/L3boSZ6qi6bfnYnrz5/bhUZtwP5QWmsUw+3FOUbA4i8BhETv1eh3m2tD4xCN1g8QALce
iRP3OgaUyBCgorw7++OzUoNkd9mQjv97jkHMiHys8MfjmwdEPsURFF74IlQ1GhIZdtbjDZnSdbJu
UO2x6rQ3qCn9bACOSPdyCpaPLtiKbaheftsUQv7FJ1tyw6iokUAiSjt2WJ7j9wLTNipDRZ22snWB
wTy7V3YJZZ3Ch4DJfyrJN4Uk1QRGgbcK6WvOrW0kQC5KfkqukQuafz3T0R80Y6voV1RyEeZLv2P4
gRTRMkBRCF+xFp1Eh20qax6WciaA8eGa2aPGHdO9rKnqdcqj/QIhcnjd+li+m4LsMAiUswFTSUZy
hHXz/bTKxyrMRXzzLtJh69FGuPUgm4z49Bo3flLz10tA9tjp9xS+ZP1HqqivdbB3EBzrMxwVLLez
MOpvtmr7HUjMp9CwNLGYO3fuocyg1Z82dpQZpuTcMG239h8RzUNtyQFMGVa7gQHFTZfPxngnfk5r
yb3tD2Lik6Fk1cYf78Z+G7sqpl/AeibZt7jAmSkCkMZDN9qHruYuYbJ/d5VESuh/MetcmRNCcIXL
AjILO0aGTOEMrjT0SIciWfMt1fk0ysR+41/AAumKnElOM1yEjDStz93XJxtg3svBRlKVTj1M5/94
/hZedp4CyczUrswJiAkvjMTXKIIUl8B3g7e0nDYbYZkBRJr+9D+Aq972BQmjQ+EhTj80wnVjgcog
q2jimH0j2bJbc4cSvDBgNySB1ZBgYOsu1jusjFFMbfoI60buApjT/wZyetPS4lD9mgrusMTtypK7
JDHI9K6dMVCEEP3ja4CJS6uIs9MaSCd5rhoo3zb6uyw9noYjtyS5p883Bmnh6xCIMUG33oBNENrU
748nVQ/ImdwiqusQjVCitjO7UpTuB45OvEpeyhMz9Wma9NZQkGcgmGjgvomiwP6MklfRG+6K1Pur
GYH89QrtuHRcoWDNNrtKtqpclgb8Fm2DUsn2zvjhxKoqM+vvkmHP26vMCHs5RYlWa8zrEMWlEhiQ
qU720hWcIIz15W/WyVm1cY9JDXBQ0ckPcYHsa4lEQLU16Z5Cvkb9KAucuEEr4Ze0ooqnPCSaUOON
wYQ5Wco7NGwpwv06JK2didgRs0CQdodQm0x1nVLO6gzW3S1nPWXXsyNe/e09oAjVfsvRdTRzbc7Q
pUG4dCiReQmrO1ZphwmxjLGiHsMWkDOEW9pbgxSqZPeRcrx62ERXWtEnBvwOQSOihpFD1CDsPTHh
I6w+Si03uwihx/b/sikkVlxJHZxgEgdLtLREwza12zA+EFUOPUySirbx8iNAO3aBZwTBnZLGRl9z
XI6wr+2FipvZWz5lg1ePJo0I/QrjGH4gTVQVF6Eem8pIzyWBOdv1WA/VGOiwuwYJwMLII05KrhJ7
Ws6+wakxfn1qzYZXCGVzA3pDuNsRlKOyqFZgH2xnWIbGBhKVtgdzDZYi/Xhx4nOLH5ZY8Ujg2l/r
mhRiKDQhmWVMMEmC4vn/twrB66bnlSrNW2fJazygkplFg1vmxdz4NAhjd4yWERqbHft5j4eurz80
nfmhYpSao38KMlaE0t1p/8nPzfquAIEC+BAM1iu3jL84Spp+ECkox8XnPZDO4NBNWImqz4+Bs6Vc
D2xtqhR8uzKweNGbtnAZFlYFnFbABxUhSkQaPWItawbLL3SvG6Y3AzCYGyN3Uqi/C27QuyNh/kjK
i1jt4fHo/n2pZx1h/mhttrsqeHGKFVMTtBPzA6JEj/i3R6sS3GR98rC+RdomwvkCIBUfvu6oHKFl
PXNitk6PC1VIHiHkBprG9S+UxCrmy3uZmZ8zkAW0f48QFgFYWiTEZiB7aFfGfirvh4BfAJUbrtfB
d4JWMMVNLVZptEFYF2Y1WEwQNzK00he/nXgSwzmkhLYQhlVpsy4HF5aiiYwV5S4z83iyDfajxsFt
xz2dxTT6hamgyKWxzSeAGMUpS+dSsA2HIC0u3VkkDTvUaQQsuyuXJaysajQMQFG7tWTvFwtAt+zE
gPZ0Qd8W40/UI6cvWK7TjA56y7YEu0/IXaa78g3L3XtxKUTRsG+34847ep00BLxk/5VdsAFkKmDd
EAtrsAjOsHbSHjLHLUdExrlNPFua+91+gYQlgCM4LZH32yNdv2WWEzJgzp4MZxxajYuoatjouNmk
5yO8jMEDMUMavMLIG09GUlBv+cn4p2+chsLAG4DM9KOaBaVYGgZopJewRO4cZP5UrmDsYHhD4Zso
zMM2ikTUx0t/h09bnXTJr7rEpI2TF1YvaXE0P3sEZ5NiEki06pLO66a/518R24imjJxzwn5nGMqT
n9cG7LAAd/chop5MqepoKgcf+GhvT6yrGDUsV/ILLbhzskcoPIRC0TPVh4Iwz3EPnQgqj/SHGViz
nrTvhO5vKsbV4pjpEIBAgp3KxaKfGo/v7ib4/8I7Dfd0PwFBak4ckMBo75hwO3/+lIYHWmopqP7y
J5g9/Fwi45ZDIwtpiF5m4sfOUJU3VY9Km1A4owNfYSOJRRF/C+kMbw1p1XGVPrt/ZpDMgEdM2zQ+
w6B4FIgmAso7+tgcVCxKRgguERZxDXt49Vq2sdxa8AiiCiDRM5SFwkm1ycZJDS7bNjWcD0BGVQ5J
eqtNSds/QIZBY8/8/zxqw3oBTys4hz6c3F73EwCyULVsKrFbGd2IBhA8PEFA9OSC/W8yvXIDka/T
ya9mg03QKtJU6WZ+NJsvF5t2U1LuciSPnBHAImXRO5d8BVGZmrPCrMTc6rZeQKnGgeLpXDGyjfCa
qCbrswPl8sLudmBAP5fAEbtFvEJCaX5hy4z5OEN86vUvYJVe32H/E5BgOvoeiU0VAM5NIF0qKCmq
KTY5pvRrj8oYi8Ddz/h4o2+g/PgGWr8SIFNhdzzjQxlFnh3DwkqmARETHilW+4YAgllF/V6mgVto
vy5ApidCAZL6qsQz3j6dBrkH/RmcrfvN14ssnewkBn+EBfjXqNAE+byVhian1jBrnQdH0w/u9JN5
pfFv8m3I1Gl2zvgu94voQL7roDl2gLtNobYTKJiMsOGnRamX3hsK0rcEo0P/35Ul5Ba3QbM/2eYd
EEVFb1wqYUTQeRpfHV5HmVS3N2QDYv41HTrpbk/7ZEr+Zk0CNsVa5/dAjP+45cLrgwySnV4M+M1a
eJRO+fVOr3YjF0w6xynhbmq5dJnpMjgHElyLuahQme4xzVvh0DvrvXrxmJUIaksRd6gJlJg0sQhS
NDE4jsPyR6mhqkf2XAu8BMRW1h4qeS1+ZWJVXLVteql6fMT8QhNP3eyLw7gj0sFO+De2pjE51BDq
ces23h+PCwYXUfmmIpEOp7HkheScKkhkqsYO3qGt5bpO31Q5PLmBPt7ufTjyBAGKsNDWP5kqbsQo
9ksZvopXC+e1SzJBtZC6t/mSjqrmvUPG80h9kqHynstyzR7zrMj6sM/AY1rpDP8AuEQ587MRXBT8
t9WFY2KkWEKZtxrJrZz/w3l09zgQZ36ht49qM2o6xcJvwqlgz7Uqop7pW2uo099nTKjqTEfVQQcs
7yRmTF/aZdwcA6HrZ+j0KKLvyLPsoDJlMVJ4vC84q32PzClXpFqoycjlcRGRRXm6WOdEY+EZU5Ll
3xp+lL1SEfVzXPRWQ4dDw/kWB/EGSY0KI+3u6ZTT+iU1wfGDHdfhJ7dbm25sYBYqE0L9XPWhk2jh
ODx2YHhRzq3YSLQ4ip+Gan2DLjylFfd8o1ODIn3AzpCVY7F3OJHO9s5Ujo5W0eNDup+OPVe2xXkd
yZZuKYvmEetxueH3Y4dL9sQ6Ql36PXQO7qVRUGSwdHEwujVFgQk7K17vcZ/3iFc/61T6aRhJBhEt
uthZV7KDgJhMH3huUlW6dyVwE1+njOsGty1mKcyDw7ErC+YSoT64xZ2cR+aXMGs3nuByzsMeCMD3
oK0P9Y9PpOopgdqMsmxYaZJmcXsbiS2LPLuL+UXPIuO/+O382zE8VIDajOS1eWIoL2UYY7JUOWpc
jA2uHwQOb1MlhM8JAtQDQuvYL5s+Dytu2t0SiSJgo0b5frOYGilkGGUcg+ugE91rV/jv8P4Ca9Qc
aNUWplO7Ow841DA4da7rwXP4Fux7nrnQgxaPKLy1dDx0NOoI1kC6XJdtmDAg7ViOZnkL9tlkjZDR
9qu9BE5bI0UivAn0QaOLlY3S2qdu7KHeiRvwEmy9QYza4lLFI6XGhbsRIa9WWJRHJS7bUuqx2duR
onHV2r/cMMeNUrXkzVmLi23EQqk2Dj/J8QmAvRAF0fFly2iMBhpSb7nx8Apow3V+nweND0euXvun
vSedfR6TdSFrOidkOKsKQbI6RHOW5+5GK0sDh2DvbOUbV8is+fDDLipWydslPDMEf1jLEAIbm4he
MpgV01Mcc6OzvkKQA3ColYZYbUOqAybBCqVL0aEcK1Grtk6pnCNlwPuaTpl+jgkOf5xd0W2egI5W
Bt1udSmS214shgk+Rp4ax7slOs/YbF9CMUNonlWVOB9qrBdYwS/wUAnYIJDaUAcO6+sJW7nG/QxR
g/KDDwxKoHvsuprjht++xJ9F+NoVLXZqLROjobYEcsIgF1+3rgv8w5x279nPKhEkMTHL0lP8CIny
Mco5gvZiHjvJaLRtNxXr8Znvt4MoyWfPVB9ajJsCD5kCLGKIwMGNKBaGV5pdMd9XUrbDF6U0WE+J
Y7FQ6h1xwnkil2JF4VPC8o8Tqmz3hzpDeM8sVicv9pwUMtukO+yvQpDdVk/PJX1cf10q38tpP5kY
+H2050ubt5tz1LMHwck5/NrOlDJEuQ3L8ZOUBLdLmtcftDRVVK4f4ULGYUi9hRV18Rl+5Kh/uPr3
ihu75mpuIDOfgtN28MxUxkF1FrAR7FlZl3ztnXFcESEA5IoFL0EMj/psPxo7lNtjG6wOURl/eYmk
sn+3oJwEmhv/hDpj1OuRpSOyWgVBWPIys5Z4+irxqE92Mm0fTcYfeAHMOlx7EdCp5yWEGS36qGv2
C5jS6SUY035YZAvXvJvf36Nzu1392Xa8GZoisqA1iR+PQvsMAnAmCncLVaj1f2FKAqkVwOPOEqtD
DU10sNkzwnO1TnpqwxH3l+w7Sd4guCGEQa4QDJvAfEzOZVk2y56vVhAxnHzkvwmgco31mE5XCY19
H6uaV+1bIZpqI6Gc0NxPyM8MUGiBTg1VdmcjagSq2yqYSE2pC5W5ooEI1m0645AVhPm+zMt6NdFM
7BrmynjsbaxJShBMBPFr1psFr+3vjuYvJ8bI5Eqi9yWGM/H83RKZmE1TqUJdyOZIIHCgZG0Bq6yH
aBG3H0d7KPdAM58fkqd7F0OkIl/nXGfKhbFpC+aqDsgjyx01fFBTezfEDq27xsvBenz5/M/Yar0A
cB6Dg5sGCtqa4pIxvqVS6ZIke7YGfNKBEm7z6CHlG5AN52MtAvFjEVHSvkID/PzjGk5OVTuWsqFF
PqNkepFjxdCxQ1hvOrIyj8/7Alq6qfDAES1JTO7TajGZtwzMX/myxDJLuI6BG+uaDF0zS4w3+Qz2
BdYtFbXTL4V8lREjfVsRsIbpOsm+9UypAFHyuN/xx0H4590EFyaWGtBVZjNRa0Kva6yNC4bAnOwR
W3Ef3vWppBZwHlnzxL92E+qBya0ObQQRS1WUHGR3+gtYvRXmsv23jmIXZ+P8bjsCo0T5D5qJuXu1
aC9zEauY82uU8oOJZTP+Chq2yD6xwwN/aLKLqmvFFca4nRJECWnIUYGvOwafftuUgfLgzOW6BS5M
Kfuqo9tP4GNkVvRQWsEq9XASZwv+XArz0hTPn1RmHUdzSnhZatdyF6Ol8lo81VcdIM/Nu53uu3ms
wqvpfiu/YBVSLAPIKUQJ/cosMYRO5LsudWMONoBN32x49Kf8FPzuc7wYZ0YkQKH7pmdJ0ltf84zu
Il2aQbFD02IXWBXdZ2jffYvStEUjQvknM9M5fJ+diUHaE94Cnz0kwcDU399AsWkUTaa4HcvTEVFZ
9wZtga5tW5lenZHyKOrp64lnaZEt72qM+w58t77V4MqewUkephWjmXUi8bYpxfooDN99nX5bgr7q
WENQGUY3Gicv8IolgVwalYcw4DBlq5rmfeRjHV1hq+qn1vMifqFRJHEgmZgPreodvwvnKjGY4Jfj
3Sww6900zCnKMmQOe3R7VKCNlXC0/c4BryrtABVjrjjU49KYvHBXrEu2p4Fuw8zr7GXDy/Iibj+5
33Pc9rtKHM+L2tJ6rJB/E8+o3bENDkOPTnCf7lB/u1t+sOmYWEU+/pDditRFTNZQlW4PiZTlRhWB
e4ANsx/3N3Cx4v40vsu0Dmi8LAkv292SYhWXJOu6g6ySwHf3P8II1ZeSzPz/CzSeRCGqJsuL9rvp
ST/NnGdJioqcDB8GOMIJ3jkocwUzf3NSOkch2DyJ/F3+nujQeIL1xWiTQckqEwTYSy+QIUCweQ/I
rxbzqBH7MIl8emN+6uhNrLrtw/XUYSRAMWcow9Nwp49Sew81XJcCJXIpgDvnyogsqqOFWwvqicMo
Cm3YweV9WXVuOYu+4znSJE8R63Lp1z7cCbz9XvHGNXv90V6dVQcgUeTrUiz8D4opOQ4XBgcPLv2X
IfgVE2xZf4R6tFYObz75PlONz8idqPNKBnD+i14TnN/JNyb2YnnJZb+UXjV3X+deibjACZPCqCFI
GRpUYicw6lmwmxUARXwcFENImX370Xap/CXpRv+ZEC3Ua06OAPWqMZCEuB6sVva6wOSvw/3O1Hx6
pJV03/aiXsIWvUDdDXaHffhhHrUyFC3US0x2yJis7JEDqfTDqSlbnHVpqLYxdp/emReN1tiUa0GT
rA3ln7CaVHkjCObFooGRQkAbUwOd2cpyINyBRHc+7YdycjYAddD8V6/gba+MtG9Z24AuFz9T8xWT
lyNgZGqBfpnVAGVnkaJO+4WQdQockbiKgJFyqumbYIURhMapvcGaOKDNhScqlW42slT4jTNxkxo3
LMsyZt31E+gLx1RMTK8EGMSHfITWwY9LhVan15BBVdGaEbubQ7Pvg4Cpx/dHzRzvTWn8ZgdyuVL6
7hdeihiWt6R8DvnnUzbCVbl2ELWnf2a1v9XBNFkCAAfwIbwKf2FnzntSzW30bWrX2MJU72SnwWdR
6MuoxwUiodZ6jEc29aeSI7vm8aQSJfLLfm7Qb6xH8RyDIWTqx/EW9ihllja1rgFVjluiHjwGznq8
oj0aD3qaVFts72D6xqMi7xu70pB8U5YaqrHzvpt7LIUq7pGlnWxmy3Y1zP5EIEnVjIeeL58KKKdX
C40LRlh34i8QMvfuvADy5q0Wh9ktYq2VhUoaPiO7d9nA323VlANWs4veI8APLjEeE7QdKhIRDHJB
8XVPYk0OdljLPF0jOydehnE6UBSmSRsSOyHPULQYyoNANE26nUp/gl0Kk7qwGpBAbp4z6O/JQMil
cb82OQGeCxyblnzfr68qTD/XM4EfyR0Reg1HaoFimU2dKy5iCrEdIZKISRGRxqsl6bAb8pEu1yG+
kP1rH/pwGNIj+pWqUK6z6ndyfQV565CaU4wRYx9D65ofBKLptvccZDwN2O6klAJvvYPj2xAto7P+
1Qq8e7DBGpDEfBHPk0EiLIvo5BUzVpPY5XaHIxKcXO68axpe8mEUkWbABob/JNAzp6SsRbZbX7TG
vcNliRLwgHDcc2YKniDo0Z1pJuOjJNSu6wm8/Qj5Nkfdx0eo8ir3aywSmWB0UA5Lep5pVS1NUK9m
iiLrkFfXF8vlONZUc/1XROEDkbSMbj0tYXj/AZqkCOx6LzwCggL6buJ1u6TbHVmofSCq2gkD6rTN
e5QrOR6w9EoeeamuT5WXcG4Ir/AShzsj8mmHnSoo9welgEWxUOsoBUp0M19S8TDL7/hzkM12V+HT
8SgecLf3wlo2GOZKY33UMIoR2D4BBNpokrdA0tzuu50WK3Pjs5Yxv4m0KyD06Esli7HeYu1ahbK7
8qLP/YBlf/IK73v4hL1jy9CHCO7b9v6Tc2W1vs9OqA2y/J7J6tsirEFAZC+OtBInrLNSZV67frZy
BR0VIHGWoVsFIHhg1PSHE6nSBpPeEXkL3+vdcTOJhdEdfPP+AFg3H+1uBGcuJOYi5yy5gROF+R1U
0BqQyfXQTnw5fSv2DvqgG8BHt8MEow3tUz/lDaOZgRsU0pEBOYo3AyvJF4gkymMRRy9zun0zAiRc
CgiCVQEBFBf8euBJP9nRISth4GYveLNfyL/D18r2JGYHoYlpuHnfPFFkYE4mDVFlRvhCLVLvVIKp
b/3jzuQcASPAo+rO+LWR/qGINVRcBVUYXLuUU6ff5nDloD1SIxgS4un+3/UFOEIXigpmPBVKgJyM
QjUuIz0bYROnFgM94gepBPcFGLAYeDB8M38IVRlpT6VkdGOdRPJpBz6V6kzDWZL2THMESvpduPPm
PmfIJFzzAFPmGi3oHdgigeeRH8jPJdxGPvR0/gEbAJKG3Lc5skMH5AuluGNNidXqLqzA7pgPWVau
1v837HDkf6lghxCs/0YLinPgl7VYWyS4ZOa1nifXF7UKlKrBSem//IEQ3VpWmhPgZTUmYWfbIuQB
R+pV1SRTCRzsZpd5Op/o5P/gV0SXMrTeCybZEcLoDddpEiwM75P7o1pD2wtOSqcinVwuJvfMnl+R
zlcwPldRXHkeIenrbtYx9so2hqZvgwQGURXZmVmNtnxTMHB+F1jYV6YS/3Oh3dmAlCCwTyQYVe8u
YytiAp6Gp88R1Tyg0DGdhD5/iGqWnSdBx8B68+TyDo4bRMqaQvE8m3bKi4fBbvYwfThjPdY9u4j/
feZSfoUIfTgknB2zLCyaby53dJtBUSotpUfhqRVPezh9wmyWxJ0KVFA/Pinz2Mn7LvWeKxOeT0us
0T2jPpN8Ta5g6dR9XYRmUP9jJFPKOIUrVR5sKa9ROBVQgVSwNCm2NAEXvobjcy0S5GRywXewF/+5
ErYs5brvVRJSekT08HuixpbCU3oZKkfi3cZTjzG332+jPUNXIv4LePAB0UtrOot4nBDXPcsXUJZ1
Q64yLKbgL3TrpkIX/ajhLqr4NRiAgxF4fqjhCgfI7P4ACT3yxwuIo33AzUC5DGYr9TL43Eb8qbK7
6cxLtspMuF5eA3urDjCobP1lDnApA9whXh1jhVdo9/dWDfG113BPH3ok2PF202Yua47OjWABFATv
LYYKpEoI3lR5GdUkiO4Tz0ErR2ptdqjP3O7yWcUNRJl2x/eX3hXKfsHJKY8Ft4aP2D+rU6tDwB7r
oQOIHQAyTjUG0Icb9n8p4oYU+MOHhU0qAxJvgB/fFXRumhkm8Zy9r/hSL/l92ntanIN3kT0eo0bV
+Z+sL0JMA1ZRu4MXxdrjeon69wQSpas/45rWAA53h4icg5nHeSJ2l+Jb7zZdbljOZKdrhLcDNHaD
gw9xQuhoIQtli0kbvRk6381UwAiorzkQLtcGdmhr683xodDXpHHJEl3gFvSKRKkDorknYlRTfxAR
x4hASTNkn2w8mgbIxZxGQxX5Y7GEk1S+h8keq/eJGcB0oNI2dQk4Dheq7tMHAzQQFqBhkM35gxjd
5IXonAqJ11h3N6iigHcd1whGdqbL+CqPaduk7Nb1tKdPiHxvBLfNrVBjpQJ+Nr9iICQ0GZMmpt3W
b46rfyUBL9zP+l1HwHMDh9HSR9Hen8fe33JAOGaRj3X7bIhHlho/aTtrtY15a1EufpG1uRgkMTXx
qu3ymfdhWAfU6AghbZxEZyNgGBo4Ta1IR7bxDpJldnons8Jy9ZC/w88AdqyPUo4WbcKdGbXVg7Vx
ncdA/yOCplLhQ/04K/IwsNu3J1RoN0cW8Qk8mjjplmkZJJrSgH8Bd8oRVJRYunsy8QXQ25zvZ0rk
E0SJ2xSZcIG8epxxYKEyD+tmFTT+7XLB8BYilOjEKzvPC9OLMQx4ee2O4/IzLwnLduSpFOrX/Vg3
eIxbaVUM0G0xtAwbNE0g5qqzaYFKWDoT71bMe/zl1hmdbEit8no96A5ZRdbT1fUDAnnNjP44LfIn
m8rCrjRgS/kIiDG7rz3g6mssE7XXaVksPyFvVu2Kb3lPGWYJAcF6ospD7sWcvoRgPYksaaXuqaMJ
4KpHqbnfMlE7bkYxyIz8+4YRm36ueo3b1kWhQKepi+wU8VUOpB4w0wFvjsRSf9s1yJuIhJHkYzR2
YCVJnUku1xwQfYmskt0iO80S57UCbOcy6RxxqRB831V3n8hfEq4Or8W8pl5aFULXnetX+bH5d8Qq
/z4ocWzy1kFp22iYFZryPVnbCsZYEmHEJbWoNrqV9DKisxH+jXeEMnet0oRphJbzwTi5eLxIcvCd
FPJ5SJjYWqBlCvIS1LoMJ8YCSGtNPw1aRPio004245NR03XkNUi1PPTf6g21UI1rf0pfApdJkwfo
39HrXpSkHgDKfOcuZJPWV5uORyOtByDF9Nk9fGuuiyHT/QsvVf1n3D5OibBD2/wrkAmMej6GpCW/
J/7+txitR8OiehHt8YM8nKM9ULxsWWXz6pIRdC1zZv4oM0XEKjSv48OzLiGhYuO+83US3AyWObTu
PsMFWC2tt1hvEoNgD+q3SZ20jscfm9gyt81CRl0J6CRaq++meEsOdJkFuUhzQQgYQ0UaVlNEcHae
OYydujko88wjpV6RPLFl3Dc3pspFRToebd34QI6uLD/VXnkmtjIIVDYW1oTvMuZAS6P95ccglEIY
pPJK0EYU0ZXCY1v6tFPPf2V1Yh91Q7WvapnE/B5LCJIgqeQMAPUvLhoSgtOcpVYOMwbMmnlkP1yk
gGxYpKHtcFO1JyYVXPE/I0DiAqyZb79Vz4eQkpMrsmvBkW1eIgOXEmFmqgm5PjVM+Khkc+msEuNn
S8g7Ko4SAqjRHV8VPLYx2O9z6yMEH/Ah0R9GeCJnnWVkw1xoep8NTQYGoUoT5lD/HTzGwxQwhcgT
ZlEweWEp+VxwlatrmGnl2SzwvEg0sX6d65RFkVPk+EV/sbLssKR7HYvb5dyAOgHpbLWxJu/dSGTY
WH811CUWoetHVkH1n6OqA8IcTfh3m1GC9AiCbdjqHKeBjN/1MsGJGZDLLuZ/oGlj81Nl1PpBx/jj
CWZqn0gYukPnqtv/xIWmlpNQ1vPxIFHvnKg5POZ7vStVZFx5X3l5JI631v9Imz90s2JiwvtgKJxa
RUj4iJLhypK9ypd6NN9tETF60fpua2bqZRaTWYcXXMNVIpq5eDQPuBYyoGBDOtqbqf6DprkdHN+A
jP4ge3g1iOJRjE0EqlivwkEffst6GPPFizijs3HMrp7H8YlPEfeHiODqx6IFg8Phq91ZOBpbrxTO
JvXN9nQtpxv0Wgkr1lcF8iCog4Bp8pOFG/HuwWANJmnM1T+kgALwWOl9x7teSduerPE/mclTYeFK
6O84MTu2FdVMtKK3xzHtf5lqsgtZEME3ZSgwo4j4sz5vf5tU48v7myKBPHMPSPh3x2YiP6Mjf2Dl
H8kwUhpEMnkO1XNBkiUpA9pcIukL1zLORupb3/wTIYQ4PphwFzfkp2Xr7JcQGzGkH82DsvaUK0Sy
eRHtvUgqBEwKg0ZhtUL/hKuU+p8xX0uXdLKI8NKyO5lejYpCpajOBTRbH4CNorWlvQrYzvEJxVE+
6pm1nY+CIMX2wxPu1WKDhgvqLlNXNOgDNPypjfYOeTADBuR3V2GC1L0Ayr/ZJ/rZFrknbtp+wRaK
ST5ft/ZyLWq+/PZe5Ga9jydxhMou/QPoZop2Y7soU95+BUS1qe5YKS5aIPZ6sY7dtNM/xfsTjf3t
/tKRwEL9DWY2xzM9IsiohK+MTfhM2xnZkvf7DWkRwN6ZohB2pEDReRcs7FJxUEHA7ab983emkoZ/
MeJJv3JkOEOrwSobRxjB5FaD/6rxoC4P1YmKlsOU1Q0KCOVDJk1C3yNlRWuiKXWwlnsVnS446p9X
z4ZPTv3aXO8sI8iyKgjKri5six0N3Loou9wjNG3h/Qo1afrUsMbeufIDBQJCiQC6wNxwqlOz+FBc
Wcxmx2gLfr7KMy/TV81Uc10zuLgBlm2YsEYBHHNmREKJzdp6iohscfDvbb8GkmmO9kGUdBILjIYp
cQwI1gHXL2aiB9cgnPbKT5+NvtkK/qX+oAhxs4Rpso2frIBthD/FmVIDEJdt9Tkkk7Q2KAkTI3kc
tWGPY3IVgUQ2JP9vK6KgTn6ia0gZttvPlTobKNnNED2kmuqegmjZ4XOwD7E8oN+f7wfNjz+4Y0kT
fWHpVHIt00qa4qcqCXgQfR+sFIskI+7LOhpzHo4BHDVqgHVrxq/sHDY8v37WwEfYCEeT7MwkNOa9
9r/X97CAuQQfhdTvLrq4hK7e23lU9aGONM/FGU5ttlszV3Dz8sNrnPjsXxMheViF32H+ODom+RW+
utwhPxtcJV8a6ZzB73CNOA2GDwCpLz9hDMf9urjI+0bkRsiOD/PPkD/RrgOgXpHdnmhL81E082OR
sVys2dkPHn3eBr7U7oC+YcdjUl5cFLWUKrZGpqeBGVkzJoPofWDqy1IKnnS67h87mJqSxOHNnwJJ
fFlFVAfgDupBS7Gh19nTvqvFQmMdBjvTSPgP0Rxkh0csp6Tso5LDCLrWW0oQq0TUZic2r2Mttslx
M3CMC50hqsBGskwDDpHcmoIFUw17TJ7n1IXgbuaGFrLfyipIhnvAPFozsxA3ch1bIamLGpcIFJQC
1wWNIg4si9B33BAqlE/nUCPthY0h7FflyFJ6g9IP5iNvp2FssB7feddqP4yfjIdffzihmBIQlt52
4vlXdB6OxGRN1SHmYDI4jtRFBI8j0jrt0Yv5SfFeDMYHmTkLhu0w7Nds6eSDzydIml4N+UUSbMpb
rmsqpyaaOFE1Ppq6a9Y6wheYxMw/Z9PhIzX7lnAoQoxvncfUOUFcWguCt4vGVN6sOcRFede6AZhL
Ga6fv5CNjPZpOG0QWmgTss24AIba7npcwnlps8lCW+oQrurSUa6AXSJR5DNGmvjG8J+nrq7av6I5
6s103dYRAGtDWA+S6m7oOf+Jgtg2oPIvaHo7akm0CIZYzZ3r6gflJcS16A6sRfNuGFRKoD1pEMGv
J4zvDfhgrRblcPI09hggVulZIpdQceEydpWwKJ6r0pAsscWg7mwW8PnCivFsSmVUX5vHChNoNL5s
PKYkcIPXA3/4tdtP4KMOn/2S26yrBqn23smxWYRSVTuXmw120djCuf+ZLku4y6ut8WBgVTQRslGP
zA78sk9R8Pr19zRrOzaIC81jl8zz059RWR2uuMHQM2QI4Hagr72Z8jL7vTGt97vefe7ZNDei5Gq6
NqMJ2MXUa5HtTk4EPddLWXC39+sb9AXtv1RbRUTrOUd3kcUZ/AnU1qKKzE9ZwikCr7XOqMrDIWR3
NchoUEEs8GkYJ2eR1JcWv5m3CEEO5RFB5GsWEru1/NElpo894MYxlLDAk0YZiNXwuz7g6thlxB1B
U+qScErFYSho1y4Oq5jzSBcW5dNYPoOPXp5jNq5QB4HoI3QkI1d9ilE2dYrlfYICllsv8HkNOffa
6rO/Z+M33FKxiwGOiFxJgBXKjzcVOMEX/mS4938tvTcXQ4uv6R680n6bVx7gF6+1eFxfQx1KJmHq
GQYHewJCjqH1CtPVutCTsU8uE7yAZDXdyu81D8N9G8FDWocnLJNE59UfusSmbYgxaK/9GGE8Sgrx
prfSxsKktaFsX3MGwvMYXx81Hp+NGvh8HJOAJLSuePh92IlMN1WBkixIFs18VBpdvvluzdzOPMYB
qHuuxLvpsuchI8jXdjh2QpL8QQkMAICpvSuAWWgBy7we8pBM0/DdbgbhRXIhelwMmuxxgI+oGjVr
lzR8NZYuMeJWBmEyJQEKVBOg2JuAMRJyj010P0x27g932wDxaR9wTHqFK8sdu1fJQ14zHDBfvIgA
IjPIPU9iIyjpztLJfxiSfrfHkvaQB3+n6Y7D/2LdoIDFtR+o2C/J+IEBWPWQetbRpwkEGuOeW60y
El99UUz1nrzEUEkWXZxHOBLTkP3Ni6coY2NEUaQl9eo3CknEuVeZsNx3enTzdRIJiIIfWKmHV6HG
uLUxHanX/IAbJkWU0eyrpDEN/NPfqWOUqWEzipL83P+AmDfgiPH6PJNeMxYAVOE6zdJt5iROdWZR
+rbgja7qGTwFZAd6Bv5Ct8OVpTBaSSeqs/2yyoTjyVVzBntNUpx8JXLy5TWOjI8nfhFyO5/wXcpp
83hytXrL6V7xh/SQ0VYN6NIAuMoIrRNuQrcDGNTdgIElPBT8rJrPi5wUBjJXIE8eZkfiBwkzBjf8
JPqs8aWYf/bn/JNQ811a90ZzvqqY+uaMiZ+G5VIB+bEBAj+6wS+brsdY8+NCUOgtTXrCFSAbxvOL
uJFiPx96ahA7qqVUHvCSXFuMTAmOikrYh7LIiJQReoMA7HsH3MBTGqPPBw9oJNxGdgrgd50JdkwM
yWc5a3HT4HrfWu35emE9B5zbxGfnmx9Y2vrGsSNNl19p8d0sS30Zd2yAdELhYNEA4wz2pZrT7QQX
WHtD84w3g+ZLfIZ6+kOIN7o9DJdrNoM7BGptPTnppYxF0bvnFiv1m7OH99RRsGh3USRxUmO7Qsg4
FDIsLIYI3LRfPu0d3EMU9rfLE8xRLcBQShW4+uuGFg3pKGKdQ4SSUaTQAjjBns7Ge4ZAID/BiipZ
pBKF5ngPPJ7Z4Nu9AjWsdaQ890Numijs2u/wE2xfsMKNuUA9T9HNrLF2Ao77MZa0G46s5oPocNgo
QRzvV8d3qiAJ1ehqrHO7Lvo9mGCX4VJTrb9HT/rb1Hh7h2qVopNEJtPV4SA61Syvq56tW4Jd2DHu
CxsIdZ7ilL4kduSp2qb/94tYJ60xf2Rp5fYoDRkDIb7Itz8jQ6CzKDHD8SZIJXyRh9CDxpic5NIq
r6qYeomchfz2PNtHtgpKSdFgnUqlmOzNA9Jvc/I3j//lfpYO7ilAAMTggwqD+9fO8tlm2jim0baI
gj2KeVlza7SeuSySYAErkMiSRAUjXr1ka1ehMiipOKgG6L9kuXFR8b1TDCTik0b2XpCABcTo3Uq/
CzUGhSCBFPvHPHzSaETg32mqhihGvCD9fbrroGNYnEI39kBBA8cfZ65h2vXmyGwR5dfbIXNUnqP0
JErfxkY/0j7mL5DZbgClfivaP6bJmBxdPZQPo7aQjsIrvl5FvvBWqK4hC7WLmyIzvH+Hms8+JChE
xcg1RsAv/VWyRP24bEsNIGsg5MRkGAKGMBv88vwm+sbx2GbJ97yUBU5KYjbPI8T1KXCKQGHuyu22
qyth3vC/h3VpBrU9qMiSsmvbDvog86WkVTxrLaqsLCreDsWFtNY43TC3Mdwii5H/HxdVq4PtidLi
ZnS8IbD+x7tRVb9jTJwz/X49XGYvbmcT/5DepwtwQekiYlv4uSCqxRuPA3TDSiSZm/4vTytJBXbC
5hVgKQPy/LSju0JQifRX/Ywz/6fFkr0VNY14W6W+WIyMhSowXnCYvxSO65wfNfe9VexC6qbzQ+m1
VqtvMsr1ZdLHVfzfd6atdmieAvAnpNj9kT3YX3QuneeHd9KyUBxf5+xrt9M8kY+uy3yiKMrqGsbg
plIRIq5/ygFNt6C+QsdPZDOMixa5o5fgCXbazUqdll17A9xK8f9WI9j8S+P3jMF/+LNZcV9aZHnh
G6jM+JtF9c32Yb2zVSxLnTpy2vbEyqYLhokOUdztlYCVAZpibloXWe1zIuc6eAtOmGU5k62QQIA1
xJrinGH+JqlFFFqfhPL+jyma5tOugJWGsbx4RBujMKNvE4V3c+fBBbJqbQgwQwBTcgLRDZVBQrby
xaN0rTwBSOjST2qC7vm7fXvJC+nVwf1gez1Bd5gqmkWGAFMWQZiiNRuitVuB1LdOaP57GFFpJ2A3
bY5wGkPd68Lw4lbP26YF3yQFEFaP4wL1+grNcwrBtpQwntlTowa9uRY0cA4R9KKz59Y7Bg45h/U1
FJmmcfo9sP73wKQFOiHlz2/0SYLM/FRirH+LDPOZ1xylfbXXDQVBnWmG6nXvBOz62h2h0bKPxTMf
3VWzhnugHLp+UycbjPeHq4Da7STsAWOEFMNjePt6KrWlImbDppduOwLKB0qCIXhkUy9/ubFq1l7z
P7zCQIMCdPzjDohRg3YFaE/iNWaPqMj9VIPcbTXztZ+X2JMYXZYt2kjarYrbcslmTutNJ037/NFw
ZSqtW5H8ZclhcoUbHV+cCSzbst81OdNI4IoUuctqsOqq3xsJ+p7b1eR37S2RyF0EQ/2xX4NZpgGI
v/vBjrvoCyjrDVNJN4qKTFzMoZALlernWRFWkZSj/pV/M0Kj6S7rJKQ+pLeBUloPmUaH7GM954BK
H0IUEPJMFgdps4f7rfeYkXAPwpTwPvy0AGpjExe4jSiyypoDlUvnGXENSGBvJIfvpjxPZUHBuGkw
kwqnAFc0nheYzHrNmQzwMf2zb54z/CAr7oDtdj2tTI8i1L2lf2yworZLKrlrC8oaOm1hE5JKR6Z0
RselYJuGrAE6wdLT12BeN0mY9b0gMxMcTvVxwfk+/0ls5iOU5nuclUfLnVWV4TJRPcyA/M63njcT
+kG5mm2uhCcxckHOnxNo7PAjp3fcbhdUlpEWMf+C8tJEZY2p5EBVyfYpqv4UvbPAjsyTb+ZlfN6Q
8wQqi1DSMLYW+iVCnPfydRkmYG7CiH+1S+b3XkIIKr096aeCeMtsfMOvrrn7vuuSkqNN17/DOxdB
9tz8c4FvD55uC49bq2VloW+C/6gCjkgUx1l4OT/rmD30ProFmShDmHFy8sPi/v02OhpVug36pdoj
BORs+jnxZKTn6KbdB/1OA/bl1MoEAlfMlzAcpo2rTJv28TleAWdc9emDhV3Utu/rJlNQY4Un9tSl
7u+s40HJtTQ5aDjBGYNztRPS8ymGIGm46p1ep9Qt8n4cbG8j0dFASXQ2XSo9cWaDdwWSBBEAuuhF
4j7O5jMBFQ3Szg9Nqns74pzkbiQ0VkwqziHl+EUIw73Zqk4cPu2fKLGgwgBAv2/+LyGSgRrUlTMm
oyuR0/DsMbHyrBgjGXnkWxQTGhwVaEGbsiWa+4UKpXcHisnk2mdWdFsitExbqravnu+OIKZ6/vjX
RsDNzH/TBNJVkGfexG8aDwfEctUyo+gK1epHGpFqf8uPXZkbcc+0NL4oxoZQPEW4ZdFWwV1jcg/g
26jbwIO+P+yrDdIM2xi3k1y2hL0hEgRo/9tj1/QKEA2/93zkgwAPDpu0lHk5q880EgOSArju0rZM
7ZxHSOEO8UaeB7+TkYHstFoYHf4XTEUd+hBlipalhgLdrxam1qCb8gFUTfKdqZhObZle5WMwcS6a
rT8hY+Kwj443Bz/2HCVKzw5+wSszGclLgLlgOuOzYEFVr3wU/OR2NrsCLWZFgtoR3IeH+I0kcoyB
NXOapIeZKEz52X/o9/iF9bCNOPRwqjk9lksXoY/7da69ZVlUcdS5+LlQJioLkAwCc6XWOqRZBCdV
zeWawyvbT3IArhELwwYSJByjdrlvbEMxdU9LmHJ81a5KX/Ko8/9FlQ+Vrl6SDMDxHx8Fm7vhaXf5
DhTW+mht2Megy8XNMAV66UzmbMl+ZIKLM0zvF7m2KWKPOOG6ru66uZENlbTpcsi7R0afmZayUQBf
AlFkJOeIiMQuT98CUgcDwG/e/07RcGnunRcMzCroEt4Blm4FPE+HReRFwgM7R9JOJuQCrj/8kAip
RPZJyx3LJWhZdzox0bV9yfzRxdSFwr+7ELDllgR6kBdm8/s1yy4i05iDfEVm37/SyaGpTJ4GpyQw
G3Q6pq4WgtwUjA7TWUHHggzdzR9Lv9ENuOz5UEC6h4mASykEDKlCT+EJNLRyPEK2ki4sAuHh8GoZ
GNw3QYnt4Z8NyYzBPuc5e+Kgrxnsyq2XbHtwosJYT+2eQH6mC5TqdACoWncAZ+m3qB1lUZbNM0Hf
2wTnpeSGl8ui6DW4kzsxUQmqQpyEWIWjVn7gYnXHRjY6taOiCrkBO2lB5/vxD2D50OCZ8pQgad5p
7GP8HKXPyGNrxHDbZpGzpIPo0g+QUvUvLnbmputk43fnoak/TzVRs/8ji4KWJFc+J/nQIlyiYyEB
w+0eAAm5j5ImtOCc+bAcpwsXhwMdLxip6dKLb73h2v/nC0E4lSx2CFczSKbL+fsv9sUOSY1uvb0t
amB098+x8MpRZg/HPNBVMq5WOiTzLNbRKQL6QwqG46NI6JS3sDUTEzHl++7aL9TLdBVM8IEGnbte
4Zg7TQIEJYkE/R1nkXxgrxoxJsVy+mguAQq0uyG82TZKqVOE9S3v4bWZzDBCXxBof3TObrDhNIgO
TTxgC6/C1Wa4IBn/z+9BzK6JJM6icuS9OF5O+/j26I+lgzWQ5wSPrDgjpdfFfiH/bzFHZ0vEzS+L
TdU88uO82f8rfRu97t3LNRlXwna1VCFnXxk4T3HtqxMo02XMhVzrYr+WFTynSyHuceDiKYy9yoXn
2aaBnpuUAcduD4SMSEZ8MTYMdjzYcVKe6qLK5nsF5Xz+UzGAoDBqaO6CegfJqBq86La9EEC1++yO
DasvHP30bdPP1123nZhzsRQsDNxvqEVKHiAxaunWcNRdhUClSBhRzkuaRlvxNpmv/drcQlZFmDVK
EkBGRtqlMI9+I0EMUGJg1mo3QwFJu/zhb1LeUybIVyvEdDkDilp1IXLNNdMW19e9RCdNWz2rUXJk
/4S11nXTrOVKvm7XH1pQegYS/DqA1Nzamu/c9YjUUBYy/wv9M+xVj9qBa5lJbvH+5mjmGuc8cnSX
WW1B6o8orQVHj9NylkwtG/nTCMkMcpcBNOQtctPRIU2O8LSqbT4t28A8/LFQdUEfc5FK36YXq1Xf
VCxBJFiG3bsq3jBgayKbi2788dcsrr/FY/NaCDg949/VhqvvO9INY2MLMc/9wxdtOyLytnV+ksy7
9wBAhGohxj/3kAAH+fPGIzkwDU/NK1aZVGV4ng0mXfFIdvCJIBuZvwVNfMsx0Expytc7pfAweM0j
SEr7ihzfNAAvZPnT93kEc0bTBPcDp2Jys5vuQvrW1/TZUKm0hSg2wv21TDh2q7lrZ0eJZRdt1Y6Z
ZNhRAblkO6Qrd5Jd26aFxKJhiM76dTSOpQeIzxSsi5WAjybQ2xpyLLmI0A9zaWG3s5cRT46QGVKr
GOwUi+XVugIL8kMdrtE+HEBbPBFPcwraVTlVnqpGb7nWAq2YCxhethRpIpF/Ii5texHX1cagiefc
3gbdDlK4c71Js7qe4Ll8MOu30It1rc+e1SUdOMd9HvzgEFxsf28Ula5VvoZR93VyWWk7aWj3KBuw
KHOd8/1gLoAV4VJMLWGk8TJ9HwWKKpCiJJ/UxULlODGMGin1R9QIOOZMySAj9yzzxI7kzQFXml2t
hkiW4xzvDe5ClavqeMAjC76HxQyl5sD1KEMHkUTskFE7tyMtDpgoc326GrdsEzopvUdHCjNWr6Es
etL84h7IxR03Wayl8V1cslQLiJqlSvPSXpar0Y+leQ2m7ujoEMmYIJ5aaH1tuRo9AZGr3FDJXg+L
AgSykCP4ZUqT/NijcAA4LWL5icdTRdO/t9ehZyeRjv4qgpMrQCZi9um9a0H9xHUQMaMTTlBLckVF
2yxoSrCEKqBzhM52F2pshQSRFdN3kDkZZIXyz5fmE31nFKbWbQLPMEtXP/noLw3V3Gq0PUR4jc1M
q+DUfnaGHW+QmkkRV+ksbrH/OfKaAIkDxL3ARTqnKNNkFTAN+vLjZDhoxTjMIutixsspVsjucX4R
O03mO3BKiAbvlvGv/sDWZ+Z5jO1zgjOarypoD4GACsNPgwGl2UZGmJC42XbtDpqSyHU4YnUuV0Zr
Fjg7lnFGgbuLbI+8OzIKcdc5xQ+L4A90VbeIY1XQFifDRvLa0pX4K+PeP+ho6aEsDqkKp/5bgaCl
qaBw/I8LeuUub0eG7JC36nMzKcS32Vsp6DEcIRIe2ZAKL+e47SQb5W5cEU7Cd7olRcTTBtV4GB50
fOJgF/wGVpiUDbcJoR0mxQTYdu1F78pNJl9YYSIKwB0/J405vuT1sofXZAxyyeSqY80qzH1Oo28a
Rs5A8f1CKbWael5sV1tMC1Fn/oTmzun3Ef2wQyEZeFX3kcgcwcwnqMm3s0xEA0szvrI8HH1wLvui
0qlzHJTsq/Frz5SDzhUDxaHxp5fU1Vo5XefhaaIZs/4ll16UJozRISzGsiW8ViRWioEOSF4AUPpK
EItBhKXnA8OF5VospWKUX1CVVJSiwkgWhk61avzygOhf1A1An0RiBezALk2e4cEMF5lHmz+nMG5B
ifrYRAuAy3JgE44Pwk9H0p+W7uRYlr0D56pfhI2roa2TJV1zErIMeGqGpvHeXn+i8eJrAk0BogXz
0C8cnops+LMWyAq+bss/rdIKSCnNbdEiKa8EeEsdDgzx3IIBIeGY8mY4SAfWE2/UBd42M8IdE9Qk
7hQApBXgK5KCCvgTl13UM6eLiMj0iQP1VvemljyZG8N1SeYok+WlFBdUJvLfstkoicAUIHh1Mm68
KATa9HVABj/mlmZpI8viwOC4tvx6Je9i1Nn7PaPWpk/SAAtPMUhA9TtHugiBqsIU6ooRm/Tesoia
N4uSHztIE3ygcM09P8W9KVDqGcXG9iATTJDL8RQF1MZlsVUtMvikLfENRELUzFnG13xy1KrW8AOM
A8Hfvnqz4V0rJJyi/9aUj/7Xd6TKz8xoIdR7jClNFAfCmbr4wiOrFq0OjsQ2dnWeYhfhbCW8f0L8
vu9fRJ0ciAIWgKUmIRZvm+E1C6d8E5Q0l7Y0BcCkI0OyUE6YI75vIlVhJHy83NSFfkqwc5mw5/yg
Y1pwRuaaorQat7Vvv/82XwzYfzs0VgQ2dfwTb41stwlNM0ZVVr6M+I1GrmTw52SvUAQuleEuDrOo
HlW0mNhYHsNMiZlM1BM1uXQ5HixXO3IiOcwDQg1uW0yOFYAJ4A0bCqJQr5MPEVN9VoVhIYHvmHlv
p8bE5y6vLbZ8NVS/MzZLDUB6PIfhsmR0YeqBpsHjrs6cpJBOwbkPRZdwAGtdtudrG2PMByuyHjHn
Uh5ZoJ1EPP4eFGvMN6+6u8uXjIXEJS2NEo9ZQ0VuG9uVyU45rs3TxMrBC6Jy61b1H/oelpJuxbHv
uoE/K/C15L6gtOQRP2ln6y7Lh9kAJrnotBc5IHZglXrtR4mL2i1q7jEukLAES1z/bFdqaddX2gm4
MIbn91AZX/6Rlx3PhB9A80in5YGT97Cn4rHZFqvR2zeLLAf1g8KmxxV1xed0v/1iCwcmkWqVOITP
69zi72cPSEiPKEltwq2MoSLxUtMsVe1niokVyb9t/rH20aN09HO5vgQJqgsZT7BR+N9eZAUnXK+d
PyStoxfQYqSsIH2NxAQmsuCxMr82xO4QqLcHazwY447NlAV0uK4+NA+2yM0C+pQ1+BHFHkaoC7d+
j0Wo+SH6LSIiW7i07W+TLaM1CakKjGUprl4NqH5W+9vOuQEP1y33+tatJwyxTt40dhzBq/sDFmPg
4Mi4EnPmK87fyK7LNyEd7wkwIrr6EXn+HkndJ72Xb0CmvHhS5OHcPDeJK56/wgb0nCLFb+CC61LI
nNubhA7paKxYAHGSfuQQG9Vm41umJo+YWzGgzSU3uttjOGSb4gFqom5pK//ANzRQM8W0vZHdoxKP
kL2IZyB/9VaL9JlrwrzHqLB7eYKVba7DHrjs+jkl43K4PPwnzXZbwAGtA6AcRS45cD18Gme6AYCQ
7P0wLgT6vbTkYZdyHyA1ygSgWEa01DoaSUdxuDJ1RxruRX9qu4o8nQeCX59Q1xVUYqtNtCI4wUKc
rabVtg8xFfT/rdv7zQy4ojYbqUJqImVXAzuhFp71iHPHDbIG6Aj5KZcD5rjOV1+SH8s/7cKtu1ZK
JMbfBsqbr6eK9fqWHkcVg7O1NKa7SkN8MDuVECsF3/b6Ejl+TdcTl2rsT2QCMOpbxt64CXe5EYi+
YwP7Z4BJgEGEi6Dfd5lxQJPCsgAfrKqTmdFvTNTfS6qyQ/lkINSaquYr6pyWjKUj2uandzOWxlX4
up5m6h0hw6f1jUTSAjUsgngL6MY8gv5WCO83ijnJQuBVO0A6keW5k6P/rfiIowe30rVRc7waICQx
AP/xHUEEdfhnlpVjyf5DhMoBMg1+Ay7HErJipTEil7XwEnUAGf3YdO4rBwLKmzGSmkpOvFwKbGyA
7aLLEbC8cQEp0F9uJhvqB2tng+RwfRSW+gLx2W6ROKCvcqEjv8EG/U4pcZpHPFmp1UnC6qDp7EHg
duvwu3t+1aRn+Yzpv05D3T+AUYeiTTex8QwkQFe6l9C7aL9dwPV6bwgKg3MDhlcd1O72PeY8SJR2
5eWmS3jbC0+eGh/Mzjonr52GyQ3OI9LtT6Bae/Yv9ZY52hivwfVelQX+aS+BXqdUWlrNMBzZaQq3
1R8DEB/lCJplpzOQ8Fm1Hn0qnc6fjycj+UjGEJwHIF816M7ImhTwBOzylT6hZUo8JZgvrGpSKBDz
NKXKhazAYFmg2Ose2+K6TQ6caFXg595EX7xQZl8qlBrRaUIBTR+6Bb9biBe4YMXE7f61FF6zB4DT
vPRUpt5nMsATuiVYDPHbfIh52bGsJMeyryOxfCO3PjsZ5MoGSYcbxJ18hjSnJdIDWOLtcONWe53f
U5ItOv2d6f10VqgP66jSsrErhgcLiKlf1+jT04oT2c/GUqzMopQ2z/Vq2F49otXWFEfULeLGXZrH
phS82pu+6ovRQoonMQ65v5yPLzsftuboq3OyldqFVTlk0A5KDHPBp7/tHZ8s+OX/jwwl/SkLoTyS
cak/KI42PK4ubyOOXk68C43X5xft6P6HS0ojk39Cj48Ydw/D0G7kcxP2jfuFkzGjgj96YHojBdpR
EFC4ESndeb7TDMS9rb5g5gPhbBO0348+W30/wKIabOn6fiTpEX+HtJcn0SGV1gCiDsH22wSM72r/
hRbkiYPyVC7dcRqaEHSKtutuM0DbGXLLAn+VBB/23OvHTuUgDBIyO2ItbYPweK6NDx0VHtKCvPFb
1zqZjAquYWEHTmWYXibY51fVfJWTToeH1gKPvPrzo471OZvlFThJCebkL1Kpa+3GIti9a8QcG2RZ
B/2izv+W3ayOKD+m0KXW5hoK2Ak2F7VEe32GtmDQS9E+Hw6BwRJ3aG1rsAIo2XUUfdjjEKdFzoUK
PRGFnj/3N1CANRUJPykzmFB1e+eY0oiblV1VcavAx2iur9be/jkljtmOXYVSthKBuFk0AtzkrJI1
0BfMTOryREnOdKZvh/sLWIiue9RxqcJLjmiAXlw2et7bQb1WwB93CH7cGwIc9DISYgAayj5a7tku
sf6HmHAJJTmeWM2nJhHK9BaLmn3HkDFw+YKMjzm8jg8oUDxWXcFP8XjP+ufhfE0bRxX9tCnalkF6
tCcgXdvWNeNIc0qkXJYKpJGVi0+B7M7pfnFFHbLSabcunQ0f2gdEZR1PM94ErYhq2xxRoDKczAfZ
MEArqiYXk0wgT/N6KLu4oGJWNL28arHhqaDeS4ujxB+mxmf/bkIysKMn1ddBU81X48zp2S+kf0D3
UwcbDmzuUlZuXVHlmbxEpZjR+nI8SNa/vZiS9vl0sS4x0plugraXpFysmp1hSpvwWJjYLKF4bQP9
IK9/Y0c3ndEras1ALKUUyw/+XkPly59l9kS08KVRJ5jasVHC3xvETTYQ2BLJD17RkDeNlPiZblI0
0jJ2xh6MkB+8rnxfvjohJ2aG6y4yL4r+ZF3CuaAOWogTw9v5Blw+Cz+dPRJfEOk4CFt7rShTeX+0
oo87DRP5AfJhwBoGQs98413KT9uebep8PP4MEtBS08Rcuc5OuDxSIXUU6b6U33Vhf9OfjcXsDo8a
iSEouPB+qhYDz9LW0q4mK6sYXqmOZsfJRi6952tvDJ8FUi3XXUGSP9YfFVsBxt7NsjjPTJCnSCeB
0O4qHatVEm3wawPoraUkM7zVTv2Yu5jd9FolUH6dGpgKSKDgKjmQNohi/Kbs/G/si14koLP3O9Gt
1cgRfm4QYleBjAV7G8YzMKL6VqiHZtqdW9XcqzYjeLe879i9zJ30D+y21nPplhZDq7bUlL2KGmTA
yzaWIL9cwRuwkHK0SKzk9vCwfRFZQiRYqjxj3BkiVmqkDbHbvJ+jQ5okfjMJzm5y6HcLS9xIbBnG
3IPz2iHAsdfCylC8y5Wz3Fg2yPqch6OEHubWz4/OUTZewmJ3Dk7AQUJ6tCCwVm3WDu/kOe4quJXW
Sya9hBD7dn98LZbR2isAt/9SVowktqiU5fZJP/LetMY42XGzI4mWNRmUzMapfjTxY+JjRPnj7st0
wUzX4jhT+ARgKaJJliTARcuPgJMHt7krUqURrPk2+pmNz9wPqMk+VDnIPT1bpza61pTvHiiZUNuy
bct8088dwtQhEaKw2UqrojRnU12eo+dPDHxf3AtIkjYg/If6/wXJgOOl7unmmOnUIVDXFe2Ek68t
wta5+fAdEf0BvTN5jHUMZ+nIO0zHShvY7uMU3q0P8wQj+tYnPm96GP0TwYgYUxwTVv+hGfsUUaUW
aHmaZvroHKX4bSQrIAphpfy4VI4r8x2rwoNKAMea/+Y32y82wTYIoUzhy7SCsWtDsks+ioE2FrXd
rOEyxDDIBhAiIY9CQawUwpkqlmQnvUYgbymzkNqyZoycxYa9gdnifO/detnrA9ZFa+fnXUJeJTRw
iZaqcLC2DSxMkYfNk3x/SCeGYP7GbcFElgNEUz7dSFDr8ENfFVkTyJ6twaJJsNT1DhTtkFr7Tcx3
r1+gcjIdBdmUck6g+EaGorWyN09OQ5cJTkAOsiKft+whLrp7idL2heVhIznyn6BH4yFEcHBQ9QzT
3PzWypCOL5ccVSJmdFoZiAzO/TaUqyRW89oeIiaGYY8tCoP67kBEIIWhbAjpggc8wmrmaF0zS9Tf
wsvxfX/QqP+2PcohVW3L5Ng0WIL1cqkTuzUyVOh/9bwDUo1wB43TvBY7U64Wq1P3N6AtcdrYwhFL
abt+UxRlEB4BRBrTUwM830TctoYXRNJ3WJk+djsX5OGvaF8/n0lCdMaEs3Wu1k/9F4BxfmtMwJbY
KZVC6FPYFapnTJQm8H0NRak/nTA6Q7r7/aRhFdBvKJspwFrKDb8PQcZtRnDFrE14uTzgrllrOy73
fBmrCZyKikklWEQ7GaAcGTXpVsptOwnsux2DlQ0inQaDK+wZf9afzHTeDQNq8waevsZwTG5yfZVu
lFMnSw9aNI0lq+PUDecnBK1EfU8ZYpViMq0JoozteL+mAPRNPiMiEqAGqvOS9yTeQ4dVP1Ql3Rvi
4qiNc0Xgfs2aTgaCTAv+c5AMsgDDOyPrP5omXmciZKy8fuoT/WdlGb/X2B9/pCtiHdVhliG7KtLN
DfoFsSHKiyv/VERnxI9S8fMVbxHc1wrxxSH2gSiBLk9zbcd3yTcLgGom9Zk93QTuzQ9AiVHYpAGn
aEBXZ9wLzIdbs3LcGemYoge/bPXv6+Y7z53KMffFMTUwYHfS8sGVjeLy/c0nXd0fX8MbT6aTFM8g
rQRPR3NUBy/qXNev1pQszfhDkU74netW509yTK92bFIe2sM8xjmJTgW7HWzWEeFdeYqMsHzELKh/
cwL8lK2gJBt1/f3cuWLIeBi1sgex60LxnS7pRJIrBmofYRXyFNvci5/HvAe6ikL6es+XIo0jLjKI
Kg679xkxpGTLmfoexT/o4iZWsj2riYO9Zz74d2upY/BlkxVGfovO970Kr2QY4HZtUn5H/srkX8OA
mrVEBr8XQbylpcwEws16zI85Sv3B2Xmxdg5+/h0rsn6yOAE9oMiPFZgEC0lOmJ4TkgBKudvIH10z
Ov06YB2BcWFke5J2JUWQYkNe19Ted3T4DtX2Ismp5Wxso77ePJspF9LrBvfYisW/gm7+J2vfjfEA
JtWSvbkyuS1Di1SinJuSwyq+82+Tcvytxu9Kwa72mnzNCwjEbOFx2RMoOfIVTc6DqTFNBX5WAb08
Dq6YpFRe++FomZzE+6ojrgYj1+sWkfYjzTmBhgw52KNFOgIh43bGetXH57M4DrQoZ527HLEjncKY
f9Hn770zkwonIrPQ6uWxPEQyJBiwcckiiV19MCyL6OXK4MXFUTpGsacGDJ9BCx3w6qKbCYTBIg7m
29yxOcVtM9SgVMZec2AiZidhNhziTsGGdjaH3UXjBCviZpLJkXcOPtxc2oYOFK1ETM8oeFLrHSGf
yxm2KhX/VSx7+aK4xb7+3dUPCHWzzQrZNx10Cn2B3HfYEwLx1CDJXRSkruLSUqas0xMO/yh0LsXk
S5qWu4rKsuE5QgvSaeQIvna5UPb5Qx5DVpGFui0tBpbJ6Q10W537WmOqxz+AjK7CUussTWy1/CNT
KEE4DDVKsA9RPmzz5ZbJ2nlGA1MSr1Cgn8BJyGczaEixGL6KUGgKtEGknhymLdoW3H/yELRJhi70
Am0pba1Hy22a2rDSv4UfPwRoSqh8BR4bRrAL+AHDYTb4Q+Sa0xvUPMYRCT9Q283PnBvSsFkLEbCR
K9eI7EowC3ODuFkDHHL75ap//qCDF+v2a4b9ZcP1bFwcphsM8+Ig02BjF+ErPrdVKsCfTCptw3+9
D3wjmeUTtiopYSy7js3EJzdHbr2YY/D4b/ePqnQ0dsOGjGVBfaV8uOhovagk1KkcixyUmHKw5O0P
Ka36FyjtjlOK/GB2XOrtqdcILB29Y1EVvPzi8nqWzv+Xb7d9XHCi6pM7wZGhRKpsHfSD945uuCGh
MDquQpH4xVZM/RSLzL9UyksHb1OIU8sVO5TBabczREez0KDEADU+QEIEDCE7NNX8hZQABmYVe1bv
Nde2/+6gZYcg6kn8sDqAY/+o8HzIgcYODf+8x5Byi3gLC1Sw5p6ipTZ1+tJuc4VBT+k1vouy4Coy
Br15kDVisLjPqqsiOXYut7zJukyeKrqHkwaR/hQ6xQKM/y7hLRnr3zwpIQWl23hr4Id1QbYhVz2n
N8Tqq9WApSKLFnzuJUct4VcM8zkurnF/1LNUqPfPwIyoStXnPCvf2xiR94GWLxhplkkI9MqOacYY
qJSZXFDlAb3tfkaVPAqTbP/kNUVozXR29dIW0V1/DeUm6qeB3uoWSuCHL0C3ZZixlrU5bmu77VaQ
19iLfccpQXvmlleM23HUOmM19+QxRSjSLeGh70z53Df9GsvNq5UqFROLr4mVZ51nbpUoIZ2Dveuy
rwtgbBHsZRfJDpsNWcsy3GGocQ0ksQcFvq5jfqtkmsd98/hALVtMcEGqy/QNo01b6pYNXLgLYEWX
DD+6IcIKM8x+BKB3IkkWJLKRp1YHMJcAYYa9jxSPSsjJDfdmiWaTorvkc3hym9M2HwEtFo2T6PBw
HcaB0xHekglYzVGz0qPgNoPamDhWnGTOaEHN+bOepfnMR/pu/gHVI39LLpRYvwGaRbcnyU3BxazP
GM13e5uLBURi7QCYMuni+9S3mrxWInXL/rP2z5KzI0OLJ8qd/euDgT/dlQtx1cW647xAiM5nURXW
ec413nDHrUX18jNIR1DP0rEZj2/yMFXWArouM2uCtqr7R1Zg42klfdK+iVQuNdoSRIBoHd10xCd/
2YMVltf+uneeGJ6/ZcSTTGwG2+T8W9wsLKAK95z81BS2uVy3FZRvnTb+RaUIB8/k0lJ1VsW7wq6j
mzhqmT5ObUJ/giDjO5S1jT92amB2frRZVAs92/G7IKErfSjvMSoC7ofc4MdwLR6G8w6RJkr8eZLR
g1d6mie4B51EVkuYg5ofRFEhyFyTepfZtT3qZyRrGCFGd5HmclrmGvBQaQUVdhM5sB5QYrzuz16k
AWapAs6gZZq8s82U82K/QZkQn2VNO7uLiF4nj3l9rd62B0uOe7b5lusKOnNbd2/0uiygEn4aKkCS
X4n3DnNAARn9zivc2FMZ1u0QrDRF6x00bI9+BSkkqE15hDcZNlPULkdNjwyORAdlTj7Ze5QmDehO
fBmRrLKFz5DHC+3A5+yU6rMQUQ1ENbRcnXC8kJkPTYgX6Zsthhmx8y5ZdSCTxBedoANeJiXQHflp
7cVsGyMKHgMtRGy7KailIDQSGFZ9VcGNSHfSAf8dp3Capvpm4v8cXvgC2oVu/457xrcPAhnA2Kse
iQWKgNzT9zirk5irhEiJrdyqwgw0qkRRwc+oevjW1p8fzijFv4cGhqDf+k/3nnkra+BmiWH6poRk
kLOh80etr4bUfPc5kpLlYacv+g3tjgmu0gbDXk1jDjSRVu5E0+goRDwfqYYk3EUM+3W7sn7DZEMZ
QP7CvKZIGxsg0c9lGbdcvnJjMo+LJ25Xfrvj4IGhE8gMUjCQOtHKdIJB119P299HiXQ2UDzFdXn+
aXxYUPAfBMAm7YeZMnsEtVneogSQjJjtDWQqMLrGsTJlZl4FeiVffmAcYIN0P6zdk4GVE3gk+LPE
u435YgsBSnrkkvtyVGd/FDYBI6YXBF8txw0y+tlKZwQ8yI0hB/9Diy5ccb+VKttjplKkej5ot8yM
jpmKwI5yn9RmxLOF/pV5yAI6xpmOes01lg8gqFLeXV2ruYU8JLw8VO2l8ovznAabTO7OZF2vsMzO
c3rqFbFEY4IDtPhh5Z6AW+adYTzO3CkXccynlKLlXCuJqENUFkMF21u0rBHHkMqJ/veMd0mKdPfD
fu7ZDV9r2YJE0CWED5vbYs3S99K6AYU9Wj2PhM+j9slF2MLtd3YmqkAUNhQlEzbWyDJqoMdI8MS4
3hDzbQJogEmhcC0x7oGc1fNP/oBd7kl6x+mbBgIhHrzP1c6TnKAGrdFwsIdf7ZaX4PrQAuSkjXev
bLjEKs+txGa/HVmslzKXCuWCeoYy/m5ivudXnsTRSHJBZPMyGX8djGVFqa9oDdkYons1BLrN3iBO
CgOXei9HkvVGsUeII+eL0HImBoq667nId4FewpwZK33Nxjp+UciPPpGkMLPmLfUiiFQ4lPYGmgZz
VyWTiZMH6LzBGpLM7ym3vWRg3PFrbk3+d/RvAeKAPyt5dCmVw7Y+wcyFhrmnwCg2cxh94bj9GkU2
HxK7jRjsXaMBR38R2ZXikqwhcoIaIBMZlJQLNv+ifbQzVsv4YtBPYIHF9XJDukMifJw9odb1bv5d
/QXf5AF3UrDiE5urjRjekdSjLCrJMVljsXhnERLfId44Def5X6Jbm0sHz09EGN+ntJYBbTSzu6xu
ho4dLB/Ra+KbZh8wBaGVDaU+d6NoAehqJ+gcF/EKeFPeyJMRy1gZZfnbEkDWNr11AWb74MkROaz2
2zm9OqUcUEmpL1lzrGpr3ql0IG07VAR2V8bk5fYiKdoWEUf1sdK4u0KiicHuNNjmhnCuftLGaWvC
Zb3juxLt+loz0b+aIcb3RcJdzZA90M8fv0TRNV7yg5j2ufc/gAHjWF+MIVpAm04LoQYrka6DdAZj
RqAQUJ3Xww/ZsWr+EKzvMiwlJlboKrCmIyBeuWIGnjRMFBmubB04Gxau/WB/3CjpSeQVFf6dENcn
SqsedgOOYpGIFUAFR/lIy9494ICyq6kOFBEuohqcgG+ls+THfeXigGChk9h0e+Hh43G56JmDRKHR
JBQX/EvXdmCDEzSbVAD4SL10vTiwJBv6xIlIiTiDsfxTjIMEf9PpKRSN7XjFIPd2PMFEufC2kRol
xTnq3CqjgxKnctop/8kb2N+klf9dowiCzupkjmb0dN/hwSDz6gV7Mv/vhgY97NS7zTNjgfxsCr66
2s9kDq3URgV3UlautkqZMpAL+axEsXG49LJauIIkHpBnNU76Adz8ZaFM1ayE/Ra3NjlMveEpcDLi
flvNj0/dr3QxX85RlBB5McBcuWdB4DKw2fn3JFhv2MMwHctbUxH6UULrV9AT+USTRTHpVdgYYPee
i7Z00M2v9K3h19gLGeePiYH+osHN3TYUGRsgAeL1mOpekRgKjtDPnxVbtNgRnEKjOGy49BD19TNd
ddA3CRORxFRAvF94bIUJktm1AMOlCyC1ndAu6j0xx7iyXp9t+lJUyeOSQOIxjB+otKYb0JaQtWtE
eHH5KQGrsFwaJFrlTKqO6kybpFFNyMEyU8gKauS99J6mv/NVjJvgy6mKB6HS41JKWSscmNsnHZdB
7wnvH9dBRySbrD0oz7x+EB7MyIIDZ2OZ1MWH5EDuwyFU8WXSVV8xyBuxipGiXuyu9/O2i5gErysk
T0dkJtl7LR28xCD6GNdzRLGyVgIC4uLj91GkvGl+9oPGWKJenHR8KsdTiLGKyxUT4Ihfds/7rJLX
aZTUK06oPRCgUc4FdeAzcSW3n+C2Z3V44sfFFmqR6z+7thIm1mkUMkec/6DKk+uB9tFYIQN3Te71
rOOWpJ0v+ZT7lhTLkjTFgLbGcWz8mdpXR/iUVvB9Qnk8daWzGLzGNVkG1pFhWaUioxxLxzVST2GY
k6e8DfqCX2xlgB1XzlCAQtJ7tRipQR45rD1cXokDRh0soiV+kpg71ogwfC5Pfbx2Qy9xsKekxxjM
xrbUfCYTLI95sGmMZRkjUqW+EjMZfGdr6pg8LRG+QEMuuIDCiKBKjeF+RER50Ai9Os+xp5BME9VS
ojRb6+K2NXTTkG0PygtEFmANM4SJ7TQNaH8YvnFRsY4Zl7cLVXeEA5+KHxjgQVb8LaHtNgLMzr5k
eocJ8/7vclJGnPvCZOflaXCAyuitw+Gh1Cib1lYr7pRrvHSDGGypNXnGYQcQfFH5IJYgcmmt9T6c
ZGen/jOmFnLkDXQOGrvOp9DqVFp4LRg/Mh7JX+TP50KMDbKFRFSNZh4BKmReImJqxuJD35HAzaXF
I1dTlXHjdj3onM2SgNBNSzhWPGmcKl/tT0MwT/F8/qNL3F66YuMOKG5RnsuP+RgPxcpKXhyO6lty
zV5w6XE6LaFm4iuc+0WkY1ajbV0H3o2kcC021j6G+MtlJvMd7CDvh6aqr9M9nLAxd+uaw5rGjSSi
4pvMLFcJAd2Tk6/H9ZKXpLy7MpEAuC6284OfTE42vzr9ueb7ZSzAnxcg3P2Uh0835S+GbY1zLunY
O7yF/9ky7KsArqfXdhlkvwmVfAQJmFvniUHbqkErNhW7hhtlS2lR4cIK2hLd93GItFC1WMPcdI9u
DQSjWBMFK5+kmXfVvNszyE6XHK7dCAjBZOu+uYwMKgU/vjI9gtjKU6t3nWJT0ucsz2ueBP9Bx3Vw
OfhZaLWSTLIH1S3rZKDpgEROzQE8ju+fIhUW1HhG8iHijlBFu98TyFINXCHFWgSFlxPjLcbGtNM+
kTxRDxTByLp7B4KIc8FPjKK1Mbfa4K1bSnEbRyYu0RZQYIOyqjjyeMGZxk0N2CoblYR5qCZLSZgx
Yq8HE+lR0qSCIekE7ctIU6Vdj+FyjDSuDNB9jBRVRdtk8FENL3oF73AejQFdJuT2VMQNmol0gFas
h9684aWbc5xL7HaO0EWuR3nJ5Eu3+KClUBoad9T4Q4SpIGR4coyzKTokMlbsXB62kWQ6jqhO1Qhj
G2utfx4JA45A8BsuHPUwrUvjVnlxLmNkd9/3JrRGeJz8BfdN2vOc6jV6ZrFHvf1NbxQq9K3KoYBu
qzdMcY9TUc0HRSSPHoO6sBolPOv9GWFrKdkEYU4VpMQeadFyRPTfn2SYx1l9eBTUUjuO6G4HH1aW
OkmiSjn0AjUhcwLeOnO8p25ce3IOfqUZ/LF/9DhcoR/WsloJcV/tbaxExHyLbY7wNankHDz0t+tA
aBbowNmxwhS2s2mAD1UORCckmUNGFFjzGiux4hjriBhmQHnj17vsSmRviCGeCFuOip2iftNpGeOo
4C/3gy2Q1/4XdbyvMt0cc7RpXWQ/ti1STvz1pdx+lI6oN8Zyds23vM7DoG5K15+nGIeB/5eHzqfZ
B9iZE+rrjCIwxfWV0ZVlp4VKtSLF84KEeG5Dc8BjkZ4uVzQ3NNP5JqzGNC2nHb5WjARTw6Vz1hFx
GYWCDY830sh5BcGlSIpQqXwpZdoVNb6lfiZ567UNh/MYuOT+m/VOSCya/vCgDTGNIQlDTEHDVMrI
lXvERaQiOoozpVOdkllJLH0moyK2i1XyW7d5tXbK8tBhg4P4dBU2i0vLk000CMu4DQujoWoC9msN
FmkgfOBSfU+AVsIoukS0HewxIjOkrTXq+SDfXvXfE3sjxd2WO3mjUboyn62Ry98ZML9RfYpbMTQL
x+qNdhYQQqgHjc283u8Ef3+0BUFGiAu3mjC6P2C+tpYruwtmF0wBL2rU0n8kYbFpjZfubDsSNOnN
5OG3i9tCQ6vYUk6kgNCEOBodW3GZRXslTiWXxd6UZdCM4DsQSk8S5DH1JuhLxg/9ackyqMs/1HAK
QZ0F4elmohk4/OM0AFzcVqwP9cBDmGOBn8uL0corGIWSlvmThoTiHyw51zrOklpxcG+U9QFFTTbM
uZsTVJQAbCjFKMRWt3tp8D1n+w2KwROAi/da+LjpY+lkEl/nTwujIMM/vHNAy/Ib8LUH0fpKl+dn
/j0kxpuJyZicXWy72rijnzemXC2ovGsDc5GvnmyMldi2UnEKCTX1PuADucjatSeKQYWtdnCVIouw
7nI4jiqUHwDoixkKVc9l3JHeRtoqgsUI/a/m8x7Rv09nMj9Unq1eaJdwJMrtybl+grhg4P9eIak2
fIBZKD3BVqIeOoF2xTeDPOCRhX/WiJUTH/b8eGjcuhACnc+7Ri1YbANbbNbHOKjM8p6Z08+al71T
mxo4hk+KYAbtXsCkUYK/mlHEoMo0pXP6TxdaNW4LEOdXTD6TwyakDtTkFYrK7MHVyRqGL8b662iX
wDEgWEO6INDE4jUzXomfhm2BVKROqbDG1cb/x2IDHbL4PJsZ5Bfs2S/h+Acu8VhZ3cPkV1/LcbJM
YrITM46cxdczzjn4ddNM4105S9n9RdGG2EsQf1nE8EeSKhUSKYK69gnDHy8UfjbgJS2zMULV8aMH
fVYUtTXtCwOLEL9yG+sc8y3rW8rQCHeEbOgInW0ftupEYq20kYIxKplCPFG23q0GV+OY9CGfZgZ1
kAMHKIM3hchPRSBz/YzTKNPbHdftRO8/fp4k/oDRpbGC+XLguq4Lm+NNpQY7GGtMxQ9jJlLFXbq4
tXgIzS83KHlrgjHp/yUIwuEwmiBUOpLwaYMfXLrq9CqNZUxQecjBmibwkUJ9eOFPtCtu9mZyWYJE
DcxO/Tcg3v4x3KcDMeG1sndGkb2exuGmuhYnzP5e9Od7451ZCzc1HtuCVxHclB5VayYqVtiFtqhF
24i7OOLYyVEy/IuUCgzxkwiQjjYDLi+ELkFLKHTfmYCDOewsnRv5G70RL/C/30Cb8kQwEOOpTY2e
9FM16a7z5qiTbgziOb7RZ9GpD+YXv0QvQqD+fN5xLe5p+myTjmHMubcNrK9aQhkpad2GEiAhnn3W
oqONxbPiS4OB20AP/b+2PMALzCmoV2cSVzFjwdkHIn9QBWSiyr+TVIeqG94kS4+fy0/OUyoQbEgU
ykEMWsUQRiQF9l/lb9S4+4p7H3Rwyyo6MqdK4bmnt4+JNsUs3qG7f+uyy986Foxch+80SX7XjILH
AGsyWu7RMOw9ar41UghLvL/9g0/B4IPMT5GNGneUtr7VyxIIZICW3Jfx9hAdjdIAxMQlzUMXy9OZ
S8KFe24mbS0LFFiUE5Lm5eVkXJhGPWavgEnE6MmAyHJo8hQDoU8rXYhSu9/CUQHB3MiQ9GBkJErp
Z/hxP74YQIJaQ9EzkFog5N/UApwVmhHl3zaJbVJGK5UISPY3bZdV8K5+AYPTl86ObRqyFQPGB0M7
pu1hMmaH1uOgYyUOLpXhDBYYHLPRl2aGw+QuefIxtHKDt1arcXCR4+d5Kc+ToE4TDGMOaDLiv15M
EHUg7Bye+SyUz+4SKWf6TfuofluiDu7THEAjTKgn4XDvO9ISbLht66g6WMkB4bKv/2N//8Ga4X4p
97FXPjRzHdsGtOTWDaGQh/4g/mBox2eg4/qVBsF+umXNrySsd4LMbKPbQh4bstzCfDIT9Jgn8Ox7
W65DhfNXwW3u7n0UeUaDKr8W1PWfsHQ2KagP92fcacdGGGetgLyaH5k/dt50iX6h1uzzjmI8MfkW
E1G1LKtCHWMmvNxGYc8d16GZD/yQAyGM8vvRJ/IIT4ozOGLcHenDXw7E1M4POkCJ/oIwk3IzsOMU
a9rGOYhPeXIq8vQi/Sdg2jcyr11VL6hxLLaZr302PWiS4hdn9nTYtqDsAoO76/xh8bWGqdF7fCty
IP4N7nmM4Kr5Pjx+iLjzwrHf9j14uIakwZohoJ5WwN6PwongpZ+KVi8Z3evRfa3OaHFOARrUsOBY
eSX09tnU4NfcKv1aEY+pgRBAC+FQQt3bkkk0bTHpS7ECa4FloaBU+TWOc7vyCNbXnb8banyvnnr/
j/j57jUCi+V84Qzn4AjQtZPEssq7jn96dEL1NCce9PM6nWuY/pa8gYfjV74YOCGnfLA/hqP5Xd9t
DDWvMHwR2vyM8AjWCqvqowLKWbQ7SfVRcNg/Pe3Xivdn5wIhlnuQB/wu6kicCJueugx5RdNdFiW5
YcgLsjnCeEMau8JdBNpHKcgulJ6jiBKMLT+aOzb117iEN3KSsi9nR4tirii04LCMNBBksaPp2b80
K/ZuWnnj7sgSKaqCeOwOUdIzZd+sCdlocaW0PgfZce/pTJhtTuT/jx3u6+UCZkV/vylRnLhNMOmy
ahMkdl2o0QGQFwWkA0I2nn+zpKMuqfxhK4CzlFyQXNnA0MHon9dLh2WHs6HUlQFI9JXpp/pkDABv
SmmmharKiJb8UuoGGqqHp75aEFXB2IgQ64GNK+y0yIPE8QXr7X2VJ96AyFrDTIfkpdvJR+TirUox
pBcWFOU1X6zyToYQ6aErFS0WZtDFeG3japJtkbuifteGYpUxTdfhsgGIxaahNf6BnvGPyGufYoQ4
/hxWwMPORVst2WD8QZ5emr8E6xVVY3NyjMQS/LayusX+FifBTQ+qSnOjazdd0kVlrtsDpSbtUSyY
BIUHQ7VGMkam4rcHM8CkUxigZYGoUCgRC5DwVxYzO8I7al1xdyVSbrFbZ16kq3Uh0w15g5MYoe/2
VZ032097YUr4BLo9agZlBR6QDc48NUOdIathcSerxxX9NhwlEzvBzZ005SHneIdBfknaETT6uyVD
S3SZeEqo94Iyo/fuY3wUC6tfLmw8o78H0AQoXpxzyZE4QO0xBEehJNCTFnsghLkuR6WAhjFLIGSB
+S8hDzyVMLAw+90sp94OY02gsa7c6UrtmYsj9+93fntPV4S0Bgmuazwknc2ed4JKOBL0LuYs7/cd
FntrNUCYcavcW2IXVcbeBFffv63KHN8ZatqYl6ImT0yMLV0XzReqR6Fm8J6CYfNiEF4Z1dl25fPL
EL9M3xFWA9sWtww3y9Ww9dEYTBPmlosqa8YRsBYRVESMDA2DFvJDUBaW9f3XsYIGxI9PJCJZArSM
3FeRPG9nFvN7AH1uvO+IWDbFYer3G4K4XPW0pM76h1gUyS49lXl4QqQeWlslFjiAtoV6oI/flazG
8AeEHlbj/CUxfW+rRSkWyWIM8Du3T+B1nyTdOQRJr7pyUY3xhgy+TdRpD2fuOe3UeXGEJ916fN2K
5LlGurm+e2Jd65DgBoV15Fecy7nyypqg8C42bfLQP5AQAmjGy/mMAhjuxq7cRO2dhvRmitBeVT0x
/0/nHi4ro4mvCZhpcZvoinqT1LG4GaFXF9LkeNV9nvkNlP94Ml9ezsJn+zb9bTzP/k8D5YlzJTYz
tt9UJ9/AIXuotdiLthD+2uYhvaKvnhyGBqtXahc1GdJqHZamIsmQykoZbdW9FaL3domWM5O5Bnh5
G73BWoc0z05NrrfxQwQknJYxkV+Djo8AyoMt46XxFQnYehQRRNRdSORyXMuziFrLaYkHEz99S61S
f9y0d9HjtdA787vMJITLhaPs2gOXACF+yejiTj509f0ILOO76vWZEixwdwEzO5mD0DxDKLSiOFkV
F1Cpx0i88B/7U+3UWC4DjZ83URPmdAOIuXmMqaqjOUW36R0FMNS/ROcNSto7SfLcowW9ltKOnm3i
DVhSCf/d8QbtV2XKsbTZWJhQRFA+o+YcDihBSxX6UIM/bpK2vLRQc+HfVdAAP8sd7RNp2y1eBTIt
MDaghT6OybNwEUE6CENVis1yIfY7TgQgi1D2hNQeI1ZwGQyasUZypvNrrgDyKYLAPsha0PucD3Gl
Nfq0tk5RnA29Sm8DcPg8zKvcafJZfxkcpdF0HjMzqFiferWQZAmY4S3jKjtJ/WnErZTLXBL6ZBCF
V+FRPpqIQpwct7jGsMeDYx3aiIPoSYzQB+VwtUAVpgG97N3OgOifK+ADqZFhCoJY774NvpJWmnij
e/I2XLfCgY97mziXKwVdrDe9j0SDt0b3qvH8rtlaa1n6+f5mTnrpXKHLCd3GG3Y40NRcWd6KynGi
jUN2+GATEBJBHmlOLCGlUWKMg/BQQie22Q9BEGaI+yXiP5AClPF+PjOQgP1D5ObEwZba596d/Jue
ZLEhp348g5afZwbu5tVWigjXxFQ856Lsg3jriQ6ftxVJ/M/XVjt66nSQrtP1m0UDJsO+yFH4TpBx
/YmQAkfCBMKGrr0Y0zH9sf16q0/YQf4my/DMBwZgo8d3Wo+Y6ISNa9bJDSRoWN7vxbfNmG8FeiH6
V+6KcHP9II7zymB+qiS2b1t/NtgalbYBeUTPK5+SIazp7TLup6lycsXx714uA1ogt+OM8px/g+WS
YKIJmTTrNNwQDebC4bCW7yiul1WZH+q1nVSpog5Q6U9nm5rizPNuC+xsBBj47NfAXvPK/oRbBYQZ
ZnpsmlyTMRn8YO3EtYFT8cpdk0K6RP1cizybwkMkNz3/PpiQCh3Aqr8cYrOOqGYZ4LvrsGZDZPg3
OJajHp+J0pnA5AD3IAv6O2+ODixRNEujs0VxckjnsgJXoBrQki6yg5E2Gc+sSM+U3zuh3dWeoN/5
/wvt/uREhRbasZsqR5HwFiLBe8Gvfv9iD4ZtAhQnaB8RezErhDPfaoIVwarEMyr6TNl51fgH3ZAn
IoHrSJB5AdeKX2tFzCxl0WXeAafk7jXD/STqs9l9ylxfzIakYk3V+KAveZRjdwbiNIV0gv69LqxZ
o/G8R3XCwQlZ6UDa9pE6aLrpJYT9mzI7Vu1qAuQMwwePVEv544jsnn3dKd+e4vbPKlj7HurmmrSB
EtnS0lNHBvVLxBWyqeOe97VNV+eEkNLtEqOXa5PZHhqRQnSqug2JMO5PoOVkI02rQ7pEPsil7lUQ
YY1l7SshH6XsYA4Kc36P/RhvrS9eXkiCldBGuV/GMVJzizb3XJdCloWVffF3DNb/dV6mkWqVAoKM
lIVO4pcN78zUHQr/FuZ9nEK4WBYejZHQVA21NWrKflrYmdtd5EQwI6JWC2EutbqPqKimnMUOCiow
44A+EXolmLoDMDK3X9DJYu/PCgpjYYKKT9zBS5G5jT/JNaxAr+yi1nKUurJ7O3BiP1tCuW0D46nY
KaKxifzxHqjelHaYTr7vOz4YA1ecLG3h3PrRfsdpw2WY+bIH+9c+SQ+NRpD00OtlSI8UrvThqL6E
9t6XoY5VJnaLPR7PG7oSOyV/mXqr+LobYPKylbSfgFIaG+TAzewX0kjFy4X3h71/6v6QwFYnZSW3
4GSXpFfy7ugPfPld+8qL0BWBbWHjeF/Y1M/3kaROSQb9rYJAnnM+rfTh8rhzTKsXK0Oe41O8sZR4
C3/drlGNX64J4jiF5ySfttEZXyJaaOvj9OA81v/0/ylJ5aRffY5rv2NBFV7pL0qrdGc9ECFLSe+R
rs8JLxywR0+GXzF2tqQgPMJLBgS5+df1gqR5vMJ8XOowLbQv8A44C5khetRoPHNBEiPAGRFGVeZF
4PQsuhIGieYtbsvA6eu0dFDFta5JKyHJ+WhPb9uOjZhrU4BeK71fo07dZ/KIHsOJ2Kzgp4voXa1T
rrIeWvzYcYOMA+SqLsl3pCdVRcDjlNVonYuP54bpHQAWdyceaiZBgmMRLQtxCextMAH16NE3Qc6f
IbRop8IAf6/rn/EOtp249iVA8WZvLLovQQITN9RXS3iRJCczIzv4OLQ+jZFyXUliu5I6sdepUj6e
KrotvGflKMyQZIDr1J0WuMxOzEqNsR8QXIrPBBT65Qg8T2zeaTdqhzMO2enpluIrxXFyEmaM15Ly
6CD1JLBHDRpDUq3qpyVMtOquP0d5b8TjC5VzRZHK7Ahp0UdupA/5L9uKbVYf/kFcOlXHoPYs8dly
9fs3dcr5VLYJQPTRBICBgtUav9oKcOwXDrxiabm2qdyIbg7I25kNLZGB6NvOSb9JFeo+0He0507B
7IDo4CELOkyXtcfAbMj3ZcUjxfCukCshDA3eGFejB+Jzr7De1rJ3VHILa3n6cL2bir0HAjDwzB+Q
b+26OWZLZMsUCABmRPWzbqanjQ5i5tXmTPchdX/9TT2YfS5+bs7EjTePBvXHyWLKpGBVHok0oCTD
0YnYZENT0T3Qx/xDZ7AAtx2f5MclztgGu/7lvtafKXtJDVZAMEv5jctY1Qe07xWIf3+f1Vo4lf7s
D5uHCiUP319zISS0KPNMbkDkB1cj3K0IdcgX1hWMwEZE3YMav6XIDoBHiwS271+Nfq22eCUdFqzN
VEXVMvUBiqFaRzGN+uuO4NC4+CWD+lasu5+N6Hc501FPa5yLYAPcreSEoC+DASezrRXwaTFZEUvu
q27+q51a3bfWIwko0KnxdyrbmmzaI+PdzXCRYC41WvYkbuOWm3kjBQA2Dpy1jObEL7jnTOqkpEQ8
YmaEfFrYWYomvdBuMfw9FqWHKyVN1vTUYltdGFX5zpCUyufpvik8g9Q3hIgTMSI99Sgh6flPShPe
2Dqc4ZqBnzrTb4PSn5thfVXCZ5vGVI5REYWIMczWvH7p5+0x1B6e+3SvFHWkgGC9YgSCCMb1ocrZ
lFr0/IDdRbNlqsaEac9fGkn0iKg/ThHumHkvzWU3njJyatY1l0DoqEJltHvL9wS669Cn9rWLZji5
LEdHUo1kKA85D4qHH62lbjcQkcYhHjZ48UyXUgYArDxqpqolaWEj8N25mgevSDuu1KLUztFl0P9L
nyGs/aDGO3fQu2/hHgazFHHEQMxzJ0173tn4l36YELGtU7ssUKRT2fKvUJmeZzZMHf/GQAT6Zjy1
ydH3N0oDos2PfZuWs1zyTtGnBeUQ2zqek92rUHEYMgRT3V2sW7Do2pg/UHaUrUNlZw8meLomwKNx
x7piCXQMC2/Q6h/aMVJE5irVXreDvopI6X7SiphwSwSbO4KkAEK91xh/9n8HWW/aMNxXiHgq0xpp
pfaJ9qFvbt+O2PPA4kEvZZuZKzGuz7GyToTfFkBwfRa6WhBbirY+GQaa6GipQYx3uSa7BZLvsuOO
8V8ncFCbckicE41hfZXgPGdzvzUqko4L2HxkbPQnvhTp2uMZLg5kOw/9gK0mT48z2qUs4dMepiTz
7Hf5Ll4knrxVe1Cbt197FCCicZc7Iw/Rue/llJyz0acxv9nl5yoI6aFu/4ALNyYnoN3dd8xNJGSD
Dht2X4Ely54UPQfmwH6sel5Ul+9n8Sf/UD8F3cUeVP07TNTZpWec/IdTfMMFLVufWAfm03re8+H8
G/2/cKGo3CT8A/NNvRKaL0QA3YKM7R/5ZyVidv8G/T8UMNH0q72nqF4SZdluIg/eFvcVt76iC/F9
0ClBXFv2B6TDzhTEVI3t6mCGcZCak4q54R8Xsl/poGSTBXc7/azOABOLYLI06+gM4GDPWGeqv6kZ
DAQuEbOGS9TDDuEvyJ42f6JU+Dmq9kTv1bOMgxqX1bnKZ+JrHZUYQH0zSrHZ75bSo6/38vX7oUpR
Sy4k3Ph288ib/P+Au2bXVIRmsfPMQKrNlHxZZS65uW8LvQ095Sj/wt9IFjMBAQ61JautfHrPx9+D
9L9T8B2fhfaLE0RIG0bLPWaGweJFO9WnT8XXoid7xcXg/2l4HE2zEbroZAvGbjK+vkomlMjh8ivx
Th6zxI4aUpbxKzs4i3j0Rh3s31aiHBObxWP9NMYk0eFKtnvCEsoO4GtKGZ3Tp/20wl5iUmx0tIMT
wsEjgmj9ulSkFGWIu1Y2OLomvH/cqoFhlZBb/Yi0gDNghFyjYCy2PsnkX2cOT2cEA+3mZYCAaIox
b0C4Z3UhbE3ghHHtGScVlZJy33THCZhHq1c9TMS0LkLAGbwtU/tQ+47674xIym25r9eUcGKjmx6L
g6Gq2JBmDyw/mFeDP7unzAA90Zqmd+63ENK0kaF/Xw6dZO2XUjR4T3kKedSA247Zz0zRKpZJEFBp
+wzFEuaTadh1wlJXw6qMieLO0B0/YJQDHb93IzqM35YJgmHqwUnD26mBPjzWq7dONV2ULt+WXcTf
jC514dX67kyi9EbQsIoidlKxiRIBJYcSp0yG7mx1TCy5zTbkhW375fb+ehqN2apRUHB/RJX831Xp
4wMLBXfAj7DAa1VIu2ptJhTIgYAebcw9A4LpNyJawwM8DApe6zomHuAtcldLUCpHAwVJ33QAm2yU
6PqY6HlCF3I/iHaMPt8ik3nh8z9yc+E6MGrXlAK9+hLktnCdzRC0pGByKv5OjkJ+oxO2jNgTcIgZ
BP1t+2d73YFkqTFWu9FhyTa/aTCvh/clI6IBvcE1+TTct/GtjK81GcbB/0ka3UFY6NY2rEdCdma0
VxtRORn4oRQoBv6WO1i12rqekbmYZPXZvCcNMHdwJ5PSFThV+naLPNpwxoeVuD5uUHcYKjeB1QX5
fG5ZY7hF9Q7xGHpHlA9I1r3zDARx3UQ3IzyX4K0VXECT+ESSb/AZPfrv8HGYZt6FuzWdU92E/gKK
dYmnuyt9v9t0Rvb1fu+HPby8HUmbN2uFhxOOERcZDzToGPTleXnNM2cKl1broX4p0TmrG9V5fqAS
STMHiP6BBjm/n+M4iigeuGFOzqM0Z4J7nLPKKPu8H57ySFvEYkqDZvB8z6epAf1Fy7k4tbzp/ytC
cc77M085EMFn40LhO0Rx0nOgWGl5BNGi+8L0v4Q5wbAsiZuuLSFuxnVDKyUCc73CIRxmg6JANO5c
JnTOhgFsA9Qaj7DafmJ2Kn9elkjAqNl9cMXnmzSBwatGI3Ht3RcrOKvhvyo7UVZfKWGd0qxVqSN2
EP5/Vhz3ovh8N1Zp2wajHltVFlzoSiSD5tnsUDeOlMIaovN3+qvh0yZt0/jJT+lWkum6fjYa63s9
RkP7cwwL3CngG9bPB2RxbRNJZmTgmMOUHyfUFXfM5NAXOhAsQcR0IRx/1jw+ealKtJ/ImkfnRQpE
mxj5e+LkiMaoWpNmG2tGz3gwqDz6cB02lJ/6182v+gPhA0fzpV9bd5WYeXhvicnWn0aWCHffU9KK
uqD1oJGGcJGzCRne9T6vbUKFZoZkJjRaE5Z/6vn6C8PPQJ1TMzUAJmalwNst1DNj47Xm4u6MHNYL
ZPaEfnUCBt+LNuRfj/CqOSzQFxW4/mit5qv1lTbrMTiiO6k0jXmJgzT85EFgRtZBVqnLSexbXsRm
NPwJNeIOr0vdDRJDgNWrOL7oaVAMosnEBtntHtcwP6SRgN1m67aJc9DwwmxVDB7wt/lPnTTyQkdH
JgFyTg+JtdJULleAytVSKcUv1Hy9sJXxyWRqHMt02rqsIE/BfIBlj1GiYC+a/8MVSYWy4gdpNpFb
sz1GOvwTa8vRppm//m6ic7FM6Njy3IlfUgPiZLF9eDqLmRIxmyDj2P1BYI6Y8Zh2h6+SgD0ZrxmI
aSO1IK5a9bwT2kz7wVSgV9ntWTYqNaiQieKPbtaNir9QwBKwxz2qKZu4zTQ+s+TQscb7cgRb3RRt
xLlAecR+tAwoUkuqJUXoChSTK7dOBSETRkGNL9LH/5jFw9otZ9txmqYSJNrmsOVSzhv8uYoQ/1vX
9OD9ZPiZuSDPUR0erm5YLVE6g0NBOm7owVIK9FYpaozY6H36utnQCzA99Cw33T8A9PQi9H7W2kFi
1cCBmA7KUarLIf0gxplDTEKUpdAlPPVRUQCrnVnUKBFglPVAKeHX6fX7NhghE72JOIAWZIYo1iLF
xFbCs81bJlWeLUYejqYS65fMPuT2Tze+2o4sHp0N4a3Br/itTMM1bBrKK7b16Ls/IZS9HpSRui4m
YpnBbJuhqxAnqUEjZq41Q8Zfx4oM4wwsb7BLKc66B8cZeRSb/KXbjMPPp+OKD0wNXhQ2JnUwpz4I
/ln+LGZ4u1qZ0TMjjm5+s1cxAGrhiInSGbFjXiovT+WiFjaTA4tgkun5PdC6SIJEu1UA9lYu3Kis
+r9nI2hO3mcY4HOz2/RXWWGZ/miSiMW1ilV2NWw3y/KA/zRZmeHxxGo8JZSnbrXKhGAnojtt/ggq
jfKlyxNtHgUCaoolzW/1mzNzP+YLs+MBgeCoeljBrWAieUtIILD7Q5xh61ZyB4d0/mk2V4znwLKk
7Gm2YPYL8qgkcHWkfFspqGR2dRSvNmvTaQKiMVjyh0N0hTa3HZnawGNfkdNvypWkWt+Fhw+T78S1
L7LmWyMCkoPryMilocBbz3Kp02iIT2NNQVXeuca6WNsGRiemNiEzKraykK76EHV97Wy/WAV+cEuS
p1qLQAsCB4nPwYbqIh71HHlJDxO/GkI7fYQiHShZ5huZBzFE6VxZ5dkUtXxjVfgMN+7dAzhlPq7R
uDJN002VLEwM+qLK40r2dGqRm/OMS4xHtoBv4xb2Ddjk9wT8hYWtaQRarp+inhCBS6SZsR+JiDN4
BYheqkyWq8aGJLebz8LqZ6QlTzqWQcdFUDRI/tBoNuGxSBDrVEngvpKSn2FhirRKJtzfKfxW2Zrq
WSyR0XfSAzk/iBcD1e40xBNTcg10QI3fBuaydgeHfEVGwJ7iNmQDIaojFFngH0pG7wRE3Qei1oFs
buI3NrtB6XgD0trOiB2Qc7un5bn0Z8M5TTlq/3vifhi5qIM4XGSo0x9kdYsdLwzK2rfQuyyRivVg
hmUlWx0eXz0SbfnBjiJzhPraaJuAlgY+/Fpik/dWwJlS0Txf4BVCGAW5APHKG9sYGQOOBtq0a10f
NTEgiyKEPi7VuxoiPeAraAumoqt/vC0uCinKqJcvK8baJOB0JWmq+WuEqpGvuY0OQis5PttnH9Ug
l3Qmn2fCaTryWwTuPdSG20SSkD08iM7xceKbcExvfLpuYTg3sd4ArPutgzNJgjjel0Bywq8Oz4Mx
DwiaVH4F6OYOGeEZSYPzPnNo21duRujTHZjhDA897Rlo077g0gNa77kZsOFzNC+PoGRecRbBBQXn
yPIt1ZpHjMAwtQdpKRK3eTdA+u5D2+lAt09RCaW3X2Dt+b+mfijxJ+9SV26dq5Ovicnz85Fn7md1
5Zd5wWBNZfoHBPO/IkziX5gZs7+fD6vqm5gbipqJP001JO2CZFQj46dt+gcShtENPZdfhu7mfTBG
xJlMtD/186mrL7pVJNED80j8cISMOckZelIy4ijkkEs/aCO3NGaiEPiXBMEbWab2h0iqUow/KdEo
jZfJ93ApE9ndc3FcG0cxhOCmhH23x8BbXP0J9tscORKTb32VT9vCKwhH4fpntblzEQDT6THCHG5X
mFa6eqBgwW28YQ1qESZLxIkGZycQIazC1a88CpxvFswcW48RMJDIbnHQgvtYMPkrv4vewnw1tKJl
tKGMlNnQOpQdTr2b2rvJg85ECZq7300Purcb2Xnh0IGwGpoEKnIqfDg7ogrjD886IAnAkhS2erpS
xyM9X8N/uEjWtxBkuL5Yd7USISGlLuTlVwJrFzcBSYw6CY+udX5Gr13AXpKMIrSzXKiWPh02qMDc
bbO5Woh0UOJsXs339jjk8OGLc//C7qZCd1BHu6IZa/Oz/PkvOHyyYqDl84wzV7UiXqt+ozbMLHfB
AEkt7VeisG3ci0lQdPpTu3aZCNJ2qYqZ9R6OfoqSasIXvQT84CUKA+/7hEhU4rwelMrq1I/OuHqK
nPC2VQD8idJD4vwgV8ZA56zEtnAJFNHHXGyHhLZBv4QI1USReCah6W12A4AnAtEiWSr71QTOS65E
8ZevO7jdwsYXn0rHXsHYpmz6kb0HV6k56+f8GUCYAYgpPLhqVHlm6Sqr1wRib1sNAKtXQbTBKozI
DSdNe+aKlu1B3ZcSd9WP6rrwF6Vblyx39zSbhKdxginIiic202guXU1tCe3ZFM6Lx72xTzsVUzkk
+to+2CQFaaVv4cg6NXU/DHjqWpOb/qzQoDAyGvqoXEGD6FSDMcCeNeNU/SZ5jGP1ky0dGVTovVhh
2mqeTOkPm2h/aIuJRL6m6kjJXwXWeeuxxBDr95U+cjGyGm+9GvfkV/kj07AWxCYb6JTbeafgdQO6
seMhB4L73X4jZImuAYOwEZfWtCIOgxNvPq8+7avZ1h1M6gequDKr0tufnUZKZsBt98FnbLDb/8OV
++WKeJfJwNRu4Y3wKWIzDCKQY0w5+oTGLoufls66Uyhplv89wshaMYizpFgvLQc9fPAX3JmL1d5w
V8VqRGZ+s6/s0/TQGrF1zRhxgoLRaTALGqPJqiuDoPMlOV2Qtta+CgNFmHr4P/m7/ws4L6ViyMDP
9YkafGnu1i2rB99mJmpMzftTlj0wEIw9xGQ3kehlO9zYt+f6+lmXy4eJfstyAGIT+eS94bzGJNVS
XpHAn7GcHuObQ0WUHoclmekhWmXHtrxbM8Ka9I2VeQjNXgDxyMShRVOkpNe3U2Ft9JTsqSw19BcO
6XcJnI1sB9+FI3hRvVoWXv3ij6vH6qZlJIEkhnkM9utxEwEXR343IN1hX2k7Pvt8FGu0qyaFQkHb
Ioi2hPFqXbU9hx6XWzJL2/Rb42dx0BUF/5mBt0srFAwGKeQbMx1EbDGnU4Rxwi2crRj6kqqbzkk6
3720IeWiakZkITXbcmnDqv2MFZcwSQj24TspozLl5P6zIKabr2m9Q0XgI2ijgIyPUvAQCxFmCV7T
ZCf523c7ialhACw5f0SPjxn6Ck7BZEIZx3gpv2aNP3MRR1JX9ll3yEXXiWEfSMdP8idFp6/4VduX
3PdNF35Ox4QQ5T4w5ktjNJvoJyUqLe6is5saKt75ZSkdFP/tYPiwTDaaQ6rij8OF0+XYExUqclXY
Y/6kqr744wrLjqBdvH0vgIYKdlSaIPZ/AL+3y0CItNcKO6YCEsLYrhanP6kweyh5EFCrS9bNbG0M
lR3lB8gxOVqa2P8yMgSS7romVN7N4grVnV0N2wRg5kAk9fILqRUk0/D2XtbdbGPoYrOeY+v/o8B3
cLMGqB4u3VjwsaTU6e9uIDNYrk+ecg6E8SzgivLlA6AK4TrSkoR0ZF/q8UGkxNptrGwoaK5+sPMI
NzWmr8PD4YpVI+cbpmexuaXg/5ZSECDwjGbi/eWNoVYch87iQiBpGdIeRlPnTokKFBQZPkDXhYWG
xzD/EH2PJNj3rl8kWWbw5/qhvSprmcDlpHtVHyYuPywj2+Yh88FYw9amfucfIIwaNeSl4MShycl5
1OHJOG07cKUTbRh4/357Yrl0S1KNBisCB8sTM3gpZXaJ086zR4I/ZBu2hu+ewrZ7aObbA/hXQB94
Gi5TSXrudg02gVAbgETpG71LqJPsYP9C5tKsvjz9OQYzYRQc7JOSWSbz+S0iUv9n5leuCcW99Y9k
feHhRPGlWtVnFvN2QrcsHt5f0i0JSevDJHU1fAUkrVUApm+xXzzRbfjwHXkik+FLaOQXESxQjBMJ
rG8wMOMtKfFkXRk+4DQqy8Efk6VIYYtoR6fpiu6rph18OruRVjQvRqTVsX45gb3xQWwsCp4t2kNC
VjbJHTIplqZ6LTEhXs40y/pkpSkCQG2wBaTfIAwL7FedGQJIP3YhoO4xlaX7rnXzCIHWxb76eR9J
wUqRp7NhmW6K5ZeAWrlISzJKwqFgUX97PghvK2Gc9rgSvYkxrcXfOC7FTOURqKfdjfRzVz5kvRyP
uwd+5N6rAoJ+d9Jj3GpHiuGCosSmxYbyFHAhCJmpfc7llQkFHHcUQJ12T/7rzCNC175bjybjmIme
EFE++k/XVKhN9qvoMJMI2YP8BZ3dlT55rTY2G3lTeJIARmlV++HortJajAdh+AcpnH9X7+4mhSeI
GczzodG2/+OWQhjw1bes7eTvs8oArDvwPV0RuL7HZJ2hKJ967oOe84X2jMZROtDaLvbGXuPHdvvg
yZPw2S6omt26/hRoLBu8iV95tppISfqOqcYqHA/je32ymYs9rW+Z2JhwBkgh1NFU8WslvyCVVTFY
ewCfeA0ZsEyPn3SPtdwxgv1ytKSwFq4Dbzo5zih69PPlPR+orpku1OdCt9YSt6+4NktgCZkwvYac
Kd9l6IkuVmiNtI2usJ+t0SFOmBgKHb/N+I7EGS/KDZyFtIf93EdN56Cz2LSXXV8V+6deGSTCT3Sc
s/Y+5KBxX14GqLhkTB+VTQ6dGZqi71zEpV7En2jFqV6pleeQBvr5Ml1vBokEMBB4a/s1QeGBogxK
F47W8frqUTp3+woz2HJSew+8weGgocnA4iGeZ5GZyiN9sPNacuH7Be/4ZoWF/TSvy4r9O6/IhW8s
0ikFxGsOICjwQKl6K+BLrscGtrP3QK5OVkSUmjQbRJAd8FG+Nt/QzoWc52yuEOVOlIFqUy+JEyMW
y8+5+uWALSe+aQSynDYB82d3NNv+qF30IQw4UcBcpc7U0GYTmF5puuhoNxFe5kONsSljROVMGS14
3Ee8KBk7q3ZMzSNX1yBym//fF4rUA+PDth99Elqq50OJ2dIIJRGZ64sK8PsjPmEDMsuxc20a7x7g
YFhC75a4ufGXAOxXloUurj9Xwt9DhAw4Y22Z1mJcAJrUdLgzHgFRgMUP33cn65HPBgvS0LkjUfJ7
qg9MNMAgTN+XiouX718EQ3dkCuWejwxgAuwK+dqS+KrQq9Exua/zGRmUX6CWSVS9Veo9rwc9wzff
2ghHaS1Whfy3NouQUu0EaubL9DH1B23a19O4usFPdDkBPhPNZsAPFAtsMSlbF6Xn/XjXFmG2uCqS
tzMnzR26n6hTtJ9PfkyN+OnHGPgzVFJa6JJUTRaihIv2PIihVe3Q/XfffXK8RKYn8TnOqW0vIkA2
xiNjVIuBJF8dGU85q4O1ECWs+Pdj5bBfRm1sv/iDXC90/mcGrDeNPkPD+BYAGXLregMfuHR2YNi3
3akOmhcKyq7fk0wYIV687yVg8uoD5aNcCpMSZA3ULQY8bs9thSbz/pTfoKnNAIMaI1ZsgcXMU2xi
Z+zLaFSXER/oX75qszlFnhN/SwSxT4Xs4MZvv0FtGVAgaiMeqU6FxJKDXxt7aT0Gp5icg6Im4ie1
XIu0BWLuB4XeR/LIlav7320g0O7PwdeIiJZLuu8bzxComiWScPFk+crWWk+B8bOKlweTry/iO/RX
iPxPLz3yqMqsmjKRsMu/9qrcSO8FlA6z3SccHn1T7f+Wi8NIyBgWB9HJFXQXJRyuZmrusaI43G7+
FEFstTRfAwLUXYDFlQIB/ZcvmVCCkrqxxZsZS5qbPN42T9nRN8Q/2ixFrT0i7ez3ibxZtbGM8pFK
ARCnZjMU81srHAh2w4yCb2oqd2XzWpRFvy3ELN8K6iXVZybIVVAHADIuI4xuv3DotJsAc5cK5LKd
r4iUdHKnOgD5WuPCmYsWNsO+31tDMsQxrejX/VP8/ai3nfQ03A4/r268qPRlAyvhu3mIULFxHGmh
k9lIDUU0Y2ok9/RpoilGrA5g6g++7dZncWpABEHg6Ofqkkvhh0I3PTp1UVfJdJ4ZoJcM3KrgIepf
cHSLz/+yJn+vU+Qfjk5kzc9JtdKRBbMOLxSUP84LKWh9TPG4LSq9fTxeIH0BozWRfnEFTP6EbPUP
ZTWKNr4lvFEth7+Ltwdd/fz4O7CKtJEGe+N75SrvP4QQKGua6fXQ6QYG04wuFq973Us54QKjEtvY
QrHCJkQdGP6zx8jdFaVh78v4oyj6ugHqjtDZQJZadlma33ztb90Q5NEc+ixjSZoymxI3cX1WhaD0
ORgQ9Dicy4V2FxDDDPkmOUWTgj0nd8oIcLafcXyaIxyZj/bS6QOnw85keCLV5mxNi1jPXP8jTFer
/+w5/t1bMpqSAnKMc0TfVLgBZimiwlprfg5Owzxgd5hMEaHjFDa8rk8FcyFciu+lhsVEXeDe3MaV
c4KPiNfVV9WxxPIrwg40hg4Ag+bKBmokF7JhwKoBCVIvuGsdYxKQzWHe3DLLpuRAz/bIUyiG9MQH
qiFF71T51KxtpwJUziZRrYMIJr9fXIqDCUYjb0n8IqYvH71yaIT58CvnycacLpfT+PRPE/3jEGB4
12NF/hy5NfNOKB5B48rxv5niudQYJEEVNtIM21obJYB3gFWJbqu0nYylWetEXTDLBMUCCtYy+KXn
573rSejhUXIhCldaevXXkuFFzNYPdQ0pf2meEcKfIVo5ba9vf0T1rMTpmfgcErjEkic5HIWkQ+U9
yXiXl174P1AMDGLMFNibPJ8M6gsdFsKghPR/cRoeA/ZbYa87l5z5uWQsteqTS9XiZIasogquUiSY
HG4uokS+ITnnC2itbdRtceilOyd2NxZIMNGOLjaLK+C+W8sTi2PuAIzFtqAvojOmuMaRe/4y4tCK
TOG3WhRPKm9OTfm4+E2Q77C7AXdjxY+YVdIw0j2c47PKyCtQhe78ixPtrCGMeytRV2h+AyNoF2u/
xFb/vSN9Pwdyyf3P86AtudU6lndlTpRN77+vECsX49mKWLdKuIAajXk//vREXW3Fnmd0X2mQvKRS
dW7WPj6vkCJOflbTIta1PfWF1E2DvLBNQh1JP0MegnUAERuHigDj8/ZW2ykU83nteMFiHoGTOcqb
ujlWHqf8eo96ptFwn5OeCf++7X3oF0oeLzmQH3mb2211wf/AHSwd9OcjO+8SCTzPoYJKRszmrYFI
xPTfene6TM0vtLHK4hxvTohFXFeo6/TJU5B2QSfA3J5I7I1/umizlgIxZAgzuUiPcYGA0PQIasvZ
QQOe1Fy807PPZrtBt9wtX56wWK3u0H7DNvKMPMPp9ESDHK4/NRuEnfEDxcP+oPeBAh3U+l1aDOyi
WXz4E2oRU56MwQzskkIMtmIHNsw8oqeH9f8CBM6kIDzCiqnv4Mp/h2Fs40J5IE9AldvLHprlGI/C
vqaNN3em53dh9kobXM1kYBg2NmMHb4apAE8DPMVObi50ZvD9axXkuI6h3TKNAhrDmZd/4raSORSd
QeuQNt2cU7c8SdH8YYCTCX0BYNJruscRHWjU/o8G4VHE38QrMp8FTuCJih1QGYtKJU8b5jBbt85P
jVHhoeW+ilNCtNp02F1/EkfoMEX3VCVfcKtwMozKGdPRh5OkwCS9wfYh0oNqs9ww8fJPN7xrTZMl
xGZ5SqSzzpAfmguq/PjL/k8YFiJLZQlVwsW7Syc2fGbYMwegSadsE0WRxb4JMroj/+rshwhHktXz
Z4sqkSnmG+VJ0sRWMWSF66h4l1vMuG3OI/MTrw/IA2fQEAh2hopbKeh4ramJzUpUlf47ZlJ0pDBr
O4ShuQiLTuGYgWlOSMel3hslBulA4Hk0ZNapQkI3Qxdp+hokb83buSCmuPlYDdu386aUJdtnN/nx
m/bHNOWh9TgqeGBsTR8mnqNXrjS3othJJTjBlQoBgPID1Hr7QR/04j01K/D4P6y4jorLejV1Y+E7
No1bVO3wOmmyKnZIBDBoXJfWlZcspiy1UxKSGYst5XwvKdOw5+wqhV6HaQ8s5mfv4v51imy58Tk8
YrIB545ENP1s6thxbubgT4KV+to1pQO/m5EDi5sBtmq2suTPClrFawmZ433yJwDMEga9gKSZ9SxZ
9HZ/EtRgjGW1fi6UeluaGebb/FR3M0DTT8kaluYfhyb83ZiW725kgU0yJxvVQKEHvvRgjheiWbiY
tX0zCCOUgrIGGGa/hzsQYG+uAfgQuRytEc0G/RYbBcENgroNSHO3Wnue+S5lomSGO/IHf/3EqMVj
kO+7pf51nZxoT6ES6CbJKUq9JeS3xfL9UxuGMq2jv0jOoQ060ByaOZAfTz8BsUOTaIIbwBI9kZc3
pTpKuwq1k8IPcmTcKwzcWWqbQ6Who+luOksE+7GPQBdUcj/1qKXfYKEbYEcceqa3FZafdD3L1jG9
r+VD+isrnmMyf7LYOmwI9Jw8Klgfh+uyy8CBYBzRtiW3nUgEvP5FUz5EIPzZHkL5EGbWLnTYhknp
THdlDlyR3SbtDM3SPXmc5QAGWettqybfkGLQCUJk9lR/Xyhb6uF8PgGGPHVH9PKMEu0QZjAdXCNh
D+OE/K+DI6Gv+HdAdQEGk22qSTlcW4Eqxq3zYoxVHsSPnch71R4J4scClWMmAGrky+/zVEovzYJK
BBi5P5G1B2WnmcNoLlfb967Zf52iqrVaK5iaafYlGkujgfypoYdMsvJ+54mnxiIZEqKDRT9EvVDs
OBN51CrI+r5SSAglUOyeQdGKO2HXkIC2RIRTW+C6JIOCueDp+6u/6RP/fvUP1XtyGt1UouhU9gxv
/mIHkFywRgcnXaN+U/CFaWQxL2cWH/kddkL2hjb0q5mq1zNu46JQEeuS0JIQwNx6a9+qrB+osuHp
DUL1fFOcp/kHp7omKAOZgoDTPc/q9j9ejO/9zhDfXibYbLvPN1GhvYRkZJrIzEts3ADWfPRYQlhh
pvTyU3S5Z1vOaiHBuX0JMY/AqpDqXX0ud/E7zKteo90J2PY2FRHkNFu846XTA1Qwh+Ek4T5h6w1b
14FWbcjWwIGdoeHFwQg5kIzF+dro0SvT5y2+Guww9R2dU2pGk77YjmM864i/ePlNCL7GT9UuIc7d
3ECqVquF5DkXAdBT8d+6ISN68TcaQ2b7G15qMSL1IR1HsS7bSaDV9eNJLnfzmp++ESclymV/Oy+h
51nRpJ7z90cGcBK8qJ8RObgSIS22qaEPoGh+BV3iBereIpSgPl2RimSNBCjKAiN6OdaroW/13quK
2mYGoVaSwDB4SuJt+8N5pRwB6zGHNXvL6wk4s3TwYL8wDhTextNqgrPPLBCRxXJX0g4V80BDEQVB
WK5ju4/1Ainxld1TjV8VSoDjN+jBT5stFJJF5xbZORAzx7wtoKJogLyz32kYegmTm6acg8zhO/op
qpY3cNxVxcwNDM6MJQnFdIjfRsP6T/6n+H1N75jlYWSRWVSEOfLTRG1YmVOmYwOSdj0sIqPkWi0k
5An5nk+7W1DKpIv+XU4NT2vfSeDSWk9Pe4tkmKchUwvgLUfzGFBj+oR3Yx+f/VPxVdbPZqeHqMWc
3cDUlO/mut5h4ONKMAQxuSxb/jqs2bOvyNy9YMbDdF0EP37QrhgDMM/d1+M5/mjp5SEMV0JaPi8N
XX/BEiZ8nXitZlrcMF5n/m+G3Ux1hTo50oM0fQbuF3G29wrFBVMHqoemM8CjdzCpTBwzE9Zndr3f
tQfLkblbzpCDGU1+JLp1EsCKOPKeMxhCPKWT5w4ywHPypc/meZD7Ukl0m/FNZY5/RoQ6zq7hOOdm
/RM1H2Zcy8kNdtTRHi+3sxNjyyFrKTmmG1kMIYZKajroMGk5vq56oD0cQgrPi1OHdbo+zDvxAMAO
2nKQfbsoNx5/5t653MLLXwbQYXBWI7/y59ZvOtOiRw5HIwJLtFkJjOr8gCPFeIGS+PQ9PF/Hj7on
BOrPvpSyAy8OQDrIGsQLLTGDBhPOl6QBLPyXmUsjYi1/wCDBdcIMnSys/k8dlIFlfZxOgYhNnqD3
5YukDMAax4ObUMmBxjio8rK9oeEZThwQTYP5iQYFEmP/oWB3Y67keGJKm3qai3HHg52+c+2A4Kpa
DHiRiTC/GYHl4ACLjhwpBTvIGHsZ1RaENzOUai7o9wpjJRsxLob7sypIf7hcP/l6fDkh2FCJwZWB
8qDYIuL8zM5HCdurUMpYUsCfw6hIziWkIfA8tBufFhJrtAlZ1vVlWV/UAxjHwFXSC+P3fwBKVywv
gVanAegIbIZHxF/XyIxG10KzJoOsOsVwjwhZNEmg/ovYhWQdnln7TTi4clcGHwC51rsBhDaXRT15
A7N2YAcVAu+6Y9qBq4+A+dUvXnIUBnqB7TcMGVoh6tLSdhIvqTzoWZnbqgsDBf5Rpx0MSc9nBdSA
M9U3Ee07DD2PyisPJTPs+vuQPGQOQILAJpF0Po7BwvsD5r8Zx34lklYoRUZNS4yyT0wmlK7J38gF
bSLFudzVt9Ayy4EYFyPJxXL2/hGCudN/f3TmlPLHLRXdgacHZVcauO8x6WMGt5lCZRTPvQm6/Pu4
wZOhS4qOmS8e0Xpp2Gub5/7MAP9APIPqSHBmYieZ6QBDS3pE8SfdWCXhqCdvvLh9NBHE9SeV842Q
ieex7c8dNnRVOqv9A5qQNslBuWUFssiDsudUsByq3OlolhnZCz1/cx6hXRHIN6hkhndY5IKh4EYn
GfDGI3D8K5yzAaPNeQTwwnUhRYfr8s2IMSInRtywMg1PNTv8ez04kKJgIVyFzuK9nuqpYloLvZVD
nxuHoRibSXRC3632Cd4xiXuyvLKyJuaFAtDuY4tpuG7BANBwYgo6CDAxi2Q+tRQzgkfg+Ze7wFMd
cNU4rIGN6Tg78OdN7p/kq9/XMHkOQp61nUPvVC8P1Vg4xMOsUjC0Vd26mr7Bh9/xw3ZyzYpOYZ+m
wC6nFPfZPkeB6e3br0eWc0CTJzP6Z+5CPxkfS17z5N8ipz0FinxO/mECBtGu/wFvzuZFS4lAV/I9
d2Fh0KbjGh4TbHjNOj7mbQwJZZahDFwnVROuIbyCv94vfGGo0RQ/BcoZPwbWKn8Y7zUUQsZApWvl
T++NaJkx4l30+pvC5rMoMNI51RRumbC7DbuXhle4sI1FfhXmbLq5TBvwm6ovI6hUPvqlp0WEAv39
X7kQyaJK5jq9njlQWO4Q0BEkWx34UUWgiHnB1Kf0ClrgWA7e5fLSbmAvPuvEQh0Xd3CyVM9XgbuM
Xn+fWV/Q9UnM/fpFv0btay935M9Syc9NMrapCSzjuk7ydrT1cDBHjIZsHINoMfRCsykxV6d5j5Df
Nr47S+vMulBj7PbbegYqweiqizgjW4O+dcPnLFpXvhBFFA3dUIsx/3GhUAtnR/xaxNQSomAkq7oO
zjPSRiV5AtnP3Uf+Z4j3k8QGGVFgayQRrEClGogwsoDSLuFRSFaRXaJfGRCb7x3ni/MR46xPqm+C
r1jL3/yJu/IpfyYBQZOfSpSaGE8tiXY4+KbuxGBXV8cjQmBOsxCtX2SkoT8ikCe8qE70RBy2/eBM
ApmUKEYB8Nb+EuM4XSC1MpoPPvqqcO9/kolW7V9AQH9R43wKmS90eYn+hc9sCMcBaXKzSInB4HPq
cho/Qk+LdekoBgNOyejlg9djrEs1wmbIqTB7547V0sduGdfvp2uMKzE4m+TSVfa6pgfjqpWIkX6P
zHf3hAPvkOkSkppukeVJks2YcgyIzEYyvLb7pV0w49+2uZQfUvZ6/yd1qoqxaXFVVwYcE/KMWMan
Ga/+vCmLIHwcApe21BWBkhOZwV3+fpjTzTRcrNfdrdkrPFxvitTaqGXpUIvKsNwEafn4WqKbtRxA
9CRjJyKof6AZbplNQk+p1Z8FyI0U1bstA8ib1THhFVQOFYmA1oNeGFG3O5bySPs45zO6+dGz7KF4
+rE66O/CBmojiJ9rmjQtUbIvFNHqyghs2sGn3LvnIh4yDDYo+DvnvYpZKGFbyR8VvPZ8agPV4Tlx
E+qbjqwGMlR4tDEPksZiD0Q+7Yxqz2DuhLb3LuRf4jS2OTAvN/kaSgKAHbTSjteQ3Zcvy/N2dl4L
np0Xhw9kP2WdGfGUKk10bCKE+lP/7OiDbASC7n7DLUbpqWQKoRPeU2DbdrZJPoet+U3ekyCQ5jOx
laZQM2xzkPywfCE5TwX/mq+7xnEl/NX7YUTWwJ/A9B/iR9VIP4nWkDEDdDlm+ZlN35+xnXMgwVue
1zQE6CvBqlfaah2kPzWm9gR29LWB8VWsvX8e35yyikQfCpJkn7ZF5MooEfcG5pNysM0sFKLMz/uP
kwzfdo18OkMZ+ecy5cQSpwtwNk7nNGZW1WOmInAKiWNpPuTCluEEoPN4eONs0PfnZrdKISD/xKzz
F7Qd4t0v/npljyZOsdOJN0wVZfRfbezBDq88grPfI292P/7ima1TnwuJg7wmmjDYgX/1gIYWxX8E
/YRxtm+CVza//i/EAsmGZshN3yfQBhmXWNhjGK+zYm9Vz9XIBDX91ZfOsYXLUT7Id4QUuTTqub08
/iioMi2yPPCA6pFCnzsJgCo286Ggiwj/X4Thap72U9oMsLnYQQL9ZZJ9I+b+srnc45limxy0hr+7
N0Nh/EkWimUTdh6qJhlCbXGwlXZYwSLzrEkYeQnrdne9HkCld3qptmrIXHsvb48WWEKmTwKhkilL
XOAXEf48Y3vK0ptW7+iJicTb3ljQ8lIqo4cGWT/WEqWt3RAWR6V9mULDZEzWHkqCkCu1NPGfJYer
svo5LTnm1ru6om6uC2oy2dVo3dpUPFeL08Lf4c3RFZEboTULis1mpSnsmXDgu5rOpsH9TJ51R/Vw
8oHN5efvwVL38CPt5Lki4NTMl37FqIOQxf0NM0ghc8i2YQLbYqr03zZdQVbNDp+fZbnwDLebionJ
Fi+K8BjIgb7S0LWOeI34Xl8P291/9LhxB93kup2xfoV8jgUaeAju6yYE7Wzsv6U5jtdAP4+EgCx5
P/OVsxjQirdz0FsMPozM+4TEEcaggSURj6XwKjAYaEmwEmv/dndZkdjCtgHOUhOrWTfoVjxhhoID
k7HGh13IUgHvnPvw/HAd8Gjd/LdGACd0BC4HBOxoJKykbbUgixCrpV5N0b23JiKUk7/Sv4oLcREN
QOPw0FPksAKvYbtlD/eTMGhgyNg5LwyCgolDhOIqO4HS7EeiIDM4uWLHeCoKIeXm72eJRbZ8uJoY
MIUOiXtcfqrVr2Ov7EAWr81ZVgfULhvPIBNf2bwDlX3lTaURP2wh0agPb5+blRQEPBpcc/eoqlyU
kHNuP7Sioq2uky2xR0P/InfDwuNSnsIg7rgcVOPo0Yr9W/TzjC9rY/pWURXqJJXTFCWEdq3ZWL38
D0Td9rM+2+UfaWuQAbAjxWt98xG+qAftkOBJAFrlffz04LnFRKhSQP9poZ2NPsVJUnfgkBz7H0No
S2OPK4jVPGNMJNQA0XgK67UEM6xalCQYfg3ludgepJJm+IBnWdyRrNpo+VkwFFj8g1NgGz1WOsa7
ACMUiIYZ2k2N9sXlwLSQ5JPACtVALUXVKAqCewO49U0Bbmp+Ainr6hsnTEwlr8dkDvFcNwI85DpO
fdJhqK/imCyHia4SzfEWmfC3dsQ09rUaGYGH9JQaxqEOpiXu5zZQJ0QzyfZBnz1rK2P6ngu91SMx
DLhzW3tUvuGIAdF2HzPXPG8FoMqNXAkT9HT4Ra/taZCD69b45QtQEQOw/4XA6NZ6CxlmeSlIto16
6Njk8lb60xUKS/qiNUL7ZHHyQTx6226eo1SljVJt2dd5MjqrA/+W9QE+wyHPDr644JEFJnEkiDNV
IrF2EZvWRQSwF//TeOo0Mlkg8H+Sn2eHJunFgXM9rQHBei04n2Rx5PQN+6CCaF90AaaOVJWWrO89
xIqW5URR7Xq41dyU3CfwsnDQH69kiHvOvIy+kHf1dUPaLHt6TCmfmds2gytPrXV8lhuC6fBgg5mj
LMtK4VaRX06k+nh6+2ev8VdTD316F0Iilk2NTLk1LjZWxIAcwFWC59bbXRkJ4OJbFx8n8ZcbN0Di
psCgQj5xVBxDzg5OLGCTbQl8e8LA78ChAhrTRMqo/Hz8P+YeEevR3FqwkCNyIOCF8e7AmLYVsgXB
558PTP+2BjomPPmYJ+FApciJSuvNYyuP69XFqB7+hv/shY4TNrfzwLNfLkxl6tf5KAbI1hg02aHN
C6A+S0GpYNpQAzmoqyu3v1hKiCEwxVhppnp5H3Rc5/H1Lkbajji0ZpSpe9pGnv5cLevbERncTlrJ
/Yx04zScMup9Augmr/5PUK7axMFed5AoqMJ9Kbh7bfQTHEhxUI0ozUsx4Ar94VUcd0uaiEe7ceuK
lZ/zd0n0g6NaBy9IVM2Z2FhDUmuZkuWPTNOyaUZLxIx8+P/G7vppztbo0pHL2loQ7fZOl1U7KHjI
jI6xv3BPsXTfxUoQ72yZxGtKx9sGShBPuIyOlXWNJ/3/Q41perw0CcygtCU15x0Vxqt0Ftugga4o
TIc8Knyc59KEjAejWHHtQVT8EdgAJNQlc4dTewGNSMqYLXiDl2z2WQYlBkKmO92Tmp0HHzh82kvx
9LdND8Zij0HCTL7CoGBYCfD3IjofCFXiu0QwlqW4qqPJ5uT3ASL2xMGHx2gme96OMxY81oBCqlmg
gPc+MY8jQ56Qwu6+aIYgbB146BMrsciXGVF4iLNyHuzzfgCELoDbcCQ8miXIdo2oEQ4NRiqqnwQa
i+RRwRThat8xxWgpvUoiFdXHGhTVu7ZqloYNOwjHYGHROAGgCsaRmq9Oc0qL/wRP3tucZ3HbpWTW
gEnlfHexL3JmwvvbkCmDw6pZX97aUIK9BJmNjUbMvT4JC1sdqqgRiD/XkIPcwmUGGzn32L2yd7DB
RmbzgOsX/F2hMGkvfbrM737OjHE/y6OWXZ22AfPP3XngOWwPbrlNjWt+EnXrrwiDtngDVyBimoSt
gi7szBDkDu5NMNQTda7irHdNHqweNTSTAapgrSolw4Y5sMrh7D36LVnwjSPTv2f3T0GhLPK9qTZN
5GGmMtz6G2XtzuGFv2hDWROJ0ey0t04Q0gPJg6vRlx8AYTefS4wWqeC6DJJU93DPdUa5fpPVdlkD
bOEcAQZA39Vx9ZnKMnGKwENK6W5aLHJyl+JlBVR+voNvQKS8hMVgYvtllxdS54pAIB61QOEaXZm4
3agrdy+QjtI2tBFerwHW4th3Q0uUYy19c5b7cB3QU3hZZBlSFJAS0ld8kdOwgr7j4yyCKxkk05C1
BMa9oYFvVx790/qzdeTR2X118BVlpFdmR52rOvYsih7lrVVyZsgEvZ951YQcUxNoz7gszY0H4Qbn
qc4wEyrH9QkQ7rkj4F9Ezc5iVcknRoucdZrY6NX/sr+ztQfJIH/i+VraRrxUMsO4TTxB0SA9u3na
xMgcONmSfJ1mnKMvihOwv/vwnZPe6SXWDy/Sr0fuiTtaGoswCiaN/PfXzYl4I4mb49OdVBZps6XD
5y5v+I7RtrHZNGrIA4EMaQ2QeeDSOWDqoBflgk0vQY68RXUt3tshca4VLQQ1lO/iiwQIAUKqQh19
D0sDI3HnA3+37ndlLh3aKrsfZJfWNRsP4x7IYq/++LBNgB9i7R1Ph2ZSGVTq8cmT+jcghiSquFIb
rL2yRzxzk8pXHsNfye2wTWE2t+e2JazpKWLrsEm/e1DfDRMZLWIbg5Ci+1ywJGgxe+BaveFQ5YUx
x8BKzCEoM2Syuxf5GvUYv5VvN27tfM9Z7n763sKcxuDoKN4V0yOrDXzv7/dAex9/+SNFoO+mJg9X
0KgEzLEagEY2wAiX+Hnoyx9Rb0A+MuNuZQJbYrVpc0ASHYhSN06yjYpOj/R+msnqgBqaihIdOQXf
+6Mghbh7QNf7gtctvvvFXRsHqayks/zVyuDVqzI7/qlxa0pKZAm/D8iH48L/0THRP0YhNu3fCwvG
EsRQSLdS1C0+XsGUlRHxM2VIoqNdT02kj49Cz/E6r7Z3vqEtZ4VOWFUNZnlc2DMRLRd08pzcvFbb
j1b1v/BtcN7sSUFduFyXThJifZOIBTp4/I+d4tdOoKTls0RqT+Uv9eYRW0MgquX+uWv1EqiXA/Jv
dovxdnPrfXbjmD0mgBGw+V4a/w62qrtSqVUqR93F3gdYELFbQwnvaiPO/CH/PbakspjAecc7gUW9
naOcb3GFHKcTG4lhHfsmD5BY08tcUkg+vIKVAlrYoqmTFgm3bU2TunQMwu+klxK/oA478FQ2LvBC
/q94EXzk61taPr2a7BS5VC/OXytRruF7EYdusYq7AhRd5gps4jEEAsAPVZ8PmgX3TK4vax32qoBW
920+GdpAs5t1J59BvT8+uCEKKqXwHy75/I3jeRlyKYuKq3A2eIdsuBk4Y6WOmWYVP3DRh5qF0vUR
zWzX2ovt8j8nLJqhLASB1sIl4U4iP8EyqFQjB7JZpKnbd/E4WZ1KVplTuA55YviKLhUc3+HBNaj3
pAVfCn05Rbtj2aCZgKvZMRIcMduyhFaczS8Y3AFHiQqEcGMwZtideJwP0m7WhSRfnr9/k6Dv9OwS
GK4VlwKNgxge5rgYWBc1oIjA1QB/gBkwcywd8RmhWAxo1FULv4MSdZ0TXAU4FgT53idzIUVASJd/
EkR6fAmo7D8OACSK5IO641+TQiTaSfJS/6BE62BXw2ahHnVzerm6Sg0LBVfPl66HTe5/FAuHqJMc
IaS1+7Yt9SmI6RmJhCcmKkuEQSQhV9Lp+vzBpbbE6RnMrRkWQYY97MDswyI51kzMQ+hjUsBJb4V6
OEhTIxT5OM5PEuP/6L9uVdr/QWYWRkDt5RHWhRYfBuc74J4bOcOdi9dggYh6G7mKxQ+DfpVyJb6O
OkjFnzHIJqgQiJ6DFezNgD8Rss9gKkkAtuHSBxJ3lD+5xz1Rc9St/1yQCUpnFoERaz5eyP8EB/I2
zgNtleW90UYxD9uwjSHU81yTUbwqcBL8vQuMc2qnqRmdmx3pYuKMDN+L+ZLUOwDgEz6DhckM22h6
TneS/DPW1ORDVrIjPI5rlpjMZdvKxre5Gv2hWiN4owZm+KmTysHzAz3Ps6wIGukWgNQZoKDGIGU5
0WKzFmyeJ31vdh/Wit4bYnfwgMgvEK+ahfui858BqzbTponSBONbxkCsUYqPWbCQOjXjmLJO6umz
0u/7/pklFye2wlN6I6HGRFqYY1dzgn7msY8w+akNsw/2rYgVZltovjC9PAKX6d1HFw1c2B1Ce7U2
8S5Bo2bZfUqqL6WxkUa8tVbBw1DWXbN2Wh3aIjo05LVwmsJqihN3GakxI3kCOLr6LbOrp5FYcs5y
Dh8VRkFN09TjeyDAe8pJKN2FmBxDGIXauOPISNC62LbUYptFJl9rZbCsyjiuiLRTcDhQi7CTOK5o
getBxokMumI6HXwFyaDzV1jy6WttUByXSOaX7uhOIyUcYxewoUW3xa2t0pNGXDSd1f+jRQyAbFnf
rS1eE4C24RJrSX+NdHYtPnqtXdeuMp8WXGvQhI9q//T/ydBx3O2rtz7/NJa256JkgrS+dQ874EeU
arbhCvxyoMjEMINqdu81TDNEnJzjXUC+UMWwGYzUythat26R29XdaqaLWV6NFIbkJrXBXqdh68bU
b3dL2/U0RlqbIp/zEEKI0qfECyIM8Ft7CeJCpwdvu2z1pcpf8bvCHsinJk0tC9QeANCpeHAvkwUU
Yq+X9M+Et0Eokdh+kdBL3Psr1jeXYez7+BD5HyjHi1MApZ50+ps6GCO3LcIvW8orR8XIa/qAQTAz
Ps605pEJc4g1aIQXb/zUNPxnhEtmNd9rcNeW7bzehFeYjnLQ2gObMuFYlgB5kTbaHqG3uSDje5Xy
psKWLXSvStxByG2Qf9KKnl2BOhxhH1b3o9Sxy14NysZ1kTdOliq3yhqUAbcijw09o15vcefCyii4
TbMeX0/yfeyQ4O/pcRqg/+a4VmZW5YAAWYl+kfzs07ODC5/L+aPwju5cBQpoGic1Ki9WcIFHyV2F
RJB99RpoJj3ciQUDxDETlzIATKK7r2r3rR9/hfduY4T+RdsDi7Bqau1rme0vwKKfFHtmfje620UT
NH3TZDmEgmwHU3yap1fb4ZhtYrfGwjh5noK2eb0e6xItRgMw5xepLi+sFBoeq0LZEl5sq4IBJiJu
ZJiig4vT/THBsTpSEJMFI2h6inCAqNevk/CLUq+bF0yjUmbjRKsvvL4YJG7I3OsR8Zrse02Z/y8m
sArOHHwinzJU9HDVJNviofS1Y9LX4tusfcdQ63xzhjxShuQUgJia6CKzNN0WI6nrsTYUmmZSt8NT
cmqY6uBSZN1BnepXPF0wSp0kLXQ1hoF9riu4u9wNrR0iA3AhbDHV1BrUgJazrk0kUlZZSCGNx9l1
/BlzYk7H6j1IEhT5WxvB0sTo/X8J98fIjOgF2YpfgST/AaGTTKWdIo2qrosH63Abejt7HDfrZJGn
Vwj8W6GyzqVvEJnpu4n7VpvGiIDx9GGQ63wFBNzqylmAMxFACveIL64YrVzISlVzh6ye7UPDURsx
38DyblNySoI2uv7BtxORY0C2eOl8edJ/x83qCBZnqEz1II+QRW4R1gGjbLtx6ythhC6xSEQWDwvg
YpzhcZ5bysdCN+QAnVnnj9Wf79OUPuamHj+Lzi8UxREAyjfETD6hg7LvzHi8DmH1NAYMysJOVy4G
6Z9TlBc+FjbVTA0HiBI/EXATzRqbROzvMxc7P0oGEZPhq9qHISbvvFxqLXsUCMQ5Z4ZMdX0ehTO2
DRjiVu9B5tYZvnlkQ+X2Y4bhyCQUC8oNrSgU+WI3iqid4c9qlLznW1hQKN626VxQRan+c/UuFz2Z
IOBZSNZvX6rOCpGuUQRbIlTJb2ZSm3WlPYwmPevx0qqo7fMWpFgLxbeMUM/RqVExGWXhvQVOR9eC
v9hrH5v0awG/r2H+SgjbnO3CQIiuSm9orpaOvk7JcX59ewBL5ZHvvcUokcLnoKM784HLrW6dFZvu
9ZRhjjT1595Yp7DKJhgRQFAsUbw+Ru7gl9WJ6gjDv3DHOM5K4p5mbHR/gzK87F6xvBv+nAMJ1U4p
eRnjBqCF+pdDz3wS2U2Tb/g/o+ljyYgibf39Dkf+eCMaesiBSkk2T9cGBBezcJlWrXtqpvf04OYL
PQPUt3haQ1Bog53D/yyV3awpeo/Gq1Yy0A4vi1eqMF7XShdtrEnnRacZ0r6E/JJNk8exE/GaTrCT
aaTpqgfu2Dtj1Z0bGnUhOvQa6vmvHtrMAfr1AhNSqDQtCeNdwwExP2f+mlX8vB2ZnL3fVDwwrEgm
HUdVTM5hpxuDP/9oQOHsCL1wF1ajrMgrSfA44rgosftJXMbFfPdqzOM5w6gflHerdq2vkRcaJOIA
FW0vZ42BjdMpXixJgtSOS9UCgz0tXrATDrXhsX5O5kAncsDun5hi40QVbay0D7aT8ufSoimwF6NH
2t29zqlZBrterAI8zScKrg4Zk0y1XYIOuAdKbuxcC6w3T0g5hWiBDtmbE/aVxiOjiquFgSI+tGJm
AVL+zr3xWS+j/DqhetnvPW5q870ptZObDLpCPNNga4/RGScpQx3MP+fMvSIBzQYku3gTYiGn8F05
6DnW6yE74Fo3OBpS1d75u8eI31EMOhNaEvDBYlWKYvYBtS5C7MCRYAuxs2HFdm3GzpwNbfm2AeGE
RsPsCVAKks0oudAv5rEZfFB4S1CZ8BRXUtnpp7bWzIHH7ZJRTZdmJ9EgjFPNXxplbjnJdYYBmRRw
nX8y8311nIiAHK7Cx9R37UPi//HwE9ZrQ9P7NPjVQ/LnTHgyI5rD+VIKJjS3uFcr8Y3fdaPUUFoM
XHTB4L340gwoYhtTw82rtV4vKqrcFxz3j4IWsZgm84GoQRSRQ4q1RavpdMKvTxO/MaeqyFGWWij2
d+4mXnuOe31bgkFUz5cEDjCqpefwAZbl6KJJDcxxrCbF7M9KohxlrETS7H7dAxymgGgw/PYCPA3w
7uusCZ+V08mpjsvGHtNModXVK5TA2cALqNK9asUyvcdqpu7+rGEwq3cAT5GSlTey4gjoEIsoDzRG
r3tENrN+NjCD2DQg9yCSV736yb1N568cF6F6anaohaFGSgGcnpxWFfk2NWyQNH6c6I92Wq9HUkMA
gC9u+WAnFWuITXI6bIQM2dK7hWHwuu1WUAUrI2hqFONLH004OxlbeY9aymB35Zlj56l4xFlDqcgH
zINfU6OF168d5p9J1K51YfUVYVngVE+vtjpmCLcRPmBICmLbmhiHU/30PU1CfBGkufzhsMjkHdai
/TIR+ToI0WV/vLs71c1vjgQhIMX0W23Yz4afdO3tVrGQ+Q2GBPF6s2dnoQdWgzwOOIqVF/p81CZm
q1CWao48/0IaJGwerS6SPgQZu8N1v/o/UfiUg8T99AwIsHIDWrH2fSwtCXmXmhi/PoNUdqT5GKDB
/e0R5k4bXYVszBQQ3M3Fh6GSnfIKDaUKGwCGgMJbPsctXyZPYB4N3fuXB86VNp0r92b+x05u5uym
1rvktD/S3HUu82IMRpP5L3kiI7XtGQuix3IuBRQ8SXSKsX2icOETLUdE3bYLK61zM5Ss78OUYFc+
PXJNb32yDnAP99lPyUG1adH73OB7nd3XRPTxXvWWFusbpFmqzNHkxd7TGcoTldkfZQHki02P6gS5
DLej9sCMQh1rBYVVRUM07DoS6eJrKTbes12moA760eNEr1lOUXhAfNAjfLgBDnFaXo0X01BMATq1
hlrBzvX4q/dmrpv4AmGmaQmpS4rQKTVKLDH7lXTYR9vpyX0VFXRsf5+wy1apBNjchXiF8YESmJfL
kopGf9SW10opltcIXOlZQY1KDhvVYAZOYc0v8LQd68EmpPOzvJa+f73g4BP3LVuU6YoGUSJWNugQ
cb652UzI0XKfc3nr1OcnCJD3IzLmpzvV458SfvcHOlW6BJvx++liD1z1LR6LFxe/DUPTkTSftm4v
Qg3Fs1yZ5zGEC6gFUP80LcsPtJBqqJFeAMT7QJ3hiQWHTpd8V/Gi2qB5UoSVsTfkBdofkKVEHwHW
BY4E7IZkPJmm4+bpQ10CUFLbbJAhmJzFatuP8ZX1ypkf8AMIX2gXnkMo4YaCuCgx5vvTMaBfCJ8I
LXEKZks9YDBYXEBrKNHAHevgrMX+d2it+NcF5xPjLukK+WHJhnJlUKwrMALhkXNPyZ0Cimwj1m2c
kpqr5xp2F+4T9/FFRvszJPsH+m/Orbku/2P3Rm3BbbTcmc0hf3Fa/othP9Y6if27E3XU1cUMUHqT
QmoXs6P/4a/5ox4nmc3h4bPaWfCXj1flE7sSg4vo8601c69DaSIGmV1c18OdQygqVgRdjJYxakHb
CVBrbqUpkYjRInsbBBoCGDrL/DfMg4oKddi8y9VbZrcUPAkwIbmUgrCbylMkvsVs6znb42sKBPWs
+YP/HLC0GbSftgglF5/K5gfysSIlaiHo2yyKGAD1iRKvBgEz7JPri7gjONA40W2ULHQUubFTb5XH
N3doQ9SUedzywQR49t9B2yW9g7YoREJXxL/0Ds58ojTWbnX6nvpoQd64UD7J3bl6/7mS5hyCjCe5
etxYWQePdHjn/KDtj9fyRew9YdjrtSomSC+6PFnOPTHpNaOLUFVqr6ugTFZMAOlARudzhvEUY4Jy
d/OO330SrOEtzfihcdkc3ivkkz5JWUoxUzAdSTst8hF12Rq0E8lhW8y7aeUXW8mkfQLsPkUmPTh8
xokctMVVYneidKufIMWftFF9u2WwohewYEZhhwLWOHxW3v5/IJU1A5ylGo/GqR5oeVXDMIJuLuJc
ayeJCxrv8kwkHJBDh+ORPGd0C3DOsaOmiq2qxBlng2UZXl6smKRTTcbacixVMqHic0vH86uXz/Bj
+AMFijav+s0BW5qrQyDbEGvBEdQ27hKb3dI3Y0YZ7oRqkcuaANmAVYvGEMScJoyfvE89KqaW7FvA
zAUarfFVSVBgf8mnGWR754t3k5uwm/IeeTrjEMf0Gpc5CXU7sdcF61SSX9bwJeBcPPoXHscJHLcl
+OgB6CcPCma9Z4fQtWksMKLZZ4wLbhE4Kd8vBbXf01MrMEq14OoK/54x3fLvj03BfkNe8ZbnjqkE
ASoGIjFHHlhuLhjv2TdZFnz9/IwHgiO6mI7LMFsN1bQ2OreWaSaW45iye+dwfUMLYWLkAc6dI0hg
snoCYYZ1d3X91tSHjRyVtbyi545onwPHSiF5IzPTANhHbpszIJO5A1XxP/05aZyTbYB5dE8f5iIt
pu936pjLoKiFW7ZAvTz6aLdFvGQdI2Ij9S6rVIhSQCTsgVSGEEVw22xluCeTnCdgM2Oxjq38OSGr
U00Rn1nlvOvdxA6F9sFZHQ9ikgGoXLGTPq12KIQcl47U7v/1IZshr83hU5LC4yqmgXV3tCOU6yQV
SdjwkLitwC2KWLxNx2vCf496Jzh9Zt2yTh1sO7290PPme7L6zI/3q8WB2WN4xsOOEKYXweX5VlEO
dsquJp4F4CgAUne8k8/UACof6IssUjEPk7ISnD+CLVbQnWHdN1QBkcUBRLjn8JT0efnYyvyZte45
clAXL9czc2TBsBAkOiYOG5VJFOBoPWJqqGzyuXE5tzPvaQubxYVKPV6FOkI64koyMBLSItO6g/h6
hoLuHXcwB+oC/YS5gFOP3RquisK/HIeHnT5m618eFlXEJkKF5D60pIWvH/10L4s1jBj9C9zUpVZl
e+ndTsyPdXqnK0qSQNn0v/efntQoAhTpVwUh1WPr/E2WfBHIedYfHJC6xnyy8genQ9tqboorslyI
oSnhGLeBG1aIe07tyNDdtPGK4OVr9iBOD2DI+wSD3I61OpaadbedxrmA6KS44NrKKElL0XrAfK8n
KDlURoQWwcKhqb8CdR0vs/hl2NGt83B1qhGHT3XKBobcD4TCZN+Vez+kmBHi6lFy4HCCwdBciujw
vusyy/wpfwpOANek6w91sWByk7PItCstdPFoP2F+6TBjk95rwMRukVVsZGxFM4yieUx5GD8dPGlZ
v5ihQ+DSpdNE3n17YaO4M3A43ppc7+V/Rvfdu3t+Hhtj+FWUeNkgjKYf1mSmIqqNqxHkDUIQR2K2
+0OJ2r4Q787xVXu98wC4GvrepJLoOR0YGoF2YARt/BakEdBG0hvGUXHrjBsJPXVouXVEJ0X5gtfo
6raciGeNcPvfYgV9X4ITADxmtpDrEGqC8Ca8OlykLsbwKm2dqxp/h9DHaaVlD9aAO0J+qBPqbqR0
4s0ZWjiOh2MaDKakiDailzMkeatPUkM5ASncGt+PerplyaCaZIjDcOmDqWSfLRWVHNmFmgfdLtq8
Iejb7/O9r2V/hDhQ/hr+AG0eV25be9bviuzZE8TjO5niwjW0Y8PfrSQqJlFg8iQw5Xu8CZgJjM3q
IwDa8YMBWRK1JmNkC57dbn1h1rvbsFNsgFkr2veyxMKe5wT6Viirtc5jdZ5yp+xiSWmgbVltTof7
N3knzlGH4HBVTAb+cdW6pifcbITh83oF+ww12CDRmncsJzU4JPnfYa4pls1NLfYXrXtqIkehC28D
ob+IWzUHaoutNJI+WSbuU8vPPe15KIo3jKcwz/VZj71qJhDk3WVu5q5zg/JhRZDjlEUGVRkAjIxZ
X9WWvB1KzQlNvvvtgpTGmx25kAykpqcfiY87guxFPuNcgSSWU3OR0FQXCcLQ/kDC5E961fgqg2xU
NnUxk2XSicsEJs6zMn2RIqr1NKXbHauCkl8sPS1Ktk4C1nKP6uFS/hVz6a4lMzRuc0OgT4x9Hmi7
IBdToP7/ukkiBqu5dSDZfpFpocrjj9Q6eGOad9N1RkytaS5EYENZTA2Uh83PJs8P2eZO8cotjiah
yOHPEEvSwwsqmVMDFHGlbWfhSt1BV34W8Q54oJpCESIYli9FJ0eMRAK7Lk0iF4/FvI4rirrax/pd
XSh6JHS8+zDvFn3O+3U27IZoj/L496MyYJ9LJGB6sgVqLLAJH1PaA1VHSk4+GnVdGmilKHNfzbLc
z0uCdnUHVmGbf6+bKiBWxt2XpR1x2YJgCg9h5jxeSFKupWst7qOUAARYg8TyNIgYIw0uDWywgAd5
vel7l7Q8fSdCu3+OwU2WqIqcf+knzBFpL+S/LihSLsBCf9aUn0RGqqecurLFgz2sZMr8zCgO+Wqk
cdrEISuDmVRh3rdq2E+3JoOSTrwy1o/04aBfnW5qV4mGDNgDk6VZDoyJyILpDseSNOnIGlfV8YJg
+8Ioch+3MTXouJZ4I5vXFfc5kZ87ioV2MYWO6w6OVSGY3hni3dwTz4g+rRNBbEdJN/7gPuAnagzC
jFykz+LujyzdhjH3p0YZ5whLMpcfB8Je55Oc3FgOvZzzHNra+XIaeSdL5PwzC+kYCdPzzgE5wcDS
f9vGZrdprs22OIoc/MEk98YLGsXMs1txTZT9bb6macU8VaYeyuCIRFJe3UG31NPN7M5WaoVW0CD0
fG38EdOdeWrlarQmdu2jW49knARVvR64jmK7cVR6CCRym2Ucr27tFTapi0DuE4YiLVtfyTiHZzKe
Dvgm0XsOTZ0yeys6GYkxNUby4DB7hlZIWlCoW0VkhfK2iMytBFiSlkcv4guHNGl2oCkmGHrlpSM+
VtVFO65GsYNJHtZdwZp+kG0Rk5SK+UgrhfbhY0Pdn844I0RV8A206gOyvrk7amJlAkcMYL/0x5Hy
E3+XJ5WwWXV9XWkXecdZ/TrPyMybBWv7QnrWq9VDm7GVUzHkYiKwToWgS3RJ5y5QCmIB8PoUP3Nq
g8TZ9uz/9XSqdMaJCNjKtKur05eNcoPZqBN+ek+ewsKbXXLRVDDPTmS3O/G4pTeCM+eYHYUd2G9Q
qiwBAucEZ+AoXcA4j42yl8Rjcw/ragnpCC4pXh/Gud+z7u6x582cXXuoWRrLI5cLTPYhdJRla+gb
BThkKDnrWWw0ZsFtYCjsSku+oBojgPUpUMVwgfW3I+PEAWdHMgFju3HwYqJYP7HRtk3OKpAAKnAn
i2R7Y1TQcjpPe3Oiw667zPQhykI0mbL/naTUeXFcc7s01PxAk6d1izj6T1UBbmvJ1+BAAZpPbOtV
of285tzbDuH72VsNZR3RWdGq0TmvLPAw0rYl+fxSl50mMupBU4WVxTitf22vx2/3PfTHwf/hzLm0
KF7e9shwdOqwRrwTQ1bFaA4LMOIMVjR73S15qcOHPHiM3BURUKu/qgRMCPFmbVnlaXNWmJ1tJd1I
pgVP8E4qdzKiYILVw850WZ59zVEWIGfEPBPMXtmgehMQrXvwmjROnDNITZsY7QAFNYhl0QBYdn02
wZbCpdqhp0CT8HP8DvygsSfEHyPLsq9Bay4aVCfP1Utmt1B4tOH4DJzsqShRfvomHVcizwhLsaQc
669JyUpSED5viGxDJTzCai4BGddmQnQmRy+lbw6FcADRvIQQiAeqh8chfok7sODkyKrlp3Pf0ZbX
TjPFt71wj9ILg4fxvv0bZF4VvuHGWLSWwtB8mbwYsRYS7lW1FAQGNDXAPxPvU3MFboEiahoaSvgq
aGBgA4buJeNVgfenep0ci0jO1TuDSi4sPf29lZzwtxJa3R0bo+Kr4HEBvHf7G/zR0so7z4t4mj5x
07/6bOStLch26DLZ0GMlGOX7/9uqLDDKXzDMj+OgTMWAPGELcKeXCUPip2joTUy2Ixzzl0mr8fgE
5fx8zEkRE4UXO5Pk4FZJNMDXdknEu7PgA8AcIg2rjiwMwGS19X4sGvLzdYz1j62up0NTAqME1/lC
uNaCu4A2z/xAYdCYvh37BQHZcgOi2/iLroj9XzXuGgLKIstziKcz4w7RVeiW144ryB0iIlcG5DLB
K/xpCdommnRIxtQ9+57CdiWSxSRMHCLtEKLzPvETKilf8mcZcd8iI9wc1I+HOT+dJuTVVJTiI4x5
VXyUkho02KF2bAdb3S+zIW+6TFk1E4n4tbgQfLOw2ukl0J/5uCIxP0QHFDRLnbI7BWLcGtiC54t1
x0uhgJl0UAcb3ij9L0nA+khHIGCJqFYP2DI5RvIG8xCIIXiFYKgHMDBIX5txQbVnh+kjZxSOTy2m
cRiakoZNQ5BkpABVq2T99sYWNJLPUfxDCCHNhV5e1Um5ppOw8OnICETQAG58D7tMrUCOLxArWeNX
tOirhojvyazyOPUrHcv4oZFt/nudkcu6lwtfIiBaVuTDvFu3QywB3tzpQ9EDtkj+0y3huBaeqcFa
vYfUKzmfEJslg7g+us/2yIXAP9mzQdHoSlF6qX3EgxrK21+OE8nnAKuCDPJ+YYN6ecmcF5PjxgQ5
8zrr9OmTUbJ6OefuZH6ILudc5nVt6yWjxA3pPL7AZ9JGqeYTI1vj8P3CFy5qvBZw/S9hQHXjaCWK
Zaib/0w2U8LMUBob0rU0QmAm/nGQREYkazhvTg+IFFI4kTufTj7nq1cpac/YZO433Q85qTA5A6Nf
GDnqAz+osUd9LBniqvIBAuDOtUbiWq/csuzl0civH6/VMpuOYGlph2lmZ2YnPCPE2J9yW33IkcRH
l2MbHWRr/cqJzmg5I2oyN8HDzzVzWwLnwv+znp//BjyAHnIPk0QO39k+OTyDB9Zjh+KboHgY+T9z
r5RPFoYzL4c5L51ozLEJ/pTyNvhFPZyLgphMyRRiGQU2xsyAaiptw2E5+vA7nlEmaWoWePuZkVp1
LtTet/Cr0waHdkS6uVycVa7ofatSJPBsZOgITMFTEyRcpo5vCqBATrY72YvIPrL0KUe8ipsWILff
ndayxc5BJEhDrpvSFDUVlKrM4UbVvcN55bqw1fpAEtZChafVZyqu1g/7Ds0LKz7ElayEeIff3waN
oEjubrvs49SKx+OlTrxkw0S+IE9hf8xtW6ny8eoyk1LunD2Y4EnAoVeRYxu9RzhfM+UPZl4rrHCU
aPi/BT3UXg5C5NCP7SX9N9s8f813tt4d0dVM7zfDqKutxizRrL39eFkLQAKUVa5B6f4axIuOC8MO
mYFd+swnFte10aEZx/UAQzjALSZ9YXCVOmBNA+c9oYvEpZ9PnHFqRMgq0M/FEegv82TdJuqxcuie
rF7EAXn687dknEfxAYzyI+YEaZNZrdYEY+IsEh6y78XZ8Q57mgP4BOE4topS9pO6UHaJEYUi96Hi
HpH2JmBiMZ7R3e5WHLEZdtJenc1t4CaCCW1rEiNiRHpUlfgN3NWqf4XNWLdvvVcs/dDj1OINPmZ3
NgiHRI0FwawGshBCJj4xOALY+hzXErlCENnbEkqFxDAJ4Y9mLIcQdiyDN5+3SSlTwBkWgvaeIYQZ
IN3wxGf+n3TOxWfj0ooVdreVkhhvP2J1rYftCXVM65/MkOiz9a3Cz0VbK1p0ufg24QCvhUaOSRBD
519TRwEPhXPJH2eyBM7K9JPEOFmMF0Ik6UscM5hKnjFzQtROlRmTffHkAr2NvwDbHizNQ0dfYVTR
r5l6AASAk9coXdq7BzjKTjE0aBpGBjK0Prn/2Xlz2W0Hl7QUDjUSntLrjIBgUBAak1xeDaaNpHRr
SECF9FBA55q/AsTS2zIL1vx86EHORICFNh1H+mzkAnUrBBYC093iEWe7N1ic4diV3hmx++0XG/9n
9kRTP3Ch5lOX5Wm4TaZ7apDLAiIWJWNdHfAUpptQ2sHnezMjk39+T/gJiD/1sXZtwqF0wbk7mAbw
zp+2cg3TzeYNn9iGcbd7JkX60geOlU2UussOPojI130VgAq5N+H6LdCx0XhFoDXCii4eXUaLuV+C
1KcCHmRIvRX2bY+zYme1bkbftCgz7vBe6lOZG4GS7PVaP2pENEzC7tMcUmYk4QqwNyfHedV3H5sr
oXjwth8+gbPrVNG1OyWV9GJf2tdRD7MU94CRPABlPv+nWig7sW4a9tcA2R4iUrY8XlX6G8DGPix2
kjMrmZvDtVvPzKGEzepIbXGjx1hvxV1vN5PBQYK7T4FWUombshrRgG84GPt+zTTDiYUxjx5uXPU9
LFygxEsdo1NfULJzLKTmXIc9j62IWHsKQyEr2bfmDytSMqPvj/WrtvL05zLd/zydqIzDgK5rqb87
0xZbK7Htwv2Caqkw3c7uFl6h1On3JFvMyNbN+1HlSTDCBwBs7IBBy1p6r6nW+IEdrsnC1rqVDDxL
FxUBvAhCmA6oX0gaAgEA+jUi9qbHlFsP1fnot3yyu/BqBHMK2qjLMkFEjvbkJUGnOPf0M735GHsh
eCHpGQjyGOVd04e7HzbvPN/TFmO8b8mo748/orOMhQcYd0SsPWkE4jeANN+1X4mdKOubfpJY77np
7iuNKzS7u8sJOWYPBjxHSZvmxvBQvkxv3YOFmW25p0KVR7UtaJrWpylmZ3w6v5SZZ0CU+29Ls5RX
TtoPhkFF3hYIqNTnKhymM4Ia/AP0/ggl+kZDMpbXGwGWUD9f+4TkvRFyONnpOrKNl5LlQhocpz+R
wOlQs6dSHjXmckEBgRZJAq8k0GI1g7nPhqX1UcrT6RBZi55+5w3Koa7IjCOLiSDe8MFDa3nVPfJl
boLvc60/4MZTNMcPSpK3Iqabb6CE+lsDKeVi2U4wTFLq71qauF/+eJte2R3UbRGp482SaUCbmwto
S07bSYjqlQrAKcIm0IQAjuCQ5xru6vj5jfXHMrGIgzhQy1MZ2OrY2zGI50uF5ElTkjlD1BQTzHBE
iW5IRULnjpKC/lxOOSVchPsdD1YQsD4MfFFs6LQcEriMsVVO6Xf2bdCOzDqyZVDf8LjhKfG9Piu0
ro/1Mo/nWxRfAB5aTezj03nkN8ve9a4WiReGSQng76XlGJddyak3wRakrqnVx/UO22eSP+X9xpXn
2b7tmtLN5TF4WIVBYR21qDg7vAhBP3seUsmNOfdJJQf6lWwoP1TOmyFUUoQAuNtGJ/OI2yGOLV0O
p7P0Uq9pLXyHAT4/v6c5w2Fy+vR+C7q4A722SpNGEsFGz0Qx0Q6f3huEuNOJL4UPEAPuNSqC392V
rMPtKm/UsyBIQdapkiITIQ5IS4U1cF0xbuOi5bSAm+WqFCAVqUDY9/NixTVURd15lRtlUbnHUEIp
Ygm3HaGbbCcDTlf2vluCtSKQTIL+K83RHuITA0cKc404AOj7dQVF2Y5Xe5lHqdrhZLcwnlnFPQbx
azQR1Ks51aXqzoMU/bTm0QrD62Yp7vNJxfT6F2Ixr8YSnyKae/kQ3dQNTAphwRzsFC7CIKpVGG1F
+ODurDXDH9avS4+di1P0J7ar8QlCaJ/lBMh4vCQlITE9rdv7SY9+iKCw30wddSF0QkVjlM+fZ8zx
hBSxd29rICrt+xdaK0OEzeGchsfFWeehz8dwuK/X6eR84hj50seVhndNx//tmGgX++Vu6ronQkkP
lCqPi8ZXv924Y8NBtd4CKA0ZraE0bhTPum6YlH8GDxx9XW00bNfHBkkfBLQBhFfYzbSBl6LSp71Q
+vMrydSWaE+Un2tePGmzbpd+TKeDsGqSRqH+o8aOX9SGMgLLWR0BBhD+RKuyDZb8ljvxTumvrM0+
f66jz7kozYwoPqtsTfYpmU5+kOVFCAWQQaO/aU4RleBdtK1U8serTxLRGCbmGx2gR1VUX1UuapKy
x0+3xVUsMVHI06Uo0buvh4CyUW70OZDhnmQjat9bha3A3TIQfGiX5CabK75nHMyc3DnUnWocrpDQ
kRoh2NCWtPTxjlcFEuZOfB7RNUemi718iUmsDLYDGkdlUBDVjnfCc++c+NmhKqiM8kIrefn0BoJ5
XFaYzkazklTCDNFZm0beGpCWfRduQYhTlmPgz4h1uiCujwV3BcQ9pcg7YCHDEQmk4UkCkuidAF67
eZolEGwd/1zK7kvNgOXSWcEMHURdCFO/t76DGYRfJqF1WGN4dU+NlGLhE9URnWHm6RFGYyQ1yGks
x3puQiLf0Xyjf4ErWg4/zGFaV/C9Va2vmmUIvQFM+yPZ2xVcD7OKAZTNClMHBvVJJ5XzR9cnnlqm
zdXJaMgRbS10o3zHjISzMb1OhfGC5OyIVOSk03gylkRZLjZ4FXwmB1LQS5wIojP8bgP7pTPJq7PC
NMx0Mmir2UqiKHGCCNGBR4h8c2uTlk//FrkYEWkSCv1Fp7oZmDTEzjn8orN2K0G3GNf5SoLRgi/9
mcQiLHV7AZq09Z5Pz9LZniV0HtB+5b3Qu2HG1+H0kyP7w4RGGNTbVMsMtd+2Own1XP0oxzeOM3m0
Y7vknnZZj/z1sN9sQH2AeNElaX4LfelAS4q/rUm+sWTydpx18ZaAdFbirzotXD07+D2CMLKMZCzW
vU/2gHOIB7elC97LiEyxxRe1L40XNGhbyZeoyKx+eG3rlMej4Qql0wKpky353709MergYY+gzetK
B6On4t8+jzyKQUlOUIAj8Q/F6rL9MRe8zTNDKdumIfXQHT2uEkIfStjA1WTs9+excsVbSH76yCFm
U7Uke+1fQpdyY6OzAYYy2tU1UzhC+S1dX47W7T+UJez61uZ+Sk4JKrVvk+AKBpmwnIewi1+Vnp8j
Op+I0p4gOo8nvV1ekOxkti4cTPPUNnOgmYywi4RIuPJ0bJZsYBV+0F4OlrhRph0wdBAzNuk1+59A
81ZkdW+oMBubSaHhneJ9kB6XNvqW4EMhGTGkhMa/olMqNQg74HnqFpnKAxTyMsKFJbt2rkZ2I4As
xQfC7tTW9unfoM44COhI9UlewEtrgSLhox6utvphZSo7HU2ELqUAIT4vrq1Cb6TVodwHiAvG6SHv
8VrK18WgegL8T9OwDt5TR4lcbfZsalZbL1YpiUoL6IpN4WvgL5jGhg1pNRzYDb7kQoASNJQnuKbl
SRpe9j7CgixyaDVUMnJWymwdvfBeJSXHedYcH2gUjWos/M53+TyeZabwrFIELlhShVs7rTKQn3Ul
CrRcCkwSSaktOb/eizk95xvK67tdAopAb77iAkr6wIA8IOmHwt+ujEYtMMmFmu9SnvZz/NXpc89F
7Zh4MZCHExLdxqYKwtHXNtApIevTiBCKFGKZ7lCq8gKVL6RlPeAwWAkc1wuRK8RwzIsNs/GboG6g
+rJYVFLn/+zRHgoDjV5f42pSg0iAodIru2lxuDr3AvWaeJnpCuk6wxQtJooyQ1W4NJEDIPkKdLjK
BIx0rTfE6IoizDR0WzrSjX60CnAApnB97jLgb9/lbHgsz1Ft30ZG48fVmxCDrDtuTAwPk3dl9Jy2
TBtQkkdmvAThcmdSCqmAZAIifQMO3i8bxHqSqLArjN68+guoM6DSUNAzpe1eRwaKzVCZEr2hOaXX
xH3JSAQASTaSC2CKZHqqPJIXlqUMT9W7M9x2OeZSJBIswVUuDyjEe4aG97N9Oxg1xQ2+hH0Dl1pv
Vq3ilkAljqejHD78vR/5tcqt/CiOMiY4X0v1IpjEmOZWV9KmIe5nKz5VJPzI0eoSCcvUKAKXLYVY
yoKF9g8DEmJhpi3Orik5wZLFf1GKYBNIDcPLqJaS1iCMOJVZZj4+tqu8IkExo6ic6G0MOPb4N2Rc
uXuw3H+r3nnk7KXybNXpS8W08dtMiLz1DfC1B2k0dXUaGO8Ipo63hTWn9Bo4uSBkcBgjZmfFtKvt
BuaNQOfdSvEt2Uo/TRlcHM+5zJfsZQ0LcVLaaqoEl+y1xjZJHsFHezxKDfBkVA+XRt+yo3QkG0I7
dRL2B3kPwpqumRwUHH2jI+ZmkWqxViUdLHzUGH3p8WKvDmfm6xZIeQa1utYFUa/WFVcOKbGIfwdZ
x69+3OQwjD/fg7HiVfoVC71UjUX/cmGtxBboNi7OuCZJ2AE7nM22tNyhZf/dCc75tmsBVqjlgqrv
BTMgZjDJLH9ipGrCkcVqh5x8GXOM/gHxjwVcOhAlq+QsPI5ARG5vx2vNDxGOgTViSaZTKckFgtCy
bIOHvwjssS+fpsgu4g3HXr8tMbsAWvmkPeg4owelgztqkYEL6RZtmF+GdYX0cLUZhdWO0cTwN5mF
BSnbai76VH7fgsgCQIGgPQieRTSg2a+CjEbmDgAqD8ytfXt/Kv3w+EXFvohXQRmY6DH7QVuEjkEE
eMyVXqXZJFKAsiOWrsKc/mP3KHxg5V3SSZgSia35X8sgfz90W1i5U+lwhlQFyqCQKJ3wUP38NdOs
e/P54TVMNUD6/Qebgtigxlb14MIevzxjFPyW6FxXmckBl7kLwPgSHzLkJMMM7bWq6vSmM7Q0SbBE
/p76ws5WPfAuLj+G5VHKJD1LF2StOH7RJI0M1Rnc/s40gp2XWM9N4uxPC8zmK9hvMTsLrh1eLM/I
y7v0sIBjjRjiMGt+0o2t2tLoiLx1KDtzr8WYQL3NcA7ZWAKCCC3E703Vl6QlmQNKdcZaJKW4iQO9
39c7NAM41mL/7md0Jdx2rC93EfpreSAk/e7HU5oOxc2V3LPdU9LIgtRfYVXC2QXPgBDV9klWZurQ
Wx4ZHWAg0u+aV433Ify6jO0Vz9UHgxsnjimveJTN9KvfMWOZ8oeSOl5xoP1zanvhG3O7QSANgMmE
JrR+TdItVbkkOwPXi6+mfzZ6PRx+LCUD1sjSf7mWxEKY3N9N6g+di97VMbITOMDzjTVAEjC0wXBI
CtV+3hhArUiPCaEq9hXSqa//vdKj3AzDQ5sxtS9SWKzgYrZ0AlUDjm20rCcOM10CU2Pzb9YlWrz9
P8q63v3oK/CooLr/hf8EOcXhVWW2DYGbjsa4QMbrq7ChaWn8gPTr/MRkPAnrgO6VFNtVdGnxi8UG
fXPIfZxceT0WpBPPJyAEQ8+fmp7iyIyy9SD0oIP/paZVIjl0SQIoIx8bJAc7LHDFFAW+L5+9sZSk
Nx7AVwJ58Z9KY5uey+VDXQHpqPPzvdl9vuoqkPbGHxyaBIMNm/6YBUdcXofokVQzkzcmUS4ggf3/
K2XgbMCXGQSx1doVZKERoLFNYLUh6yy4yylg712KLx7dKqZ6RfYLu31jONfrFAmFPeN//w+F8TpI
Z22rxkbd8mCpPLOU1IZbOTJt29WL+w5Br06VzuED9gXAvFtEQvZlc5TeWHVwq2A1fIk0GMECoCUo
H7mkfDSyAq/TrudRddMH73AuxzJ/deX3AXa9UpAb2RsnfNQN8S9nW9rSKKjkc7ONmViMlWhaIOE7
lwWxoRN2SqYkSo+J9Q3NWgQjy6uNgxYpnoxT38RcrW2V9zqVvM3dRAn6/aTgQ4TmnJZeWQbBRYDg
Y/XW1/U3CsFibugzKJi5Fjqcbljn07iwVD4mo/LXrTw75Kcx0CWgf4USAxRKqPbTCBG880x9S2+9
3nDkkEIpQTWIrH0bHgDjnxI7PdGiGCZnY2m9B1C6d2MHfzf47iamkHs8Ytr55euMvy3loSHsh+x4
PJu4VN7jNW/ti2ItFmw+XmDsFvGV0QCeCBFfAwVszYrS2Zb9XvKP0FDgtwj8ufjPPDR6DZHAKDxn
LQUZQRWk+jXXnVuTQT6UkXlGhbQXvmoNYqTjqVdZoksJo+xrN98BrWQbQCUUVfpWwVrp6ICirghz
O4qRHxJz3vQxTLpk3aTF6ltelipjKHkidD7R62l6O0mEDbMV2MU1gVCh6yLm58ixqHCOHt0U36Ok
eR/KzageuK/3RUdEE0uytNcT8BPsi5krw3xHvimOhevSrxY6OtTVILYBeAwhMK0uvlXkzefq3hc3
LxZUiy8mzULjFANzPHxz6GPI//zcK7D5KuTq+dhQp6GF7WuoSNK8CtJd9Mfmos1tPRGpXXfzdn0X
aG/+PohzfVCNWuyy94Su8Pfuzn66PiKdFspeDC5usn5+hrdGszkcN4e056W+Jk2PDsd7Pk7kFc3n
3bltnkmCtY4ryEHZJ05rp2XvaSfzsFpu+lDSjaKzPuZjjK2uhF1UgnZGGD1ubdu7XUzOYILDaZOM
ORg2Y6FmJ05SnZMeDJulAwtfwgZHBvvjCDuUk5eNqIxMF1PJGLo0QA8GfZVwA97ksQpEyfm5Pgoq
lqlvGeNinoHWrdp2r8OBHv+zOehP/PDfmzapAEPJRLn5YB3ha7+PE32YYgziawQJPbfXS2WwCP1+
+6oD4nCpriQOVMGcJaAQIEAsqOXACpZjLwIU4Gf2sg7JEam+OQIX8tt9rxzU0x0INu/tA4ODZbb7
TSHE1+DM/nFRDLW/eg+i3JHLpE7QEEkYroYQUKh1o/rIo29Umh7d00wuxDqjsEx4wdu80oAkMTmo
Mdz7SG+rZurn0y4wcjWkDKmxpm8EE6qyHlTz543zRi5Clk04dN/inHbelre00xmRG6dxQyyzCMop
oqd1mtQx7LEVz8Q9FXJUtYLMr1+suwpAfnpMF5G6qfaZmc8Je7wHnjVnSimpQFypomYveYrDzw+Q
dzDG/iLCgsb5lhFF1TrAXvdslVfj0eezKb4NwEiauPbTGwBLfcmWUsgxsTLhuR6cqaMwbQ58v57G
JjMACKtWfBafCZLZZEx5ed+iJbpSX3RsShDReTxAJT9HNdf6YCXcQ7LIqA4BA0FbY/f6SgzQuXgW
Qoxq2RBvVUhNrcr9fgiXuQK135eCUsSZ/96SdoBaeoC1HBpSXSx1QSmM8ileIdGz7QOCZjk4/3P1
eDhNowVtdLGGumtpr1OYahTWUpgzL5z+Wa11HpU09X7ZbYs/zKYdkI/m3s2WE64Z0rbjB+XUJVZ5
aT+lBbB/TKywlFZ2SpzxhgSnknrgWCGc1HHJNe8QxQH/tqY4ckow4XQlwQbnme1/N9TLjKEH0/wm
XMkI0DhHfn08O5H/8M3GOBIcLUjHJlfDeXtkb2obL0CzR66BmKiOpU4tge/YX4YYJS7XcyovWi6Z
5g4QiNfSJ9n2LFS9sCn/UEcVUeZLGd9OIX/hLmu9+P4L/L+YvLqeSCnyWKHbMG9pce/Oqi9pQS76
P9t3wFpjgIYUCB88ViJqzEqRtqIxbfl4lVPY3+QSjn8mxn695UJbvonev8Dw/+K4BXYjTl82J/Cu
Zgn1aA7L6jRL/oFQsSN19mYAh7daWPzPLwMEg7weZZ6v1f8YtVGsuAnnHuXAzXJvgfnq9BBL/QKe
qc3SkxcmdCVH6tF+knvLaXxsEnWXGjMUeIr5+3OMMhqSon6Kz1R2ATHvxrrzbbJK4fYQZ+lxG3LI
s4gnPXTXLqkEccr6DslS7ISRy2soxic0grCrXe6jYax6d7xYCjOvXXBn26aR2CL3fepajtEn64gH
SQW21qWPq96lo7el9+dpSk1WTGHNZMRWVy6M7tp4jor3HSqfWXmxGXHg7oNJTN1KbMs2JR6puVDK
+Lx79TIBxwUf6kXsq1MeQ3gsXLqw2uYUEcKW+/4PbQOaHlM+qRbXWUnWvX1+E24rD1r5qkJrW0/J
A6gsYjWJLwI11JiH1S391IfbJRMO6/wr16cw7VsaGvsW9EiZSEEfTQ3r+3TZfOskU7Mf3HSLLAsW
+HPK+rLRQ3tZnyUokj0DzDZgSNUfJs0zLxASih0Cf/K/5xaN8pP4yKVxpAPtKJ7Ie0KVdqHTQW4o
Oi8vLcTwR5ZbgbPPzMOlkwxCl6WZLNsy9QGxn23NxpCPBuGn9Gv3mmjIop6bJwuk5FScXjtFjCpX
IoOTJHKp2tczWKgOZl00vgxlEwwGwAKnCkLw6U46gM0ma7giVpcjEh8aHsNTAXAkJPeA1QvOvN0w
V4ZToQvU9JqNm6kGDazx9HMDnmWnxCn9Sni7jYRT2XlOk1s8RT90lDNsdosbX6+fpF4GS1w7jcRw
NvsotHr2Fm4hUxDwFnYEMXpPlajMWJB0iFCFv2QSPcJokBC4D5OpXN/bmDVps/ZZjCmRcJ3aWLJl
+3Ca+hgqUZF3x6pxiPLF8FBFcY0HcynsBx7ufv3t+m+4i05oOkI5XEOm1U+didCyreEWWWKRnv+/
WdZdns/WbQWdPuEzG7PujWKgi3nJhUIKpMyGQMsPfgSLdQJQ8HC4hsV+YQeuWoLdp8GErYCkrPdD
Y0QvZ+wCKiw7sxgh30ambuX6y/eLMMzsjySM0TdCF11UmhgAi503rkZyTtY0nj1z5nzwXBrZOR2D
mBFjkzJPVrs8vjCrDKGnS8w1lcd1+RGFAlUN7+FtFvc69YHVBrC1rIsFAmcsu/K4S3FxqgvyQ8ye
9vstP75YU+fskN3xrXwBRwo6uDPrcouCMojyTn9phuxxE7WcKN1yXpMvXW6ILGs1Bhd3N7Fy2NP9
jSvGshdr051KIMCv5/5vZ3XIE0/Fch/rWs3ZFarNpmaAGY6weAS0TDcIaC6gNZQikjT/6BdiF5mj
0pKG2dQU4sC34upzn/1kUNvT4cnlqH4UA+MP9xcccsolWMqT1BOAn4ZDVfUSlMC5zhP52SeGtI4S
o/xZqOnx4ziiu2CyHLHC/T/vJtnyvpW6I4uun+4gMJf9r0DgxckOtxp7OQDMFK1VJzt0uDAukNCj
3TarzFLXDjUtHIcOYh134cpZeh5Fgi6pAOfudO5Nn2P/W3G0pqUZUN5b/qJYXvoC9yVHXmUPihZD
w5yAJiVossbrB7Y91FXYbTcmK4ZMW05sGK11AqpCXYeYDHIp/5VgEZJhu11dOuCTU9LWtBaLHqry
u8CQVUiIEeFlG3lf2/Ji4aFyI+yRqdVql/Zy8FZlQXKovNGbEZXQuuRzm92vOYNjWsNFHnUC8VAa
aK5/l6pZdg0jdR9OlEhVmHbdO/c/bLLZs9Iwr3mbXW5NoifBEkYwQQMQvDOh3KusUOrZHujLd/Ar
DEMSyvhCFxg9IfOrYGnMhMQPwqmi8gz9Wsl5W9hbkUvPUFNxvCSu3m88lK0FTCxVcFRGlZXfYSKP
kxcUNsL8Tup/dDjvNb4zOLcMTQJJ68l5yzBBPJLgsra6G+wsEDN2Msw9uL3vS5oCdIfEUNfMy7RD
q68suBIvWzlF1WBwE8VhLlFDnwnCaw8GnFOmgKwB0FbrW9tPEQ4sqNtuZ66u+7YoxR7daGc3X0OL
GhAHY5LcudC/ALMUDbtE2kcDDkJ/nYHZMZl0co2rdzRkXq0HX1OtrmaxppkDlKjTdwymaESmJ7Pp
DgPlsMUs6e5b2A+pr11ltJSIkqgkoKLzAAOOq5Ea0wGd89Ntkm9o7WDoUDRTAmccBjnPP6aK4wVX
us2Uy0RTzmXLGKbHJ/5jZ+ydwZqXdiUVu/ZtL7aSHHEHZuPv2InYrvS+50uyUl6XaOcFNoUJslLc
lG9tD2xgafVlrbGY5iVLlfN709+MsFXxanO8uniaFFja24bcwU3fHIfGl58PR7jWeFdmVLXbRCv7
8DLJS/OO577t0SydNiNyAn2kJSsfkvUeih+VBelYZI62qD7ne99HNf4E3whrlH73dDip3JlradT0
yGrzOByWLwv52yWztST5acJux51idxFb8SAntqd0qkJD9egCbxrXVJ+h5ZHfhdH+N0wGD7UVx/QK
dQElrgPplNgwIH6yBNJgpDrg/VGtDAkZl5U05Tu1kysHxPB9PMjWnKKKHZ8lf+93Xn3pYDnyGvzB
co4kkQKaj66GTbaU6z9kF1dRtI34C8AGIFE8QliF2B5sh7IftHmecusjcMXQ9waxezbsIz1ec3hQ
8ZTpBvJyaevvTSpp4XVCuV4v00bUx8XCTMj3TBnGRmNPc6zpn1G4paZf1MkFw9rnMd8wcZP6K/Lw
sim/UMAkQpl809NQTyolMd2qFfjSFfb60BMkRGeitz9ttie/Q0LxeHdnNCklhdx999ZdrE5OufhE
cFJLie4Aw+qDXtoj/9T3a0Oe5RIlgp80xnvEMjUto2xbDVx0ET9aicb0ZPhXq9XPNwGCBNReDR8+
5G1bu6wN0c+U7qntOlkSgZ5jJ28Iuo4U/6w1tzh2aLcYa70bv5K4fiTSiMo3BhXdss7pHCUa+oXX
0b6V4CPvbYOWjz5B1xql6YJNCCjqnQFst9iT8sTbszIypeYT52ccAQzY63YoB2vtS0+Dpm2X/XF5
TbXPHZEkEOnGpmgJ0jnUUgs/Xn3iXszw74Hwresc4lLnhjxl8FgWITNb5SyCfQQNy0AuWYIjoSxW
MM0/xoybSclfxaSCMYpVIpxmZjKUb7Z91e8usdvaCK1nxfSVSwIihzV0Yg/xjBbQz8k7e+nByfmi
Il28JRryRv+hHc6fhOkoLgQCb16Ya9k+phcZZmXTiZUb/JiZrqVs8i/b9kzTPLPQlGi7zVH4x9Qs
tEeA1J4OrE393NCZrMgtf4eN5zlVsYwtijxRNphDgMrndRE4Tioag2+FMojyOKQfPUHk6UonMr1H
ZPt3xtXH1ahDh8gZD9tfVu0z76oxTbKLYulpppBfl65chTGMgHNY69aGgjY28To+iHNIY07N+FuX
p6FNJGuiYMeUSI36agZlCKbdRqcJDwPU8rgQDe9IHyYfMAnGFtOk5OBQQLi0Uij8trR8n5OrXTnY
2kVHPqaeIEJeJFHTadmlRfhgDzt0sPWKiPczefniEizvvsHs/H4B2WnVH+mVI9BTF/Tj/lsumx6r
mnxM9i9awlQx0I9WZ2oBskWvsl6FyF1mlHuq53pySPfX8F7rEYcacqRWiwqbiSkavL1mQJZrtIZJ
+a8IVFSPakd37/W9/Jwox23M0J0sIRJSKf8bNvFL8g0Ea6mJcwKWJFRA0dw4iX4yDhrFH81193t1
1JimbjOT/EyWvGpk0FzdTW4DWcmaYC5OvgrAduazITFrWBwd9fVAzSWoUd1g9bmjQBBc/E7t3cZL
+6Z0gLHm7EQcbWpdAtpIkcAIKoaR57eHEhsvveDH5bBM+iy0STAi9sfN8BtFvuf1NtmMTKejURez
+GQb9YAs28d00F15An77sY4ZOfsCzj4Cgqoy6PCaVLhA59DrsRqsYxoO4ugBlECDzagqbrAEbtsF
AmN9XNus1QdIF4JWqrfYlQXE1i7D/XQJNaoG19KSNRVK5NTAFD0ixOf44sEbSUQm46t7vNXc3EN0
S34OziqiRsn35osz8GpVhQllN4ffdH4h6rUz8PZxdcN85RxpdVKQsDLToDSzEctXZ+/V/UXuhiXc
D5LAeMGKAK2cp8vPVqKDEFJckW2LZh1etwNsM1qjdJJ3BUvg2Y9aLuZ1fubsiqCYwdSz1CuoS3pl
LJcTFRW8Eo5TDgExxgwYoHUPR9avreDB8jsccUzoaACB99jNCJuDOmdq+/Vr272htbTw1uQ2hV34
TdVAwFMyUo1MT5UP6FI7aHM3AEAhAhixp1YFCYxlPXbWVCpm8rcMO9sNxtTA6pP+MEB1FG+mN1UI
rBn78a57ZUX0/goH2taTTLozgubkNmO9E0nlpz1iyBr+a414tULskGAQhWVL2xiHOC//v9G3hnxv
qtJrC0kUq+1rVcBiZfQ0k7qYgtF3CAmvFdbrkkzznHr+A8Sk+i/gPR4gJiDwOnPpYSnsJdF/3nQU
Iii+1MryzgKazt18T4sBJvNkQLjY1Fm9etQPwZmlrwh6Di1LX9lGT/R4algUIZ9CK65p+QcUoflz
U/cwUE6bzhxiyB1vGivHD4ZM0ZoyH8+NqvL8KBJKAvq90iBuKxlrG9RjiYQ3mOU7KwJOTF9cWNlh
GFBfUo9W+Vi/E0esKP0p6s57Gqkx5b2QjC4IZeCXqQ23Zv+yDakw1NpWeS4wMKRlGMk3Hi7mNALV
BcgsZNHXVbsm9ah0Y0dNqDLFSNUQqWLwd/BHRVUP6jQI9jnL76Yv01yF+KijOQ+9P1HuRl02Pcze
0X+alijeYP2r6ehrBWHWVCcbRdIts50N4dEvG+7zNDubSebzVIcNeYihhufpwjqLxi1BLTnQ4H0Q
ewLO4DDX8QNzIqwI1aWxOE7YTRUbMXn+dKxW2rDkcOicTk5t+2E/SsG/k7xv0WVhAEle5V3GeXzp
EzLljOSBPssRi8blUWtKFHj2qpbGuIq4qyffDV5/ENABhWStU6Oq/Bq4Mfb2GRlmMfdxtaUCmxQF
NF7li/Irjsvye4tFcqwh70I+OQn41xo5iIM+vQIeLmiW4huGD4Rf+0C9/XDtFgTofloqWmMuTX5X
jkuUx9LXf9B8ixVWIxnBqAE9/QZG5n/4XN+3DViwt1tKUbF81KUpaa59wQ8eRMCNDMmX6bQMCZOA
jDlZ3nv57O7cXxOjCEg6XbuoddEyfDEeKiFV8gsknonlHBW6Y4tR1TvWLyj5swvnTYcJ5dWwCo52
Ltoc8mVh11fLXTFBt6gCMSW7td/cntPzkbfrRrQzcFJYWDmbk3yG7tpOxBykddWwX88UD+DcqYME
iqj6Ft1mxqXf83Z67lSFdnzJB/lV3647l4m2+spK+hVABxuXPVcoeNMNB3G6tYdseur31999DW3C
QtxStP6zAK9Mp+BJ1Inb0b+1pVhMD+uxcMNbOmIHCsFaz9SB4YUwhYJ6EHR7jUUB71/1CgV20xpm
qqMNDzxU2mvbDZ2+XqjoiAQ9jSmPErPlYtZKSSZaoalv4pjsPQ9NqOvKmYPBFz8FfKWqCE1FP2zE
OcOmRnbmzSS46VYifip6pYJwHq59Jm8DcUb252uY44JONGH9/iJcl58zdZhuX4PPN+xo4amoz78q
+HU1viwMJ/4ocoyp/E4UHwx0yfH3NmQbmoo0FRH2VBrJjIehTHldUe4ij4DjDpMnN3yPkT6BY/pp
aTDDic6YrI5E3jMHs4guiG5GW96QM1QYnRhL5Vspg7to4DlD9zghFAQ7mlFtIXHuu5yhl3TKQLbF
hgye01gYBu97OLEZO/euPZfswRaOsoLC2ugVm9jAyjMl2dRhDWlJ2agFr5upVfgBdN/z5XKOAvGO
KzVDpgO7n/w7Z4Xop4CQj9xv4ZtifU7a2y4LHZrU2B2Yuqyj1pX/3758o4z9wAGwN3JAVa5oZS48
DnqHP4Fgwlv3Mz3bgeZuzD7dd/Uhw7tr16DZbvvcseDRQGAtbnJQqybTdiL3Yv5WJXkh+fUzDzyb
vr7e16PW3ErbKX91e9ap31FecuINFNW1Mq7Yc2U/jh1Ankha12RC6Mv7mo4iYOYOewzVPdUylk0v
ToK1srg3r0tS2ADjjniU1qwO5nUT/MC4FmYcqEmYMV63cDgn7nNTGopiv0tyx/XYlHE8VlTrI6dy
JpMD/RkdmFs8ltlnJFSUi1e1qL1uMQ4tMJfkHr8Gj1iSJPuzoYpwmbs08oHB16KF/fRxUeEeSIaz
HussFWX3D0EjXGacqLPcz2y0FnqWzZ0RfcCxey83x+nODLR88vpfDWSd4sw0Ri3mSD0bih8DutFx
pGWAJhN43W72Vu+UtPhQdn8xyqyTo4l0gQecRXtv016ZxO43EQxYbVdsDa4g7Fnx4q9imsZB5gsD
WzzJvMYr4lJLYidUghR/xm0/rTesHXxXG9Q1fODEFJX0mKqlG8VfpWJhQAdBHtBKGYrZAj9JU4AJ
EY086tra6JimJ5jbW5+wbKCotTps1zVjTfOwQ4OrCxsMKdRIB60VIUWa8hyKJUzucrYz7/C+XCu1
Et9oDnZMFTEVN+netytxgFF9Z8EiR3QytXlsGvNcHuJwcBsj1RpF1XLG6+qF7qvQnA6wZAWF87iZ
rjoxPobrc6cAQfjC0NSQpZ+tkmMAZhXd+JvFO5WJqM8eYQisFmC4hktzZv+W+9JreEE9Vj40xBX4
nuNEMINkq2mzm31cTaR1uakBZLGHkVy/i8xAmSdDese7PLZC9Hp3mjTeQbKBtukze5R4H+6baH8p
41YE9ll4JWaavkK3k/VMZhsUmxojIgWY/lM02ZnilvmF/aiXeR4M60aYXwhBCPbRTBdzDg6OhNPw
ojCWyx29lzGT46Yy0d+W2dySRk1A3GFEJ9wjzpMEoObAF6FLPzFBuN2v53quHayuMW9WfW///1Vs
BwEWePJlRIlj2E7DAhpkJQsaU8O0z4YEAUvKwIKSo3PJKSvhpZQK95sQE0NsZJ1aUTpvFAMRriaC
e30ovGqjbRJSZXxV67StgpX4P6pblHBvP9m1jjQJ1RBSfJ1YdhrYT68tp/b8V9dCAMLDRS6yc/H0
CZGblIIcyEE18YsF/7Qi88gfrFxn0uiEy+QbtvNzbjNdUyj3TZOU2Q5yRVf8iS/7UDf4BJMvZow5
L85OUOPZ65ibectk+8KznenR+mU0Wo6a6mG7BaHjXtKyK0ptAESTQW1tIfy8k2xWJ/StddbbAeLX
kx+LiCzHprCFzhlbclUEgEOHmUujE8edSR5Apo66gcQQXNxCrENY+cuUUPBIAWATMifMN+nYwrkR
QSmNH48y/6t7sg9MCn/GGv84ty1DjeRZOHH6tZbp5oyTy7Dtqd3n3p6npjLksKsjFDt/aMlwOrQJ
cDG5IGKJpIsw914HXZd6EIJlOak4CpdruXOFtQfR9tYkmmDsl8ytDvQem557+exgwjf14W43pU6R
aO9PMGGdg+pQT4/fQxk2l0C9zJt6FOQ4KYoviTvnwpfaNJVDFf0WMp8+9TA6mvoFbjBIFi6BtWK3
/ODDlSoR2c1RwkCXs9aGP6qdMXqRsQ3CTWHAHE1STz26D9j2asET6M1IIjv31MIZSNYSZUaM5d3I
Nvmwgqnyqr9yrGzGwIcurqkWhexcKU26dpdvuxDgwYc/zdKOoYIZkPLJlVF3/p/RUjO2uBLz5zZT
92185zgTPlZ8TDQCAbmPmG3kJCjKhpl4iWp1MBD8AKJvmFoPLBWIQSUQpwbiksMGbglNRykRcK9d
amb3Z58r+Z3W3YgzrAIHhlEpoPvmWwc2QAGlpJ4c73w4p+nNTOFM8wynLzX8gNpwVaSSXRhaqsCn
KoPiQ27hh/GKFkFtsAFg3njsIp86hi1l+2Otz6cxC8FV7r4PD4IHei+IDKu12NGkJJMTtBMkVzVQ
rSQhmZkt7n283y6DzhTeS9m2zUTZw3nT0xKivGdnn/yCEef55AJHXZ8A/WUrQIFxscmDZXXB0q8F
aeoNffDJx+jfOPwTcw9/rr9Rr7VcgbKH17FDtBkQk8bpCWy4y+pTUtHTgXBFNymPJ6YOknQhww4a
PI08nTb9HoMtJyRIi0zoMKv5PVGzFDTBaySd3ZJK9JvH261ret8FgiUJapqqtG96SEB3X7Fqa1j2
7OMCa08xLmgNrxS+FuDjK8/p3K9Uin0pSbS2+ryXLyAPQTiwQC48wpZ2TUZOxepJvBjIVVW08hm3
vUaIbVqgvjWCPYuguqtGbmEQ4a48L6tCXb/bpdh5n01Ay90mxjolHpC6PstIpQAQ9DrU5cY61KUk
S/I6xp9AyaaN2q4KbUAGAK4l/1QdbSnqHuaeUvRF5+0mF2MXXcqqDmcf8YQaBPCORDLz+Ib0Jx+V
L8NWvYdE+SznD06rwXDC5o/JaaSz6CRCqgTLZa0FGwZ597o32WAGynpzEiNhSbvIBbt4y4Y45mTN
2Lxn/rkoFhcjIqK3pgHidwGbdRR1ek7+AQT4syLt8veinc1JMewxvrSF4grQ1o+CuMAAQ7JvyYuf
0VE/BCT6kZ/E/JVlYIXBByZlTHN4Ctq3pmh0q03uxnNJeVe346Qj2h5qJa09zs+a7YTUwLBDc5xl
wEh9Rfc1Vt4XkvAQXAe7NJ10h24GJjUQfjaFLRSITIq6eifJD5P9feq8pJR6GBV6PH3+50aGEoax
4k2IFSfS9NJrpbeTUCmYIJzsIVV/y9xR7ux59LW45qegYTnaeWaBoInh5MfvyoeHS3H9tbPCnkJ1
p2Yv2Xk6mkbst/rl7nniFWDHpD5y5ajNAOObD2Ke27bNCbIos+0M/f/TyHHJH/JkvNLNVi26acRG
JFkBv6hETtfNi8Pj3P3idSYdBgpQRp2731FnLXOHZBJ9keb46IRttkDvWmnrZIIQK4n2aCACFg4x
ABwoz0L3zwhXsTO5xw3IqojpLK6SyTWNGB5lyJjVydjSGqrkSs3b/sQXar1ogC/w2vg2JHWfWe2w
UqC06nyYEh8bzWQHzT9Myb9uvdgrUrVK+VqXiybyPMzKtuuh28F5td/8Vta36hIiNMbDNSEGK7NB
8SCjINzGwWrIYiTcEjkYB17QwyEi0acCbQT3/RgvtX2SyEw1doNSiFdN/aCjxUYmUo37b65Jhj4K
jKhyRfBXTg09eQURZk+pzBDmdt5fZqEZXmzOW3BQsyhJD/69teg/qJsl+5L+iMnViXG/sSQ60X3S
bVeEbZjT7Brpqhd23ou7nFjSIxKRWVjB3LXQHRoP5eXh1yRoGNPThq8Vcu6eq7OgZe6HI17rfQLN
NhdjG3fADuHtU5JplVxTLRBUc7NizvCNi3OJ82092FrTYzzq7lZe06JUZOdl+Mu2OsJbeaXQ+MI1
Cku1sOlNqJVX018U87BBtJr57TG165NM+SicwdCCp4sIpTdHC770J9JamrEUSl9ldxGL8wp/CMQu
33YKEKiwC0qVrE5tyb6WxbgHJivCCj7FqnhKwEQoINc4CZxmDJU/gs8pPkUq0XIGlRoZo4Cw3BlX
PztneeCDQvdv1f01i3YiqWuCMIBQe4nbnxg0dkTS2QtpXF0yYyVbvgviDWxcvW5oWo3a9Uk6XukK
4aLpYEeMITQG7a18gHYpYoyIkKghN67F/q8281ZM7tIYW9upXOr8rrupwxAzNV6um3EPYIGP3H/S
RDvlA+B3D4gfILmBIJjSuj2P5Uc49eJK7p1EsZ50gym7UcC07p4Ch3iuXRL1YvsN9doQq4owGoSA
p+i6Rqdk4yX+IILhpHqzt6wT3vGQXia06QDR5ftFjLY2m4dFaxBeevmT1hxOAWpl5g2txyHcihjI
8fiSN7JqAflvOqMC7whzJzqUex21ZG2QbX1CHHnPLXLsGNSBolLdc4z+jmL/O7BFH/nik/lwtiKd
Qbvy9Y4CfRfDEleqsYKic2CN0srUEq7mbFP5a+tNnfklwlREe76RgoL8nfXtVl5BZdG1V46bJbnn
sS/U7V9ClpXcy7pUEeWV3RDZB3+SkqyrsgHgDStlb6gAjtITnQK1dhXJGV7+Yh4zJSOMmLPWJsrb
7XgUtwDV18jaEwjY7wd2cCk4db+k2hzWT/s9RKRslLEJMlU50U4axe5hfJswMn2QqHUhBEnadaSI
GqozM8wREApe7Rf9O3nRpj65wpoN+6rOqVwG0VOYEf44Qlkh0UBciBaPi3Jdk3yJdsK2Xjj9UWZP
k58FUq9iTvLbmEMVk/D/HdP/Gx1uA8WHSvKy0PmlDDWHImcNl/31KVyUhCvJUcuYa3bdoZ3YHSkF
n1P2ryl1V1MW23J94XGxeU+8am6WWC+ucqrtMOtCnnMuASTscHvPLUzmSahlRB2rt0E0rpQ+tHbU
ecQMps8jcGtpcuBj+aXG/YI7prQTlLH1ythYwmNrGMJQRTCwB8Y66vd3szUyQBo7ETumnl2EfQYb
1XmDbyHJXX8eLEE0y1QlQNgZLJ1NHYW6kh7vUQaO00WYKy1I8FhFpPgtO2WgMEjC2XFoNFsxTSUa
AwOcPkEqfRtS9ofEP9TUejwTtBv0unNtUzPal6t6ckZsFU2Haz0iWkRddZX+syk6WZp/1I0odC7r
2e+4/d4bwH+MeNi3xcWMlY97FFToGCGABEkmAaM+asARzuxVDQgqkJrFCVNGrKXPIEb8+U/spfWR
uwY5lJ4dSswf1oDRZbpFhVHnz1Hz9yEyBmKVyXNgJLiAOIlaKPuKmnlwY3CDP7DbBQzk6bc7w6Eu
DSkvJwFrzQSSyr2DLMIzlvbQMaZar0/kvtgEPuM1Ldrcz3pM3JXfW29GoYU31JA96Jf6w0XhuvxM
RQ19vNE1GzjQwlgnHQ/nAqga7KfQSwL2phrdQgHgNI/y4INxUYK7k7wnwVvN8DdvMFktQR9G42kX
Mj+YJ492gDAxOg2CZQm/I7yaH2l0kyZGkz4GiY2+2OYw+oCtYl4BRHJApX+INnVKLPR+4F+D3TDv
QcYsNA6OeymnNq/vrbSUL+dQq27K59zIe0dlY6/a5j62V0ZCnVcxeGNoIqPFYuvTFY+gpZBwNy5y
m4/NOhu7fBB5+7+Pc38H0tPApq/dYJBT/5uUV3ojWu3vtAVzhx/SfHOgaR+W6NHPOYmzJQWhzYv+
88vet3/rLiQfmfwLgWPP2Doz942RV+QrDZjpxvCeQvNwI9EhC/CiZypUZszwNb1vV23yTpUxYO3E
JLnMuziw+Ixbvme72NSo0GB/fO4lxB9yvNdQta4e9S7U6/eT54htKk0MwqaamySGzHbwWFFvtckZ
Kv1dXlY00Np9W3Ct08T+t8/Z9YWPsSw9XgmlesI8avkFjIXP+ZazbF7r8sT9dMUJwwiR4635T9sO
59W4op+nxqRRXSgZ7fRE1VIWCqlSZsVwV9/6i8/2KRhnO8NFRUtqT+0HnKhUXlrHy4Ej8q2azI+U
1dBdbZBv5Qn1t+eCANjs0p1jc9J3w9RBw9xv1QYUD2KhxCLDfLexzdZKu12yJgkGPokTwVr4vyyy
qFYZt7zhodvuifiiVq8aLvNVFKSOW1uK9OEXCNi7gF5FY6TXxiOol2SiZOxJ2J4RGjiJBLWdcwt/
NU7Sw9xqOGMhljKOidArNFgrw1SgtCQSj59/9CRdak2ZB5rQ9Vs9XcQmxcGmd5GOQW1d77WGu0Xq
njg6wcryuEAUvPosZJs8CvqXOooQ2EJKUtMzKLQ8QtEhEsFQawe46RZkpSStOQub/tO+Yi/a5zD6
ITDQ1/EriBvE149o94uQZHsNYyy17uduPLkhf94IxtFKO+6TSt716RrXw5OnGrKuRv1N3tHeZ1eo
t0tlTA++5/RwOQSCoAkwxmFzqNo8OCQcjT+TGxV/yZBtOhlOmpCr+DyRXPFWxmUb+wXhYKFSMmvz
qZnLsfmQSX1UxEYdrkEeHaq1QqTjm3bVIi7R++no7VWZ4S4xZiLmS35G0LMKKieWha9ENl7wFWJe
/dUVUYVKH0XCjKdrRdStJY5zFM9s2013X13jmJufRxTVV7uQDmGpnJpMHwew6lJRQoPNGUjPkFtn
zfWE6cKB71mjtbLFFVeAW8CG7dc9juJErksBohk768C/n2a9IdH91iI/dDr6Rovj1INfF+Zognz8
kaMTAKg1ss0bD0x3+wd7uIrgSeyQIc3qhKtH3rqr3yMVqn9gPzniYYGVw7C3KC0ANP4d04paHEFU
9JMYBVZCPy0ZoZMpthc9Cp2XyUzZSyQMqnEgNJMV4f8xYBiox+GC9/CXH7GPGVfk3Q9WS9Qj0dUK
sYW7n4SPqQUCUriE7WCmj9KYuP+Dgyy2slguyYz6EP+JoT7+EQ3ORdcrNr0RCouw0hpW1MNKafk/
/HRb9p4TxMvHDMbAp2wgmOX+vn6SOtbMuMWPUwePBGLf6tUO90y4ewT/qvi/QT/nLXyk7ptiQmR/
Y40NI+w/mfrWLhy6P1B7epEJJ4cBpWEoFjVP9SnGB48ntdhFtSOYoY/CshG1XQKsjWaf8qnenesw
jqKsnk7kcNSWkgfM1naVyYxkoJjwvSWswUZTCRz9jNg8Adc0y68gS+t2jFL2zWW+1GIXkB4tGaDY
cZDfVp5gdC8gUVPWUdLglqOyyNhigavY1SjrwIvOzpongaSuuXsYyXT03IlVma3FSRzS0iwuFqG5
hEQlhWpwTAdNT1q4UQGHbL1dbj2/CBBhzaBXKje9tXJxABlKamgFhoWykXUlZHaojtkWnP7x0T8D
OPCj5xH9UDfeus2L7eE+yXqcmXAKTlleJJXC+HN13k8X0IMfvbqsSN0hqazVWViaE3gdj0rY78Zs
A0ND6pse1hvsTW6x07houk3mHeMIfNSPTaZ6VZGAcS77jfdRu5EjWfNzCrU4g1dGBiNE9PP2era0
cw6v8Hx47O2zAklGeM8VZxrcHxuF+qwvBhvlcEPGGbEb2edT+Tl54YpfOuwMChlsFFuzpH/ZBwXX
OPnxkPG/cGjb/JMy8t9D4a5Zzdfz76apf/9mAIv/Mjkt3FDesr7C8OFNhBCooAJ6i9yPssJTdIO9
5TBMLKJstA2Anq92xheBBlkMSH/9pIfXkmewEs6GyaQpb1Al5+mm+djSLMlI9qgW5ayp95iEfFeJ
mJgKB5miiojIiDX+wR/1dXMB9rFAsVuWkiZa+w0asRPurA1aMqogp5lEcpaKacL2tQNbziqf7tdi
hptJxb9HLIUV4Mu84yCy50SP3R7W3F3yLFUCnSWFxSArRsrhCgnYHLtCXDO1pEuHkaeJryXUfqBe
1pH3jYqzqJ4x6Ib0DreMn9M9b9PJREVprRjLvOwZS/r3ykYjPuHSh12hdP8w+0ors+d+/GJw6EM0
5D6MWUF0rbwIr4pEApvhTvpKH//NOHZJG9P18XPDYkJzr3FdW76UPOUulODdl+IN3+YmO9z+3M+9
JUb7msPsAhZiRT1N/2FwVbRjMPbHRaM6Su1U61ESGqBuNqf3QdjZd9wT1tYd/kZ31bGruvLRarCz
QQAEFqleBq4D7sZ5INJKb0y4q3H2nLCv/oHZUyhB+xtK9iO9cuTMgT+mBDUrBZGd9vyrsogPqhrT
5H0wnepBF2x+wgKVDmZIlJMzRZonOnB515nunnqxCeGq4SrFXf41g5o2EjIIZJ7qPOpWl6BvjOD3
rBsWLtCzFxD70Iq6mQIXNSKiNI9EoRqWhLhh9giuQLquLjJI4AvWeI/7219cQ9wvX9o1+RSDPI8d
H/DNH/YVzxv2Onr0uUkOBo5zbh/ZWcDbuh2xMrh3tFb4nlF/91deB7coxHAiX1Uf0uFXD/i+WRA4
qf6xNW9j6ApWdfZQ85zZAWVXT1VGWTllzuK+fnbOnTNeMNuIJg1eR8TSRTC+aI5fDAv0TXMPg0Ya
JLPf3ipsTINaxexPlQ3xvgK+AgeATPQ1gSJ0tW2RrzfhGUcjoqOK+2t14LkooiZ+FbWL0kss+0Op
Qt93R6E2oCHaOPcgjh1c5T0oGK9xXAdr8QDpmyEBSI0LG3hyr4S7svojI8khJFGf5HhkJpUiI35S
o6d+mpJSTzeyx5GckUgchesOCoEAkA7+e9W60LzEVMKq0Zy9UDfYTLoxrd2nVLLip/fgggYxig/3
lGWWzAQziymRTnVjuXe2L55N0cucVUwggqFh7/rGkyHxNCdGyaUp9XDte5Ba0d/6JDw/bbyFi6r2
8z03O8e0oKkYqOTgesu+zoaI/LuzHzetN6T11/+Cj1ypXT/vgbkx1MMq01C3Sjn6vcuT1FQ99TnB
pxm1G4+zvQ8UcOYB024MfwqB6u1Hk6wxTcrokrjplbqzZ01EoW4tVfQ+1kqmuJx+r5jrqNqSlYeM
F/OfxFfr6NCOAoiJUTqW4VJJ9mgKZE6EqSmCXPgqKgF4tdro2FeZ+ln1NqgST7gfRU6a8xNC3t7y
EK6rxAianj5HxfuxIuxhdVGifGMZ1tBxepuKzrKwUX/X7dhX3kA/7qUZqNPypV26yEPpUCDoInf2
pFt7rUEM3GXxLR1Nzp6wUnrjyoOq8CdSP1gQtai+VcHvzElVPFi0l7gu2ur1UzJ5eQWwwlXIRdnm
qvyLaCil+jYqaULvvXpZrmMP3qJo8/KRBsLDzCrwzP/i73uOgt73YbSSxlpOc2ozhFQA93PaS30t
R9PZax+LydNjWSbjU+9MaY8DqlsctRuwG1Ufd7PHEjItLsOekv7m7tsW2L36F6UKJ9bufCmeksxv
+pFl/3C8vsyTbYAXDyNYJyLpuBUdUgD5LulI6vuU0rMWpW5c68vjye4s0nQbCA4TsS2CxcW/WRtF
jz9Xa3tod6uFXUz4wtuJ5hMKEYbTEhZz20tjkWPdRTGBmIJtqUUndAUMPKHnTCAzm8kiPk7221n8
jDYL6fIPYoQJM09I6vH4kAjGqvGVLShRWaBRb3w72ARmRPMJTspN/Gg62Rr7Ybd/vAr12LwnLadX
zX/86vOqyYZ2GYK/atcNrF+y0QO3KCWNBGYbS4QM0rIHtCeox9k9IGY7VMslv10vzDThwUVrua5S
E9ODy8rt7yyyVGK7LwvSBKdzKdj77EBZxMBsxbcW3Imd94OV4fBtcCj5+nX5ZCwHt4xFueotYepc
ycSiwUlZR/0Z7blm4M7rQb6OxkiDuxbBX4NKjLB0H3w47miru2iGpVXg0QkvhTHVtU1iy6tftp3G
TGfpjX0EWS4yItTSzyUETb+O3yh8czrdbJdPSM3WcInxOyx31JuM0sbBOCig/a0GV7OOOOgEHFGu
qe9gzS/c+uAHnzgAcoro/pH5bxQvlHYqOuViPMYAC9YzQnV68ey8p/3wJLOUb5Gb8WuFEhehPlsD
PKQ15RD7jvm9VsJTQ9l2jVt0C+ry0waxEhkU0z1r23l0g6Ewcfrn60NeL3fLm7/mAk9x1lxUbHwa
hEIQtWl+q1sqialFz7oAwbeGHsQNsZJr17yIlmDFcHEuldNzjNN8q+fZg/MDxXFN3fKyGvkOxFKv
U6LkIrfaAYHm9LUemy4yVjVPqoj2r9vCkmy68cDFBbmlQpmm6+qtqUqllt17K8d4xIP9JRSpq5i6
nyswm6jyjHB/ezOJv30vxdCHGhRrCYtB0pKB80AaV74OJjWdKVf7/KOtpbYRJZzULaPe0TT+HM6P
z3IXKeqwCArc98+sgGXtZhtdTq/r2203POMUd9Fn5dd45X6YHhwZFyKB4HnytJEt8C062YHQTjub
FDz8qTVDZb/K2cGrtpwwubvmroq4snOBQmc4bPVoUjBkfFlbckiEcpYdzLeWDqj6hgmQe3sejjJr
NNG2BWlXNQt5T/58TImMVZqs95Scvla6UkihB42xutv+tHsxEEPavO/xUpdCN//2tmuYwlRyEpQG
lsr8q64SQ6WMSqMBTI/Q7g1xFDDTXwv1UH1eH631njBHztyvZzNYihqGqP5qjZTrhDdf1MDiJ8nJ
h8trUS+l8zGOijrhjOk/9cjAMf/JQnoW9G9Y8D6cz4IDuZbkU8SAhMFMm49pfnY/+TRQOqaIK+wP
lKn/YLSHnsDCkxg92xMewMNaDOOBWA4LNjvS79GsFg6rFJWkIvFURKdzb/mt5k8rPRzJra9xaz0y
jELID1780r1aG3hEE/Z/zXmu+DHJ1vwMGYykR6vJ2RYbBabFB4sKeraQz1ZYz+BlkA4UIbNzGVIJ
l7a6Pn5qOu1xs8TAv+m9OhFvKMfENkLwzvh3dyT69gLHPrtpe1xZHlaata3w4MMY7FeW6+6sbYAJ
TcTPJqQQo0ZW7oljN4zzVfWfFsuZofawKIFyVt/yKH1t7rGuMBphuqbmuB70n1u4ZB3O7zEdo2ca
SvgsbRw7wFLBo+fzvKlhu2g3Ld5nS5eNJ1AfEQ+l3SPhCf6GEUVpsghzKOQjOeEMiTTlT4fl/qcW
uCYJYjjJV+onyvXW+ivEsnjDh48XEPB1dHr/0M1H3a2Sr4NHgq6Ewx1IpBI2L4MAebGkmeVS/kia
y99vQdWmzboUMOyStLAjQdH0a7s97LWp9A8bMeulg0SiD4oDl1YBHtVEaIhLh3zNU2cqfAexOvX8
aSQpBClWXt8lDW+X8QI8OYYu+DC1oG7TDQlRJR64yruuYW2nFIoHERWXeQ1s/rJp47+aDVPMQrZH
KO5n9UMt5HFWFIScBH3WRivkJ1tCEeM/ED+6H8UqpWxstpzzA2Ne7BUfea2UvgUlnumL22IMRVf1
WMmppx3ah3apN1G1A51pxs9vDBhh1lqMFkhdP56TyeXUy7g3vKnGNrs0dRNwChgrYejt0QtW20sv
6+l7KKavKGDaBSBL0CUhwNGlMlv864BUmu+06+PZ/5ujVfoGnwemXQ/p80T40xV1kNfYn8ss2NMy
fHE0twxvfIfX63+FjfxIjVYITJrY5GUzwY00kAP7tX+OiCa+bsSBarB9wz6lZrNWsO2ygf3xpypY
lBfUui5TOu5LPZBxuAgTMZDi1lorJm7PyO7sixSdtt+jJDM/4nf/zaQlREq7T+BRFS/c7J9n2o1Z
/AeKX33bSnWE5ibPTqrOn2f6r1/S/Y81d5J8Vq207gCh376cDeAQhuymyHYz4+BT18R6ekkgrLjF
6TjOhspqMTtaAmeaBCWJoeOMDdNabxsgBud7O+mZb0pfV5wWStg1ziXMwcQMzzwt3kOlvY3rlX99
DAQxZLXWvNXD7xIYM3vyiuQShnloLYaDqMGZ6Bm+yrAC+yjPtlY59jj0OXzsQvGjV2Ku7mB9FSib
1fiUuFz/cigpNY7KhaZ0fFwEi2YK2ob1u/hmvjps4tCq4YP0nl7zi5jC04gzvl7u8jJ5RGotONQP
OUJ1zcQGIUu8RKeokn1m4MHDyc46FXgDM560afAfHNmx0f7311xFu0IXRr0oaUkq3dYNa26I8bxs
JgB/iRoJ0buOJyx0RQsyGMe2F5JKhYWqKZ2khCTvUWZMVqJ/JSGpBHe8yobWolgxC63TkU0One0r
9NLdheaPbIlq9qySAwjvAIbFyDVkNLxH63Cps3Ic1i0XTmEmDAQJb3q7n/cyPZpK9UXaFW4VfNjE
C0uEWfUfyMZByvn2hoSnyAudPYu5troEbhpkcg5q8KcHJyJ+5s8SCP5GVbUqRfcoH3+G7deuD+3v
scVR48sAKcDXLyF5VHPdTNyZPGB/wI8WvtoQFVIOW0IPqlWe47kEGdCzyxKohpqarvRqWQMHKhJ0
MwUhQAXv/I9qJlnyEtBAKp/pjbuly5+qo9X5XFcQ8OUpS1a3/2CyuZZJQycsobXeSY4/VXGZLNeM
z+dbjfDec3kMJul43rv4tjq8vllHubCkynEsOZOv5b1D0G5omSDJChynCmdFO1J951rO8fvpECJk
sV3LtnLPOtI+pKTwC1uZ4Mo8kGgEUscILZb6muCjJsnEYDinPUCwD7EmVflDH6KpQg2VpNaqKTmF
ml8y0amUZmLxU4UUbu8TWIW52bpn387yWsGfWQSRHQya+qfhY3Q09y6VwKwrO4b1KL8QLhxPQXJa
5Bl1cJHf47SMsP385yPRObsxULjm14btBeawhcVXA2D7y88CrRT6Hsa7iph8zVfKr/RyNeISwspL
0ksv4NC+s94pD1BPGYO7QQ0qEzXh1QtbxsUiRAUbCDbjcojEHPtW/jTShqva6RdT52rX10TY0Ru+
iW3RAYlXBTx5gQHhuxuNtpo7PeLxdJHuLGBQomHNRuzfMdzeZxIGeVO7J8mwKfZ5bsOgsCay4KOx
u6v18lJI+EfFmKDC/NzkNQ1DaTPmcdQ830/uhEz16WxN/9CO/xIN4r0XtqL/eVjFc8CcwPpTyoxi
MKgz5E8xfF+l/2r6x8j2mig1rjZF0TGWbDmr5f5FARJtBLLK4unOLcmVUmjx4eXeWV6dlOKCHQxn
3Ayo5zMqdkyHjDyu/E5afwmmn7sSodWUI0VV9Kg2AiZ3vvy4OLm58zLYjPkWwKz56FQ1ODD5mIR+
st/mal4008Jj3Uw3BHlehJguNz05/hzctGAhhv8II+A48rtniV5qTiOOQGey8HuGNo7ktQY8wUnQ
5MaBgKEl7cfDXBW1DABttFWf8ReRFlOvZVMr2CLuunXK4K2EGwo7Um4kvEDRI8FxHVmzgfxL2apL
ML2CAjr2S0o90WqNwh8yXO88Cv9dla1l+dktzA9lYWWf0Qqo9tlPV0072DZlusxgYJOlUHgra/Xq
Y8/ZofOPh/PC0Fi+Z19F7OXuSeucsGMtQohH3GVuXKB2igG33Xrnsw/67bElHmAWalU2+ZVzMt45
yiKwMt+vTQcY8RKVkAQ/vqxGhhx1DVthHdHiCcrFJDT3G9+cvIWjnlsV+qYQIq8p0LB/V4P775Na
lAOwGA63kRDPwlYl6oSmKg22qoqOR8mCP6fqYudQKbzurpO7A9B6gaa1cZ8gRIaoazup0xmtOimU
qO3WXTDMz1WAqQyvJfgYKtJMTxcD7188tpl9Bzbksie65Fk8ggwLyjInfj/q3UwzV2LBPSXAjR1i
7nqp8DTF0DZvh4JV4PqH1DSdJ+ZtFk2x1VZJeDRPT6CE5u8ngSX+yj3oo6RWbDIFIWNdHvmAiDoG
vYJ4Nh+TJfEA82jVSEBIt78lUSzUvLmCCZQYaiL7qxY/A/OCHvLEQr9QTIKx4Ldut08v8SBP7mrP
ZgZ1N64J8ItcGtGzq8NhSnmaNyxv/pHJJDGxC+b0tH+P2wgO2RB4apvzrNSJRA1evH/ruIJ1gVu+
K0oGK5inRFkBjEsFOBJOw2aEGNi64PrTZMpI1fQAGkNu6+tR4LF8baJsWK0CYSTQbECCH2H0XP0y
Sds2o7uw47duMsihXo2oCvKE6T/vQBMkSTKMO148uRYeAw//YI3zOjTHExqOw2RlgG2v7qlxfNHO
cl+RMzPHTDkwlRL0Xh2IbZY5gvkExPC8+qUWAcI6dwFeP2PuNlRm469+nu0SDGk4W2llXyxCpcyF
8l/eB6kbDZAO75aU/xxM6POzbiyw3kKrtDf0MxOPtBh8BJbZo+A6UI0bzMMitU0XkaJLkyFfVLwd
V0A5EpiU+79aa5LpUaX9XICvrI1NSMVIh/ioRfRh3x38rJ0dw7ht+8qnnChEiINeAN+srGXlZ4Uf
L+vy25YE+X4aNup44DymLElwKySW6ygEcRF9P1mUchY0Nx9RVcS5ATr5+u3OYz07/RbEeVo6DsFC
UAgvMsE9rVoORrMHCdyhbqWFVe2x9Q2OMKiTW2iC4aA1byOuCDgCmWP/sXC7BtQOgRM+0jlgf5PM
I3LsjxDvCW2oHL7W6rxrmMGcjCdPC8VBKaU4K5PHctO6Imlz+eU2YL+UQ7dr9Ca0p5PZa5NNUSdV
RNoaG13wBLg7c4EBip5CnyHXiDZEq/3EC2ZuVYpnzK/cpUSUR6tDELGLvyqImHtPF0XUDwzhkqus
XRdrQXttj2+3/SYUzek9yekK0pq99II2oLtsDF6pA+eVIvygTnlOb8EoZN7C7jYYcr4sw3s16iHD
pR8N7qIj8GFLRy44ZNBiEmlPskV5LQUzf8eCzEZLZuXCyjtTcUqU0Lhc/Ke96ktKYLtMB2C/hh4B
a5dwPIaf2hB/emxzX3Lz/0fCgRLJ+jnWw/p/kI65Srv8m/Vg7fti0GkioEaEYcKQDa0ycKN1Hor0
XuZTFDr8L7ZOe9IQpu5x8Cr7e3FmGox3tB3nJpqtAx0yX7Th6v8vzR6buEPykAUNSDZ/ERi/9VPY
E+69GDChB9s//FY/7Jn3wt76y6KKtS6z66XgU19boaOdicH03SXA5LDq3yp2UOoWloy5OijDsS8x
O+scc6VvPEiXg5fTjpoDR3a0Tychqm43ktIFq0oGZyz7DOT0a8+dfpqR1EK0aiRfu61wyRvFEuLh
1P7kgYdaic4UYM1oJ14N73iaw2e5z6pZDEB06/onxEhH9BcrGRVsOVRlGbZ8ZjRd0XhR8VBVzm93
oTlIuDpoLv+mDlh4r+UECccxl5s74+lw+Bl9InvyRn7ET94qtjPyH7leq9G+zAq9jeK5yVcFlDKs
UsP8QZqGjZ2ZfuyWnai8G4YQAKJ98pU07Z9jiwqJhPQ96M+DVSuXyxf9RfYzpN1TvCvrfORVvqkD
gyCMM7fJwMRrZKVetYU1HahZ/USEzCHeRIBzvHlEfYFxhH0Q8Als935/QW2J69ezMFtWwcc1EGpZ
LNw+e0/6n15Ol8HOnWPPeUEHqL7KDsXap2uj9n3InL+qfqfTOmS0XzvAayzlA6YBpHc/gRtZUQyR
crhpRFdz1BV7Vr4zbB7cFni3bJY1BKf8ExpirrkA8qqeJkvlhMoSHC1gXafUh5ZZ//zgKuZ+Xlxa
Erbt3Wb02+9mm4j3GNeH3qTeiyLAbedrGy5VUtqW9rITICQsjxj2bv2gUR+jHSg+bbLTPiIAu8B6
Sqw/Q4Lb+soL5MpD414zKPNZP1VI7bllwpjCo1DHFukbKk2UHJZvDv53BcgMclQwO6Ixc18qc0P9
JQGO+dl8VQhLgADa0oDL2jmU6QGUMA8+zrcAQeXQB65e/P5tiGKa6R3EEKPlbEWxLlIwmrMJh3cv
QU7hUIIenHHWaaDsyEKa0TVl8E3H/9lSkjT7fgLpGwuiL6CAYJnJQYLQqFDm/7PWLUp6ubKXHxZb
08DP/cy0q3+S86uCSH4Ovn+r4AqusHRzCMMxT+YbptZMeQe0E8QkGwPTifsoyxR9JssjmXKPCmD+
JaHTH2kTnSEIglCJ+AvKNERQXfautMNZkjaahjExX012Yb9sY+GNwQeuuLvpy1frrEiV90rDZhKJ
sjcIKzGAPvNM6BwkGh6MpUHplZORaQsjt817QXWfPoutGhuIy2UCXRsH3nGXsyWpyG8Hl9GJ88E9
22rKThNPPY267RFRX9gdZot7/+VEjzA4gqlHQBgUHbSuxUi8GW+Fpkd6VHxi3yGx5cpQMOGM1m+E
TcMtaf+QTrX3Co3yA+RPGwH88rhffpZLdI9NSoDwf+N8oW5XRovdVTCDz8kElx95u7XK2jpU7C1a
g6362W85PWWeHEefPQy2UWB/DiLRXFdYDJHy8YpnC9xcvxUi/cb//kz5nc9fHZRKg0PQYvI6KU/P
oqQyN0XiFFcnobiyG8UQ2p/aSRdSg/7SiGYandpSmhBT41uO7+7j7c+4gh6v/zP6eUR8v43JycEG
C36zxRjIwfOg3qIltEnFFYJDkXDauMMvMmpbBw0+9WFbDesBLNygn+ccQXYXFu1uC+5gaux1yA6p
dXMz2dPpLEi29X9Mv6ldYWzwGqYULPPtpmoT5kfwAsyaO7ZPGPVYMeiU58M91gm7Wry3viU82pJm
4bG08XQZjoIcrR+7lQyynFrqGtfgoUOo5M3ZJCqI6vUlpMW+KvRnpAPSNgfMdARfLuz/X1lmUcKF
mfm0dbrnTm3ZB77oQRjTUw29mwpeHoQdwFz0nlrl+aQTCklzDAbBtB4fHVCG2jMCpfjVVPNlcoww
zDMnlEdnVA/b9xN7LMZ0+6E3vrriliRZ1IkvCRn7sV678zJ6t/392bKn9hLJfuN51Aj25k9qkr0N
rgbQza7ezwGP41FWJFZBVIrgKhWUtMKw9ZlhQuIY3MHKzvcwLInLqdEAYzmw7vwCBkEGwaobyCpN
DW8qRA2qNIu70h2FLm48m/DaQ3Qc7gA+h863ijVU7o6cISqS1ZbFydKKtTPRk/adpm96lYSXFtxf
BZFXFWurTJ86A3Y1ZgfsYrd4kiu64PiZoy7y2WF+MemfzW86rvqUZVtt/OU0n2FZi9DdcWB9AkAS
N1PAdCLa3F0V8eawTa7HOVn1akJ7ndtZEyq3//e4EQuEZ93ktrwLiKmkcN7lXKT6l64LRHERqgsr
Hj4Vxhj6I7bwbY2oRkNZ3vxZDm7u3KD70hn5UFx0DIVJxGs9AspTfWf1GZtn9q72+0+8wPZUYNGX
tlInE0/uO3cZLLmxv6ZUVv1UtpNi+GMWTQt43LtkcrtqxRJ9W80tiZRFoMoEmR04gF/+n7575sn7
ARl0AbCeb3JEKmKTbj/s2I4+oM2zo5yejqkKB/gAL+pu6wqn6h3bJZ+vlcHT+iBBSiH6JjwYuy5M
cwBFbyQRgSuXOdlvqJx0Coziyyt+pwKk5J1kLzyOxUoE1QgUjyf+/3oNkz97cBtSoJJHIG/eYCGz
tbfGR3S5IrdJtUR1LuFFj1PjEWSb2bQO5ruWSxvXrJZLwt78/QaheRBjKTNrLoPX1ofqXexXHlmW
Evm767BI/O3yc3hssOeuHI067Ir5jDnnffht7wSe3N5v0ts1RZ+awAkW69QsDey1RTA29OuVko00
BL666ooB0RQatCLB3jkzWm/26R+PIdQVd/4MSo15nc99onBbs2VwvMas+WzCYpyF5j0sa0TY3Gee
77iDSrk8nvLbwqF/V84Mvtisa+Z08+OHh5bkIHEhOuUGX/8qQc8Kl279FGRGJpI6G3ZRIqJofP9f
zLfqQCCUusA+nD6p6qGLixpX+B3PFlAiNIE842KRMgjb1bojudqn+ojZhbEqYLc2wvkNWWN9XThC
hRgM8qk4cUII9yyEhZryqUNOqbr4/xxLoo/sYS3iKklpDcRAVe+0YO2u4Z0G/25ijwuxT+uBWGG8
JLnp7+6T9682xXyLZGrCBSKvn4c5hMZRuKrakEXBF0J9zTwWYHHn//E085xlJc2xVNCN5XwwkXrl
1GZkw2UDwIi1DurD8WwsDousXtVaPz6/ITaJE/dQy/h7eic5HC/af5+IEu5orMYxT7u6chcwUbfn
VZD+9IPrLTnV7bDQJ7U1FpX4Wro48wgDtRmMl1yePucRKgEV4WX/OO7uUUneuFQRmrON1xmPVzg/
HMbMQUudIZlvcj7UmcQO7b3mO1NEWDrQ3y0W889x5+30HxvwE+jIXnE8lFFH3vrOaFjqoWhjn6lW
XXxPuJm4VPfyrsqNU62SUhMECgM3v4mkAXy+Bcc3eXcI77HUxuIfnw1w92snedz5RHqCFs8UojwV
Yoy/pb3CVMnARza+kxcU/Eg6ys536miMkYrHwZoX3abZwUx5cYheAEnxgWb+N7ahSNEsW21c1AK3
h3WClh4K3PgV//Hty6Y4l7eONMvxEe5uSBR+zinfnzijiiG8yf2dJnrID629DrsizrLp5wmtkEMT
jhzC0GWxAJHBd63ekr1ePQif8Vl1Z8A0eUa5wvdlfAi8kWxp3XWy/PbB5ub2I3zmREf4oK5nhQwO
cXF5tca4NjuUHN0BAOp8S7xasGjgz6NK9D28ACaakKabxF2ttGDBlgjkvoUcSu2fI5PkafnKBdn1
nNLs7oRDownCUpG/xsWCNQbZ8EXZ0moLYyPhUnWDabvPMQWtkK9igaDgPRuCJ5mXLMKQstPOJB3A
Obm3jqwgEoJ0Rzof0M/hv5CIEqBrpT7rvuwbMOpF1kNgVGCGC29Kwy4areBP0HdKMPgBlv+zBFqO
DAVX4D42nsDC5Zw0R4n6MCTzQ91/GnAObCI70qASi75ikGBGfE7xF7YfnbHXYZsbEqGOu3BsjCI6
YmTzoaRA6HIjbYjX1XfqHUZXrCyCsH4+oEMIoNp1qDyJtBdoUIqhhV8iwqMxtzIeNKgktoPvcUcc
I5wyvNLKGLW8j5GoqjEBc86c922bLq5L+B3Vvb7wnJokuHo2wESvW0ksJuli2spCUtb7WmCUXyaF
gx29ANFrtk/Q0vbEZUc9Mp26XqLQRYgMtV4WLPuS49nzFgTbih5w5tt2tM6J/VE7d+55Lo5wk11T
9qR7EglaZ1DnH1Wh7v48LbJUFVdOTcwyLX4HqomNk/Mxk1MEDadVyqORvEhmHZV8qBxnmrrT6FZ6
PWvjWKmJYK432LG9UT6y/AddUupijXnRkZ2nLSmbo7eQOiSjGrc3a8VihZPee57/Fv5NCuqBa8W2
vxJmjjHoA8xnTLKn1KjvwrmHu10sImvC+gl14Q8yTeZ9aeoLWq5xESBACsGd0aYfWMG2XBgmhGUy
R1h5SDbhHbDNVLHk8gh4vMz4N5zFLxmD8Ukyi5ri01T1gq29LrMbW2ZR5toe4IRUGtv/3/0JRkLK
kheN+DfkS6uu/fR1XskYleTjRh/CyUyneML8x3JQVbjxUIP6ruzMOKTu2kl5EvZ/jYznyqymSg1E
ZoCO5meJFcjdatUTK0WywQvkjsTXbeCj2+xImLtwwuIkzr7BZ23kn3NvnmekK438Ct2ow1X3yvcy
gbVJbOkKPmg3kqPgMo6+GvEAS1DTpmGSM+0+vTGh/par5UOuxpAvJlo5CfHcltWC/NIu2xbUz7l4
ncThBjKTuQDseBusIK2tfoHH9Q9jOAonSkH+N9C4dPR4vclk5fzAWR23RqDxjlsqpRX9CVVc0bY7
KIXuD7Orw4Gz8LyRutQAPfPXIL7aABZ5CaHq+o1BReM8OXblVz6DvdoG3nNVpKvmYr6wjAmlhKpr
pUDpGJzWaK+4l/TEPWHid6GvhyYngmt4W1nIOrYHCOOujCweUdwU5K2IUFZhpyhB5JJjv6BVTTKK
7+O2mFA4mvO69g2OmdmPxVMmpicKxwAaz2MxE0CziTOENS8EDoXK++celBP/uHlMF9zgG8RZXomu
e3NobzSYK779J2gYkYRQFUlrrwHk47ZajSbhVpztafx5FwyrMqrs6OuX3+zmCntNGn0ZqK/toTXA
Sc8THK2NT24sbKuYDfsWTRyRuLtKc9c9LTnHy4aUGKxxHCUpgwQLXJEswZSydghGUIoK4x41dQAb
yLWOuDdacf9DfdHF3iuqxUeNJJHbBtYGgV0+mp91AOSmfXZDC6zcMuT0G4euLKCLSS0pdpMAwjQY
ZginK1AkN13NDjXwSkiXKE73YWOnsCyYJ+wmmOnb0CuGjCCvnHbUdksvQQSpvw2y9owl+r2l28Mi
4Il3q/7NJa+Wka7oGpbCUHGwoJaIXbKUSsdHYpW6d9pVazIBW64NPtcMuTdZYdqaK+QgoPv8my18
uYxHPgFHledI+NCztCvRP4DVuYLJHdlwbTiYR92uvkVE5pTcOmZsrR0AQ6By4ozE+tTOfIBu6VFK
H8KVF+SoPzaktWRytJiwLxK1mLH/VgmvQ4XTiEmmQfcOWgAWyKWrIrqHOWEF7s6N/T0qIfULopUj
DTW7k2nm4RzXvp8FBo7Nmp2U+0+4TKZnsuIFrhNhw758XapnpN9rA2YJhn7rJFkaVqAkQ0hVT5QX
s74fwGl1aUo6Ose6/iBf0ejAssvwGRl+zLFJLOKU6DRKp/+asT/gFF4inxxczLnPStXVwDOBj0Gn
5yneNGJM5YnW8cRv6qGoDz978iVs4V4yi7LS7ZMCdopSXuEhk3jzDhqotA5cxfwV475c/T48SXAq
3tCN5EJjvWFrhWlzSKiAWbUfMG4pger7mZ86p+42LCORE5WS4Mek8OhPyqprL5JoBPuaSUUHlGPd
d5QY4V6WvWSVP10NTKj3TPWburDS0SEp9gua4qX5i/VDWDpVj7p7i9hIKd7F4dyRjccuJXbAB2ts
5Y41dhTymXGY2sKtfNk8n5yeh5oYpdd2S5Ymu5/y/yZQrgTkH2Q0aNx/kSmSXH5owOie5EBO1vAG
zKuo1UamfyTebZYO6aJJRFAksoV5nfZIVEccltG+1xU7vbeLzL/6YZLzICMXgtJoeeUUjm0LDQny
x2EIGAx9Oi5T3IEVdpgv8i8BJB8aJnQ9Uw9mJjfTNFbOjkNKE1QAFnqHpWr0867wkXDZq4VHqBYp
NVLylr51/ft5ZUszQdXcRzqvRHwJsqMm6mUbO5H4t7Lyb7EBClYTWMDkzW4h0joRO/teXzmGXAg9
9jg/bPhlBfYmXFhk1P46J0hm2AYt/0zAnuLs/io9Tjn3sM1CiJqBBSZ90y5bEmDdOW5157fqxKVE
OmVIfcQh5tPFR0nscEs/QDzUQ1jRxOxadog53RHdjxcR5RUj+qrmte5W5cEAEw4DuuhSkonxvMp5
tNHZbPihQMatztJ/5gBlhv36f3qfhRtfeo+5+AqRlKTPHBlzXobcr6IZmg5e0eY32yalQGORepCC
vawHBt/jC3JaIIj+HlIW58BbW63QKmRsDyEWDhEZBtR59rWc0qBxF/hP/T+mOdyGW2cC02f6ysum
ePUgulLI6SgLvEjaCRgjHcppLHyXebUPjm1LZRVIHOScYVH4jyJF7rbbIgv5Imu1ZBaabz+dqmhl
WDCiln2ubiGZAVYaMsjECdmiD1RbR9AlwJ+oTniyvzNTPpIzWUQUrsKmiL1uJW3ZwechTgZzZ5+1
hlwzvUU2kP/rzsnXhx07A9OtZ+t8wTWhANQDKxPpJwxwQxAzMT3Jmy90PY75zVmPzq3TTb9rclW+
ByoYMgRY6EcdylhAWhs5HfxcU0b6kXKnL+cQ0IEOdNRg7OC98Ygpvbw5lfHab9WFMeUbdQq0dlHr
Dfvf65bJtmcTkrZZS9hxyyluwPGp7aWhAJJ+cmBO9E/H218kKtGlyjLTOv70sfYRrikrJgTdMjvD
9w3cxg1YxAcAT6fmMTFXV2O+Afebe2QAAkVnqsWdRNSo7ZiktA08oykUyLY1r/XtVKKTnSt5PMRg
kSfnTx0f+o5T0AIKAs/dotpu452gyBg783OQFVrbkYHK7yBq8FzxsfvtNY4mCjSEkoix4gciBm8i
qG6c3j6rYAJ7vuwMXpUWKv4LMsdCMraTxuThSMt24NqcrDKowIuxjcwGGjd3lFlt642QWqdQt9BF
RXAPgbWitLZU5q5/my71/4HvwQOMNRMc9HsC7ZfSA/RtiPuXrxRxWE+hwl4Zt+ft59Jz/xIW7QlV
EV9WGrby7/hSmIZHVovB7sTt+NjFY7nGfSuAu6rJ/u8gsaTieX0Utc0I7gl981zHkY6EUqVYUUlo
/HHhHQrGNMgMXlXMRfJ/7Xbi4FwV7Z0QNiCwZyyrBlffaLdPJuuRqrMfI31ejpnGSCyo0pL+ZN1W
qM8khwkcy9iE0SyZ6SXlp6UZf2ZvAPbWNcY0maBHo1cc0a+5kUnFQ5tITSuBq5IAVFQPOlC2DavN
dmA5X5jicDx4lO4SZVq97L6TNBOyROFL6XcfiQcjHPOaxBNao5bS98LYa93CAOkiQphr1DKIsu4i
acsrbQ8eicYbNM1ENppCA45X6e/OtfQ7Y7NhSv1keTT1wHPnDy99Jqfn4j7Mk6rsSsSZPgkI+cKF
BWK/fzTd1E/A7RRUsHt187oq14qFErIB87HhiQPyNG20px/V0E+BrM46nixo6cyz9BI1RhXQ/MQQ
EuUXZ/4oIU9uCqyhV6GMcBOAKuJqo/HxAiYAxcBYA4+EXztcb30zfp3fjGKosCwQTSKoYRkNC3Ln
3WLiL2igMde008V8tLSvlaqU8uxKVzuacVFvR89YZZHEoZ/crwnVsQJcqjLsKYHM9ese3GOMJRK0
IVLl9HUM7mBtruU/C+SqKrxAtM99Ndm/SB1JXaIQchLcECKNwFutxYij5QKxTt2vZ8P5fWdjqLwf
uGR5nPbtDzT74DJj544F9xuilWPODiqtAOFZ8qNfgfQq6I18bismfio4yYdaVC+aQoGkIgaO+ZYy
tCzpSpFnRTuEwaVHtfhh9lN8TBRDfGjW7xg4b6NRqAMXcIOhcWvlYyPDdqUyK2vfGR436VUP3BPj
1cW2Jal1Lm6wRBgfE7mhRzyY/B4sz95T5/hoKH4QUBxyPqFDg0UK3tKakY8UX7H5V+LDOpCJYjBw
GvkA6DoMmEzez/1BdQp7nBgOLkGNwgIazOTlhmkfp6AYQiJBOkc6bBZYslS00y+0AsI68vXP1KGy
YqEOPf7/e7LXt9KoPFrjcBGOJCWE48NjAZE9xRA7zLDT+6mexjDga8PgGDWvRg4KHgnr/PeysHg7
1EThkIC3EwiJjq9sCpFYS5B3Pg7NUd/YntlY6xDpHUh+i6DL6XlcuUpU2AfXfgzW2yXyWOu+/Pd6
ePSQirHvk/29lQOMI9D7nY5ajaa6u7MjV/n4vjgN8b5W+v7wys8UpwO+UVjU12Z6AjnZ0T74QMsO
OXpttYTqsyK4LPpuAoPFHEX0zAUfl76pgW3m8HIqwHM6tfVL9TmnQD35HDbXp8WD46ZIlIQIm1NT
SaaZnI/cY7eYYzDiBauO5HX12tD85Jb9YMinCow32itmoAEv8NSWqe3aGIB6qp/2hpTWNybOkRte
Stnuqe+4XMxF3VbhDssL8Y4TMkCa7rsd3QMk+5loSdK3INGGhdgc3KC930UX3zIBtnAYtGc12+4x
4HQiTTPQR/6JnQa6TiDp6B3qGtihryyBbTHeEIXtlEBdYoLM485fXYbzN7K8xQYPEFTCiVywBEeO
6hzdCvHZgg14DEzk0Rjgg1a4Ntw5BJp52FgnBmvBqR6YmQActXkk4U8f01q4gmw9Wcy3Nm//2c23
TkWykSVw/EmWTujsax2Gf8KKFPs8DIoZOE4XE+tcoef2K2p9i9bXJlGRO3zZP2PLMzB6ed5c60wb
IWbyQYVmb/s1nw0gcqD0WzM0oQfpQGcWqpqeLCDZolArGbPhGbCXJS4gnMyC49kWCljtGA5kGkP0
KdgMifXI3qBhxRjMIT3VDNlw1JsMw8pCUY1orxU+iDm9yqBURFVpLyTTyD6vU89pAeiHNilfw2Gf
tEq0HqrIUynr3W4xBRE39o4yDeVruqMSUSrxoZDpmJtH3KdRFGdCxamnLQx/KqJ9FUBLyWRVPExw
DqnI/0zWNrLfGik7uQnKZcOpCNc9vLB+nBPf6HeRPK0DkIymaJVrFSNxy5uiC9KbM9SL/OsnNM6V
0jP0+CIfq8oqVUatV4BLQw5IKfhu9nzNw45Jhst7z/tOozxOfbeqR/iVzFk7H9z35hooPOjJ95v3
GMzORn2jr+Vj+UDEeV9HTpkYm0iiRsML+teum8aPEqJkQC+Cj6m2db7n78BgUUZi4Mqkf77otFBe
J+eLx+syPaZTuJu6ievrJjQvg6H+FaxqCD9gQ4epqUlBPmK5VjYSDfhJ3TMRn13Fprq4uOrnek76
nFbR5IfSYZHoBGV6mY9fwA7IV/SqQCRecS061cLNbMMMQIENx2Bs6CPwTYWK2Z/1gOCGVAro8aHJ
LavyOG22mLcf0OPB8P+OlsowEgXiR3l9d/JdEn+hB8iB5Ece5mOM+rH/mDJDjkzna6nLYd8DWlGN
JPPM8hr8CGduyXDENn+VEXDsa9PN0P764uNUgN8wB8OvU26BSW9lnovkAeFyDwKe/37kLR8Y3ODh
dQ+z/XPqYpMkGf6AiC1fqi8KypDdljhD79MuJvlmlBDEP5WrBQQHJb9kuju4NlXGhGL+8zuFNAk5
xA/3f8AagEivmKXk2/zLFp8++amptTdQ1Ht+Ea6f7kxFL5JKnRNuYj3WHUdTBCL2lAesN7/q0i2p
4HL3nAKeeVpfuLBOjaED44N8zxPTMxdxhPa98yq4WqujfPe5ekqpxI8VjcPMsNcNObSw+cJRTSs6
E5b9IEEdsIhkJjFRWihbiU3EJZAfcpO8BruP8oPPEV6163X6OnMq6gl9EbmC1JwcjfAh1MfV3RCY
yjEiuvlhY8yeeDwBkbHigUYgK2eYcVA/6yPgS8FL61wSkP11mc496fyB52X54dsLT9Veq2nPMcHQ
3eJD3KLpoXVfQfEOJkK2kzLINsGRnqypvhgI6uaWIpL820kHBcRdmdUfR7LZ8qn04mWZVBr17e16
qZUYf06W3R2gVCRjxE+ZLeT/fqIUxhAB7OzVIkmbkKnPJa22trkBZLmtxYdVhK+faO1ofk3FRofC
burV6X3LdE2GdZ6XHPlgxav3J6mDaHpU2tGxAVYiKHufts6LjJQIAby75hSl4cAmO/gjjlVWzj+7
Nf8MkojD3cRQicShISY2Yp7qKw5Vd7xE8hAq51coQUsBc67CnK2aC3A7LxuEkc/CEKN8B437QZcE
/tYsSWydurEzpsgp3DU8ZioVboDA1+yHj8nyGxOs7olHcRRZo+YTwKW7MOJs0Xm8QMCRbf5GdJXp
nmaVd6jDFfPgpB9KjTboTG4gCFk+yxpNKzddh7YGuboaDSvPmemT/141HglfXBYtb2lUzhul3rel
MCX6ITAHSu4Iba6z8HhL4H9Rj+lZ4UwNjlFo3qGbjIRfi2UlMzYkHa46xdRjn/l0AntxT3RFVEeo
8k+gUx4VNaMwxPoJag9MCjWjqh3OxAg1zsEdy1h6W41JT70xsAHy5nWP9pyXe7NqVPCbtxiwe3mw
8qpB9lUMM6a6+x/8TdPzQ6r1yPv+IbWl17cbP21LCQYGi7wVuDoaxFy2wFtnbxwWHiXaBN3x0m2+
bIM6is0LFIuAq5l6Qpe3H3Glu1etL1aZZ/I966U9bquCUxPmeAv6YEGe60wGpFMI+R5ANzAK/JKL
c5vR2AgorLbQGL99sRSMyZGsOFvLv4iaZXF/tn7SFD1ZxXRWEQhYo2CZ3DqliDER5Jb8ZWZWp0O3
T7lL1lKg7dmc1ygKMtR2PmJWh0/HibZ3ufem2FwQOsAzt2abJWw5f7gbJRykfI2sE4bq2maoa9iK
uoz165epfVZzZXLqjPzftFL/KuFMtT3NBbFWSboMoKkiiaVtIyryDBsANt6J1MaBwZ7tP/rxjz9Z
/eKYYPpokWjZoFqLeZnwP8XgIsfI6uU1AbhHxiKkVIZEwMjqjyCUufojRRY1qBf4VMBTg0zM/8ZG
Z0rFLejhm7yiI39j++qlVU3Xfi7edU0leOnQqzzY9o0qsv77FstzQH5Uz16jk6mtZMSFav2Lb89W
uvxiTXKDU/4JtmoDB8QVyEgYO4L7AYtl+XNnn7OkRWgegOTTEW5m1t6uol65B2exnMCMZon6n+Js
y/DGustLPSOxw8iurcMN+NWKqgnJcQxhOGuQCp555NCZJnZQeRdltP0HbT7wa48/oho5S3oSiNSm
qCKvnQOT4c4FdPArEbiEIRvJES9wbCNruuTPBZgveFRZsotQuKiZn82Pm3WndX7p7FgC7bg81BMO
ZiJUAfacIFTy09bYRlK3sBDsDVPrENpSyK6KHTuHTIME4sxP4biE3UpjPTRUVq9uNw1LdP/l8GVu
bOFAiMfEgXL8KbVFcQxUjV7BampO3+vSiLk8GtY544PIjYzRjEqTpn5B8Aq1P7mZ995RESaFwcGj
xti6Cf+GTplrbb1oU2I36joqu7qQZUwsgAReIVUzo9p1dokVwW7Qfeo9fkkdZW4l65ox0b1TEvuM
Pyv+Jmwj7FlyLczqy+Nkn6mS6ODuJhc05+3rQMAgYmh6mtq6msvUfiMWA0hF/9dHeDv8Esc9Zw/c
k+WefENDD0eFKdAd+Sf10YDuHX08+T6vsF18h9k3NnxcuBDhmeOn500FCqsPtCimBYYh2SVSBYf1
AW64JXq4pcCxNJeBNYpfRPU783LfyHY4KNzhHwUb60MDwQgORQ3QzlONG+gwMLv7Qh/G98Hf6pJF
8vGCwK16T8psaKOq+Q/LDN1rn/e7XL7IUGGd1TsgQ2Rmk23HFNqeOz9J/TbFAjDXdMdH2c6agbfb
KwX4V0zQ+81QNuH7E5yu5cHCfN+ptQx4OxodRDMu3O5mHm7SSAdJ5yoLeE+Vu+KjYQ+r9UjXvQb/
z0/iDr2Z8JnpzgMPMVQA/lKJkEowBP2ULZgMK+as0XEVE3esWtc83qQCbatgCsyuyS638h5NsszS
TY+5luzCj90EYKWHmbZzgUUrDGUKLZ4oghWBz3arNJ9pZhTsyE9Y/6j4jdcwav6YhzBjsrGbyo4A
q3rMp647KTdajLwNxxbr+CZiUijzsSbBG7MYwykBNIZqkQIP7Th6Eq9z8AkWn02nO82WVWqEGdPM
GQGcqEOX57lyV72jxjMw9jLhZ9G1Dn/i+Q/7vO4VzMuANlbxu9nOhtnQwF0nDCG9emNnVl5SrgEu
iYUUg6RsNTDQeDVSrIk2R/sa+olD+cj2TGaObrSNzIvXfzaR5o++hH661mo8YmzCeTmCZAcqEwqe
F6Cz0spbZ9hp9pjuL9ZEdu6BEGycZ7U/oJwTpTY/vPNywsBTUa8c/euk4SfAW2F5KpejHpYRcl+6
VYUVcb1hr6x/6maOw0Gj5qW7Yf+gckg7yQqYboqCvFIuPnX65bv3I2qSIZU+NMYAFrOp0lyD82Js
b6yyEGNNbmdZFH2mx0nBZgwpdTUQ/iO+Et5hWNjeGZJlS843deHDf9grEhx/tMT54B+ez7XfRxzp
77r/OQMe4+v4+kkZiUlBsY7gHE/WHQC4sKKhf6AfIR09Il2iq82HFTVC8dmIOCtcUC+CultMQzmi
Ntd/kz/wj1IzcQMy+pZhwupMiCRA6fZcklfj8Hw7/pAgBnKOB8U9QUJXjWS9+FUNakKcMJpyRRBg
q/Y1wbX5Huj9xwWGM2uZiziQI2lSR7nFcnz7KgIyt1xBA71f5AaGqyIw3oAT8ht4VS3U3AVsKS5K
c573kKbs028+b32Olj5GBhd072IZDRHwvzhvuFbjukVZiWsGg1d298z3gjnL4Cgfe6vPEC18K6BS
yvTrzgn+V2B/2LjZSwq431UuCuXYxWhHBOrZS1ySu7w6dvi1zrigfzt2z1cjojKXKSHryV3yV8wd
/Kl69+gyAhw+I7VceamFbSz1qLqcoDWZSmVn7r+ITqcnI49iZ3i14yA2N3AQWR7Gu0xx2MeHrW6r
JHgJD/Xv95nJkvRi83QPhjYqz7ay8n9FJirnBMQdWtjq6LAQlTwYQcuVQ8FpcB6WuQv9ACZVV7g3
YKpfiubQxpi1mVgvfGWJtc7mpzvKvyUXfI/y4zKP9UoI53zXc60iIfO4IhVwD2kC7hdN6RNWtO4n
C4TsRv7NC/vjQcm3JqyM1BZshmO4LLBhCJ20jRI9LbtHynb2MLWyf8UXscu6tpIaVY/9+1kd0VKq
RR127z5/8oacGVPHOJ6rwZGksHNaLqwCxU0UktcGhW9k0Q5a3WDbOoKwNMwU+fIXtcGZBexLCuM2
8Bzq2vK8rQhdGrD2Zr46/BuNExpdBkqhaSQyCaHUNC4Eb4MsztD702GoVnf9lbCOZqFjlGsaqKp7
hfbhGD4sovoTz9NuuTvua/qjPVzum9vAM1wXKTI2C6ZUzQepwDWHgz/FLkr9V8RhQfrzWn+KFtxp
8nSdnGMIDppfCFiuXynOxjIMdxAO+On1yhG4UMlGtOP8edmIFZCfsTpg7kO91pq2Iwv7VPAI421C
1u+t9mWIY5emTNpTGi+3HDS8s0m9lJcO/+t5PbjOC5fSJIiv1t4q02vuUEEz4s3Bn529iJjo1Wvb
GgGgucTHI1jz0ZoCpdrd4xXQv586AaRQD4Cyq512so5V5CZk84qnCyMkOd3zFXJ9A5t0ottaSt1T
Ks3lJfYsZhckryiyvFoBm+seizN9tcft2AR5ldbajdVnSOuBliWK1Kxzx1vfueOLeC8siVPAwCOI
HIA68X58QFCAEe5lUL7aP5EAti2I7dj0m6RGVhEsaz9D8VQkppF32Nc9paxZfL4qY45WaZ2jcTvs
w0HV1VdA7AJCXfzAmFqlTJqADvsKKK6lVpRhjncgcrEPWIJTlIcEQBReb2CqhxwiQlF6E7E9q9Dt
4JX22r+DMeK0nsVFEi6+RMsX0921rqAM/jr8fu3az4oQzMcOxWW9w7NTYMUH0REReFp1TldM9xEN
RhFF9dI0P4WTnE0gckm+W1zmQlup31icGjPjyUrdAa7y2IpivhUcw2n5SMgdnbmv359Nbrvxy+1D
pH742hAFzPYZ5UBnxrwsrMK1gaLEmxrd+T4ztwtu0jS6WtHxTKPEAj1p0eqgf1C9CHgQz6GLvLCx
0Wx5AQDRbcjfZfjiZZDLCzs5MEu5Q45JMTozfQBASC0y+KkjTWVgsNrlt4Ij5HTw5v/Q+TiiQgWD
qOKcMP5SwPzenNxFPJUqGNQd6y5dnbL+vrhUy1ENKdHbar7/vTGeKv7ibOsSLI9nW1jCgMQvIcxC
kXdrIPDYwkZc0vUpn5efMARjiCYf4e91HVBNhxwqWgROWIm1okC3Zfh00vGz+2/G42G0OlB+B1It
peWajqHlRL9q3GuM5xKtTMqf3Hd7d3krJzjy9wQIFzA1xUCx9YxaKONxNklZFdlWwLCjDM2i4TtM
blN/WpvfgJRFGDRhpeP4o0oFJY9jQtzeaBJjl2UqSF9FsIhBCCHKY3FQBQOPCA17oxcKweC9qEZ7
k3wIvPvUNcGnAW9rGmN4XPvwvfhyde17cDxp4suUNDPvIfVeUKpdVM5IgyCNGJ13mvF53uKzhzKJ
+Y1eoG3Siqhe++HVFwOQfE81StCcvhvH1eYJsZpStOhCIddazw4r1nljrLvEaZwyyHT4IxwOUYIz
bTDX11oD/tpARu2eI2rC3627EUITnlQnxcdhB4GhTwEZYelBevp4XKDiEfAFl8h+G3+Irpr6DS4z
+VXHUC4dQrH9GU706z6OKeytOZDnuVBz+Fbu3+zIzQt+O2z5b5POPcTfqvaZgtbzEHq1FNxHBhpS
cB121jZqW/+z4wx8O//OM0It1zoRtBFW/JGWoJQvAR6cjDbSu+YqkOMvD/5OcOvR1QUrn9ATdaV0
nEJ2RW877nyL45i+3AdVDdo2F2dZ5zTpjUCdozXlmYuWCWs5FnZ8ZeArT9nisQxh9eg6h4Xcq619
j1Un4GzRo4eDUulQPfNtoEtFM+yRJ/+HTLeNc7TuKZQ9b3c4oEEOqT9BvlDwAKvaH845epoqCEZ2
mmnv1CBndOhpMbzDNoZfIV1pdJ4uQVYG+HG6Qk5DUdsvOCt1pJzqlntKgOblL7N43hFfFs+VcdHw
mxFWWYTymEvKMjvfj2gTYZCOnOL9cKN2H9GegSFIQOxKX7HS9BnRCByeo3ARym5cofhmnSY9b3aK
+Nq/FSCXCA6P4KmJw+Yo4G505ZS1LrRKa9IXfZtHpR3qxCb+7CF/wK+ihFz7SAMtnyD50PvZA2DX
PIWra6Y/XLtrf/ryVKRLDImDG8sWu8gTwqq7Qv96pqlCauORd3ndxa4+L5VBk20cATXI4iVBnM+k
DDf5wX44Lg6VV0AGWRpc0NpNu2XwGqgBmkwC3kVb90uysAkj7MsqRQQ88TBlRn3a1gNTJB9s0gHK
ojmyqpd3kmRVTU0Z+/xylYP7+SCeq6jUPsnLiEzFbbzpm3W2dGkdotR3LkWfMffZs8mbcBB5Et5S
xetblSba9Qh9LDvdqbUxY+bIReYfmP/FqbqerlDELEyL1D10g9tN7XIgUF5cWK2iZRpBONGTUl/b
fCwILCNVZ9ps23e4Y47qeuQAl/qFt5qGFSDswiKmLqob8uxuYSLqUqxH7CmLx3Mc0nUPwBjAB86c
UzOvohDdV8xHlMjqix6rwvC6qyFV2VTrXw4kaKbxh2s0MRf+x2YLNtI0ZfpMXRMwJ+e3xwZqNaH3
EV/AtWOS26YjWOtKv8AXx7bPuPTOCHxomijS47QBGPC1aRTB0XY7/A73FlckIdgP1kXC07XGF0to
9hxMaPXP15SJ+VvqWdd1WSCwIuwyldaweoFOHMUF1wQafyJurxSu/jP4qE+V5DTOTz2lWz2foQ4S
Ru0IDQvLwmE967sGp//aMwKeyGEBPNrELHV4qBCFqUg6e1d/L1MowNgl9F9xFJwfh94cISp1ySOl
7pQm5haIRoFXZioc3ah54xyTcBfNCObihRxG4yXJV3HEmNZVnxWTbyb5R/SeewEAQ8N/Q30wNhEb
6J2OmFxwZ+aDaDIsk5DKTzRFvblgOm9/5EyvOYRlVrjrORT0AsStGiI2dIuuJZIkIYbecM0TQSej
h08zQe/93QSVz6YxSXkIKedLBVeRBxqgo6yL+FGVzvP3etRKMHQQ6R8ce6d8ZOgSKDpeNDUmVHjL
W/vcOfUSVQqNK5kFXqsBv+f1MfmyIOUA4T8b/2tyzupgynWDBADZ7ZMrbSjgv6UdCpi/l86uxJWh
tQnjNcK0bZIO71JTiEoGSleFrvq5JpovwYUfVydP/G+z/GsMHEwPMnp47GCQ908F+vREn2EwGsih
aBU5A8q3GJBob0khhSfPeDRe4W1FKOJ+uRkErju69FR4kK2tTahofOgCMiWCBd1p9oKNuf4++9Dd
S5u/aXFZXKrx4zgf6BoP/lP7qSBuOYhhOEZLPBWBu4mf0pul4B51IGfS8nOWsG6wJ/6/Mp5OmIIr
OJHD2BK2eOtFCAxQbNVJyqkUNuqDDc5gwDNpsy/8ubrdRjGJjCt/ptqf/IaFZrTLAEBqLPluiDgw
BDUzvsvJ1kibJzwG1x2siYtCZrIYIxSKimKSh+mBjH/+xD8Xm2HVk4dqQZOBADFJmM7odyCsiNz9
FM6oJ0+GSw9MP5abeZ5KB+yBuB8NTx7v0gW4a3DS8xybiv6aEVxydZgyAVXG9psdU5i/653vPX7Q
fiPoPn6MzVTCC13BoYgB1NxMqOI94Ox1NY23pM2dC5j+Cc5735YulEiSM9k13asKV834YJBp5ZMj
hhObfe9SlWOTv9I0hFYJMjSFYQdZyz6qlyA/Q+q2e2Aund7ohosAkWE+fmOOgYVvHXUc+rDLJTvh
kAy09VuLbZ/ROBG7byOdsx2RiJ0lyLRPLeqKA1sZT4YoPySCd3a6OaMP2x9E7557EY8coqyGEbiG
B7N4hzwUUPDYenuTVHqnPW7tW1ycUKZya+eOL1tZCpmd84RYSpKC4zeFq9hZ7dxxWx2nLzoVP0+S
jcLDOfYxQbwe52W1AOpYb9ULIlgWx6lmkyxdualZiRSXp11gTnm8hk/NVOolmi4ifPY1xEhSES2s
YOeXs4UclWhp8LCf/CngmP894xk6ht9mGTULtLeM685pmz8tco/FyvJowKQ43avhpg5rNjLX3N/9
Vp3u7yh5c+ot8uDHEWfaAcLz/Cj7nWiBU8TM/OkyoK3sbxKCxgfi70bPuBlhmA2pW8muckktn9OB
GwPNv6G4euPTgIzUN5pm+gFrpcH4kZphEzJqXsuxE/MTodEH01IRuEyOOecUYx0qyo3CVRdOa23/
VrXU03q1RHnXdJHrJOAEZOKgI11AXBC7JyBH8SettVLb+CwO5oHq5UCnblun+5FxSXqX0+KYzDHe
kJNlzuFW8ZHppEaZRO4yrOucFkEAuVVRxc8RbzRaMMPS2oPANI4kPFiPfelNb/N4/kICqzvtromA
QWeyCL2P/JxO+kh7GY2LJXBVx/mXutOvOCG4wZXQV/b3pwiSS/173PFdARyfSGdXGOc/5Nox1vf9
9mA6mrcaAZHRFHKdsuVcovAcDr+3iTLl8N7g7Hh6ejWHI5qnomMzsY5UDJpmtlWMZ1dzydXEEN64
zguG4D9RhderxUE/N+VqL7eO3to9iSEaTjkUHI95yarDsjc6MSkv1csWoiJnwUpRJUdhnlQpSkDm
sFZFbZuFr2G3zQpfNldo+JzUZ3NjArtPWPNGsaPls7S/5MpcEI6R+jTf9x8qY3X4t5h5Yjgra5cU
ZMORUXG6gZq6rOiWQ0Wt/PJ+AugeLnv9PYf10gZ+m6xjWCvTKLijRRVbbcsuBjMO7fUfUXsgjKGm
1TY+fZXunN1Co//ud8s0yH+G8Us2wqdbCQyS3j6jfxH9Dyn4HKHS84F+v1kBTVA0fL9U8PQa7u6Z
0kXjQfZp3ymHmBA4dq/HSj8K+jG4nLSxZz9k9+gFJlrSFetY95brq+vGup34TuL+SctvOQPmIRVA
Cn4vkLRV4olXXF77xyNyAiibhvS8o8SskvCQBwGtEFxDSl8rHMpm4telR+Cy8s7QB4zMPt0NwLn8
OccPuKjVk01QZxI7yX0J/Q3LoPBN7FG/K+iW0S1N0Le7bTAQXgVr1qrBvE6CDB6G+kH6K56wa2gp
y4RHwDT0jW32lIA3nmkDnGEIQ4b4MRC0tb9ABY3FFp0/sSoCxBJSkuqnh8buVC1T1Q0p27j0Q1Wu
YAa3TU1SsgxdA0hovY2LQdVvxLWqXUcJrX0ufVdp3lgk842dfIeYGhpM5OyoVACf5PBhrCkQeZR7
xDQ779e5e58QXdA3WoklU2NuM8alZNIby9EspgKkgRAbHSmlNYEsreUpWsVPJAqX3WKLW5lrgITB
s5BIkQBfjVT7TZM8gi34vMs4xxXxU4lzGMoqztvK5smVCNWA0W6lu9Sb7sLGMRdNfdRhFX8ketmS
yCv7ISpONcLts5zpx2y7UOyiJ/MkGEhZZoevsOapcGnzTNWinv8Md4QvhlRxidZxp+laaArgrY3J
H0RbIdUgjzWS2n/gIe80U+b8zQGT5Dzn4i2uAOnzzMn26WzVWalTgVh3Isc7H6RUSXzT+2dbjF+B
68u+mYX1MYRHJq6YmqENFSK+vsamjDm9Wjg/cnEL/BtTxM367TDyIlNhdNc+2ZnR9E7XYhvNhhhB
+n2yZTpE+DjJTdbztJZdaSw5TLL2UWbiqr96TtRq7rqD4JDJJByWYwMAbO3l/HuUs2tU99xsiWtN
ll5mSWfIi5OTiwVW2uh/caK4fodkRnYrbV6vrthk3UuJwE+MlJp5p0gsQP916fxOuGqQEULn59dX
0l6cf0+sdElTIk6KxLROAgdA1W+u61nEkzpjeNJ9dK8nKg2N8q2E5FJyi0GspD4uc2xxISMhzz7i
HPawjuFIAfi6VTIRDRUVH8/dLhKYWCiolCtZlC9bcNKJFfeUqXDNrDWHvf9vg33qCSjGg6fmDgSr
BJLOjJ/WfCM2xhATsoaqRzbD1ydk8duR2uCCEp3fAWrwOvdiCvVpcqe5Y/JKgdBhaPP8Qg/lbYJm
zqLSEO4FSVgyPhkpdfJe7jCT8HJLOtGTx4BTCjxJdbQFMbntrwYeItDLqAvL1I+BmAKRzB9YN4o1
TN4kcLL2bVaV6wgLOkWVBr77Y7GsS23itY+tOBmy3fTNG+Bk/BlHbMc4OdwPObZFRq0DxWn+id5v
tvaJtT2Pka20UEkbXqTbApjL16lZNUR4AZXKki+vwUvJkXb2Q0xoilmhnbkBSoGffErnmrANXr9c
r85c31CXir3dWYDUbbknNKjvuA6q9KyEU1tLCiP5dJWhaOgkGYDTTWXCbdMwTrzZAS8r2z1svu7x
Bu26K8s1RjvWRQ39KH52bZ+pVB+jQzfXwKxNHbwQQA11betY9nb+IYpC6hqUObhLNqnRFVeSjUVv
Tv+tkxkMmKExErruLr8GXMKL1JdnPvE2tiKWtMhSY3C7SZPp8qAnmdXoOx7y6M1bcXcvNNcGWMvx
IZRirk5d8lCk25H+FlWLLQs3mpq9hMnfdSTEKkHG2VZWF6MWsqbnq7h+e0A9HLVZKxKoiU+7JHXr
t5XV/cbW2svMwMYy6gEkiSNJGTUnSP/NbrtzwPgm4glSgQzqtQEsgxBiCR3GCTwy9aeTmgtVRuKd
zAc+2D98sabKTkl77VWJoiTvema/0o4VcDus8LD54pyyuOzc/q/uYH0aDVyeBheYzO2ASC/yjA9B
ocAWdWm94xhx5x7ANhpdeCFgKMPs4Sn9+s0sCPFcldVrAk3+CDCK9oKtkhdpOpSb8gQXiQLmFFCP
AQ4q83dVo7MMa5M2/e+uX5gGlZA+ikuVREOFB2TLlP1ieJmbjXKkO0qb9Rq2IoaaDG3079D1wXm2
8xQj/AMNTHAwLz6T2UPIuGoCH9FIpTtlNyXBFZntWsuDM0WuFbsGBAmi0mFoBGzdZCjmSlDD4LJG
XCbXjnEaSjhjqnoJVV9Fg3fqhe3eSvPiiTFRF5m+H83nh00xIcXAUL96//bhHn9ToMYAMMUcprMH
Fb48nWZpMJXyh1n0ba/Ls1l/rByPx22P5TMK71h5Ni439mwpCmKrMvHhOuHq3httt7svwVWnSOUD
OA7PVNGRv1No/RPlW3n9Qb3AwnmgW77C+we5XrG4MBrtdXhBKiSCyBdOd6wc4H/h3L9yTcE0gSGa
WEge/E6ttbmwxeJKBpzKdH5rh7fNzSkcto/9QndlRTbAIlQHGCzjJM+TFQ7h3DymMAJplzN1HUvi
UkKF142nFDGv8CNwgFF/Xzhxat8ppyi4PFd2FQgmaMrqnPZu00rM0kdK0E5LY++CB1m5Xp4z3D+X
Ke7aaoV0IzRV70aTXBgnNryaS3XR0fO5F3P/jk/0GCrmsL//H4ExVJKqe98UvoDisi/lOZBODy2g
EM4xNXPwN+aD7gw0PMHlPTXC1M/i18LrKgeDqAB7ReqmvVZaBj8TMWhXusHAZuTLSx7J0m0daJgZ
tcpq0JCLMlzhgX0Q5uB4nsGWLsY7me2Y5W9c97IAGxPfvXBWf+6TaUmWeKVYP5pD5USoj43if2jm
rSCSmNzZT5XSK4SwsqDN8X8zWGLKagDbxCEg5B8M3NfPqBoY8XjKSWG8B6T41/pPeTSmlgU6MUIw
dAl39X2OCV0dh6uerRV33WaMFytyIRCOr2YWKEk3E9Jm6jkx/XPivYov2wje3msvlnAjrXSkGrpK
twLzQkVa/aqh1W89/AQJe7WcpRS4R32YQejRGddf+u6KDK4aIAsdvzFKLTbOImVoXnRJs1KxoNMk
lK5EPfNlLjs7P6rJeD66TjovCCoL9POUt0ZiwxyBwl469hoM7GocltjC7XVd/ymmqIdv9vC0XonK
mrDWqopJxOLd7JRq35LFIKCE7uPJmQiQNEOWq1FPFjilDoy7GjddfQaCX5YB/u4hyXdtwXF5Va6P
fTXtfh+rZ9cWvSIpIedGcMQ7XDO9kxmlVYVumYkn/PJpR6ocedQ0JddMa2D4BqHe3PpHTORY7gJt
z4sRqGrOv+mGMfiP1lyoIBq/QKhEVtwTeTVW5pIL0jHZTfhXgOQAM1FyjegPNnQX4QDJAD4u1c/3
4Ks0xkdShK83Dk5kDpWsz+m7r67ba7Sz5UZVNtlSkAMHW5uqSy6fIy8gzM1whSoIMjJEK/v+86RI
vGiqSwC+Nc8QWyjCrAajg7zjWjIFLCpDVgQU/W8MqFXhwSoyvi+XP3l0vhDOLFP2Sj/gzoVftOs7
TM4DwjJ0G/MXA503gVHEXeO9BWy129ouEF7HXweOZTAvOtPYtQaYN/e6N8yRrFmrPUyX9EYapgpe
6z1r2JPDF4XOyNBHHOvE8R6ud1c+i27WNWBC7H4oFtIMJNwV7uv6O6EFaWVXm0vHi73G/6gccdFD
mNfRQagBZsxsmMCINahrjeoLH5eYi3oyqQsrtHXA4jxs5a6FZJ9jrfe730o1lMuC+fU2gdHyizSn
P08+BQX0rj++Fpz6NSL3Ykql7GjczwJFtQX4KfVuqnb04hNaqJGNy+LSH8NpxNsPJcA+ClulMamR
Sqkq/3e73c2i1oio8yHl4h4fJDmMlHO9z009uH/6AQ8ttzcKdmPcqz6XSLpndvsqZBkMr3RYi837
klVBl4Z+79S3h+I3xf1wRne6c9NVkVYUwnb+on8pcsZlbvPBo+RydLm6aRUe31JDS7SCLSMvKBHj
kyEw6G4l77Ez/VNx5xwPtk0R3cNeV/XhQIW1rLJcZgWhksx/+ohEJk3WEIcFNwZ025nbJ+Hvacgf
QBpXgtvW3z4mBUZSaHCFjvTUarMcZwQjblIUSrewDsWWgAb64PPm3JyhCPhWBpyaugsHXCjvZaj/
KXNDydXd8M+2s3E+3usRX2Z0ctVAgfg858rIKgwC4OmK/zKbjrajsz9X4KjT+0P8zOZWVY6q6iBN
IUmwYKTHAku+5n0xDg2Y786hLZpseWdsqZDazYxKOKcjQteVvdSEgORzoLNk2k2Hhl4Qkd5jStU1
/Xk71bCs6B60lT0xGcr/LvtOZWngGY8LQxb4JOKrgMMcggYejVvlFxGZVYSZB8fsrCH4KWg3o6qI
MvOxNPKNy3xJcGZjWwRD0iDDvmk1y07vAfoICk90bE4ABaA7jw2Xtv7ApeM6Vkpg7AMS5PglCV+y
tDh/MLFw9UDZx8SN7ZaotW9LgbgAC7h3JxHYSdE4MFZNC9bRYk/rquVYM0aWwggEVix3MoFgKKFB
dY67vYhBn6qrLYtOsVnEoMG7UE1d6hYPKt2Dgf3luhBmH3GgTa19GmzLPhslywgJKhAhiuu3o+hP
BX8M9ZLINXd9WTzQ3mw5FxPa0B7Ct4Ium/ZtlfoVqjdNnIrb31R/H0UD9W8wo3XPTpftEzDQC0Is
yl56zwwEfd5bzDTjQI0/1XmFZ2+ExwSYt+8H5T4mH4jmFw64EEyCahAM0aSAfhrZr98PPoJo0c5e
qqyJ4yKVf7px9OvMw476sdGb1d8jTGg2UZrGgPt6O7enTl4cHpQKrkpsfri3hR8wIjIkiOSCij+R
YCQBjZX2zFDXdKXbvrU7TkNgWzjRxr0S/lj9wffabsvQoILa5vEOZtJGRODlms0p6a2JXIhJMmNX
XH4XFoPrln7O6e5Ib4QdsVuLo7iZYH7Yf2IYnBk1tI30FJwTmirijzchBrLCwya9HRdJjlTiAeVk
7uRFxMRzpgIeD5j34ZTN1TVWUMWkDIfV66OorWBd4Jb+9dEKxeWciG6GHoDL2sujzFPi5VUt0Obt
AWxbq9mBcwODnImfUmWMU3khYietiEG7XLzBAVQBM9msf8IFZ+P8jr3rWyjWKdf75d2qpxexGSHM
nRDX+Df7xKAY2F7dhEwduVz+0M67/Sa5D+QKi0bWc2JHKwY36u96xUwrVm+cwUasiO0x/5bd2Qdb
gOzjZ2cFAbIyqDjH3hYH/KWMU62wvitmb8UzUn7XjuCBKTmsHlfJAfoHLtc+obrIz7SkIG/xDGaX
tQ5jioeVLGO/57k5Gkun53CgMGR9TVo5qsNxvsrOeBLJ7QhF1NQtjzsoEq2yGXjIo8TRgOvCeLT8
pRI2ZMzdFgxdiGCIPnDrRjabXSlv5U60jEp8sJ+zlmYQDuUwqyL86qmDL8nuGramu3R1s1dZsOQg
niTgAI1Y3j5Quen4uWoTvjVvbRQ+bMFRUpJEb8s1FvP64nlogGFvje7jzaHUxaYOZJtltFL93gTL
rPYy2JiHnLWk5KN0Ps3rcO2OwL2XNvXw6aYpb6xJlbDldkSwJZcC/7tsPvSiwH3z0+NZLHD/jVw8
BTvtgz/8rpyyujyDOJAn9sI8LBm66uRgM6GdYQZBwyP7aZ/SPObH9hknBS2Xs89zlEXET2RbolEM
aASSH7hD1npDQUkGdTMNnMRQ6qUxmN2hmdTaeJPCJ/3cQhzNWb9Vw97/WBVgYOgNxklwg0sW0Mt5
A83EvIBkB8Wy8CeoneuPEbFcki0cv22/mXtzdZKeJldoRuKUDJncPeelO61SrS53MeMwd/8Nfa66
bjR4jO3NBFCnI61lE3qz1KaRfuXf/JK4WW0sQ5XZ1XYAGh/HNSHqMuc+lRnJRqaH/TMHpK3QRrVJ
/dZ/yWL2u2Rb4aVE5WSXsd8qwWYj30d+1C/giw4dlcHXeb1aaFXKJmXEaWt5kVHMu5lZ5C5XhH+q
qV376qQPTXoaa/BBUo0IJKiKNme9VSVS9UVhkNZVSTcQXP9YiOHC+a6+mhi5A726aWhSYp77oXcu
To90T1806Nubq+fgyGyL0N6XiNVMHLkFdHiOYE8e4nEXSsO/2r13U2qvlWVAhzl5C/JhCOo/k7n5
j8RIYcK13zTT7G7RMxss1P2Z7JU0HrmrOowadT5aXarYzCGlKS2SF5BSxw5MHVutOUquMwgtGJIe
qeekmsPk4kh+L/QdDq+DAjteQeipdNo6MRRshStc3oyanDJf435vzrTzELz45H00kcDi622XN4mt
peeqbw3iJHfBaeJsnj0AhjdoHtq1W9lN3KTddK/fnmnI18/7sjzYo4MrsD1H9dXgq4dsNBVDAUgW
HGEfkglu4hd8OdO4haRQijQRFoJspqXawhIKyrYmALSHULkvx59MJdXc65DbXdCxik/Pr0mbdxTO
kp7Ex33DMi89jIWZXP/CDqdvpnW3/XNFPu8oo8T0lRICXLtym/cYy/oavQzgCAmVBTkpPKtaEy4z
+nXif0EopPDRn5HkaH5PEt7YTNFKBoiHMJneehPgddZuNdLbQ1sPEx8aGP4p9P189auPksNAsBaR
n5qm5FN3D+rrmLM16S7Cx0ojDl2dEBUl6LFdc+defwGTXHd1ss3Vj0KpR9633rwoNvv3I3rx3tQe
ViPGpw2ZMeAyUEBhl8oHS+J+MORzq+GKn7w3ogMP2nkqSdl3j45EG0PFspqZlx6gfDTII+aFWlwI
2kEYMqDYoehDP+FHl1w8PA/JfHTqyuduXZdl4jFnRjmdGk4wU6IcRE8CDafFE0yEQ9IAcfIGnsxb
YWJcBmcjK85wNpUyLk3GSk32pdlRVKShnKhBV5DvcG5QeMtd+1ArTQ+9D45P5l275lIPkkWNDBiB
urqAuURD2dfCTyZh8YwvWBDpwUm8VRYLrAJDbQk5G0KFxx7qNcPkNo2pYPjEgBfBGZYIstXQcnbk
JEM/I9Y2kLNaCZU9XHTCuY3PumChGKHlQYMJGHaT4mmWFj9IWnSCFkAdSYDUnCQMZzY5TQvoq0q7
wJQlXczQl1LNpdHYwbIBwLN/gKmdzfpi7pqQTZFVcjtsswFhQINLa44YPAkBaVHehV5tpX8hra6N
DobdbXRuz8Ha6XpiVrH89ucpgUPTisY3Bv/h3vv93J2m3RQ5W9Khxz3UefGAY0mJMr7DQXUGlnmY
KYLcxRaYpOS7czz7/jlt4JCuMYZBIOI1Mbvly/ZchLPoKegqBAozunE4rlDSn0d0GAsU7FWczmNI
SbD7/oAGP+zvoIVY0eNUu91y8aFHPuPcq8By3s8PursjL2rkk+XYpDf43ad4WDZkxICryHx5PXdm
eKNNhMe3lWVJtAJthGMydQtanKImF9VhJxSkQkkW0PG+c+hlEkmpmVMv/TL1xJqFYU2dl0uIZGDn
rzVXzcIN1ztZB662FIIDgsIZg2lW+k6kwULanVPUVI8p7EHN9hTQoseXeX7kEVWIddivEdNFHnN0
AZ9MZi2uDyYqGYZ/0pJxi0GegrIHvWdMT2EwYmMwWpdmTRUaLOFceXK8K6oDEQo9OfH1l06Tuy02
lYOSjcz+abGKZEizoTKwTkedZEB5bKMnSSkCeGEY/du6LVKMl4XTVIyCnd51TyKNgEHW1MlRgGHZ
Fq078l4+PVF+QQOaThhl/YLzmn7qRv4q6Xv0sczDa8Agg3jHvG8ULnL/CFUtnMFaGiD+YUIHeL3q
jociTbJqedMRzfKxtMcuzq4KmVn5rDH6+p6FwSZPDwEnFLelZI/Xk5yq221DHSm2F4BRJj9D6vxr
hiZVOmdFcCwSHKwCDniDGj8Uh5SJPkhK1cyGXG34RjI9INzQl7Pd+rfOqTJngJZ4X1rU0sdHZMku
Td2LQeViSQGSC6oIn6s1TCJCKZXiv2xF7Qgcl9ZxCVGz9jm+BfPb6q5K+QHni40BSd14KNEspoqE
kzY1bEIcIFq42I41JVOB1v4s9jmtz3bSWDuEULlnRrOU8WJUQjesO6rGSi7xOoKhDAXxxSXFnQsE
21pSRMEu5Qh97FW9GUwmHAMCAwfDVrM+U5oJiQksrsFFeethZGjs1oIswOrpq/tIrUlM751grS17
+E8BgnsEZ874o9MAzu37SP0ZjRwMhrPQE6/IObjqg7kvHg7aQVYacTxFFkYCmbCMxHllyaj/UuTX
M4f2g7YxB2DUMOQe8Skl9FQW7Fx2o4VSK3NJJpYnJ85SOdXBA1uvDdFqGSZAkxGjczl5uHV6zFnX
a5mxnQuFOMuLiOqdXqlARc7zGWmoqLiZudzFKhqorr9KIrTGqEquNj8/xKHY2Jm9gcQPumI04Z03
Xpe9ph7zCHfEIjyYgikhJ02owtO2SVXYbF22fPKSVe0nCNqu36VAyDIUUUxzhI3pvAdQrGvUD1FB
OZuQX6lhDjfgtUHDZmdLpn2F6yHwT3/TxFSoV2EsmBntVB27YFD9gIe/5QcRR4jBx5OMw1rBMg1H
vgmMpwn6IKSZZaGK88dBi8eoPJMKT8KOTBIb4stcxTWYVlG1CezRFONwgNj6WYsJ5uEPn05X3vXc
tzMpVm7VrLw5E5a4BgPIzKkwD3UTp6WGxXESAzFB9VKHM9YJVi1FnUztm5pqwufX2ohkZUlmPcPW
HrZ3cdoN9rS9k68m1m/w7oAjVOeiw5J0dEjXQW123EqxI6Bpz+a9x6bBcz76T9iZ4B0Ffe+9dzgW
T6vPKG9bRnMGqce8Jjp/R96s+Kr0NRImMhJPhV/bekuX2wPtw7iqE5t3dkyyu7ud8FXWTunZglr5
HePET8KuhgWpNE/BySm7ftKQBrPcUpRTz/KH4+76ht+6XaUolPnR0/UpcTXDtgjEb9Gh1pfbAocm
Vbu/20X9oLYPMPStLTcGSttOL2PkH7YejEBZa7JxfIby49KOQI0YiaNvARoQppFz+kQGXH7wvaI2
1Mtblrd3+Y7fuzWSRPQOR9nxZ/9rlgBUJJAlQxPL6JfdREiaPS7NAzmuHh3ziRQF23URHLEQ6k6K
nbTFnkT6rgpPCXMU9MwADzhrpENNdi9dLiUt3rnidUMqK0k2qPdj+nZXcSarvQz8xFLW6tPEbJFe
gMWMJINcaUKSNusqCamUykwjVlBv5MDmKP5FWX8VDuNhWTpmpSG7vKLLklghzRSW9xhQpTHQjIbZ
NhnT8wdh1vz0WP4yoljb7mz+AW8GnjDHyYJxmmIR4sbg51aPS58crtHRXd3Va+WoDte4vlA03CLk
ee2nnzoJ9UVlsFBb+H24p3viPbFh+60a3nlNZGRZz8Yl0rEsVLdoMpJ8IIaeR7nbZhQ872d9kty+
XI3o0LP4vlcr7qcmFNt1mhW7zzTtxAEv1TM9Qhq2mROVYZ2sNGPm9+AsZwRkEKaNskXuhA36E/TQ
18JDDnqhFh4dkU4ivvOWQPXWmVdgTVjbofk6+Vdg0206NjWVldelwx58csjT/P5knVN8cohiO3TX
FKGsOUBAQLfc35jsaFC405dtagUZ/LjpdUgHFYwjnl2JnQlqPYW1hKCS3Ouh8+vRjevE1Cv7WNxy
HUxS5kRX1d/IbAQnz9ticTLhgCxxFPPGsbbwecVJYOip5FNE7oQ+oxmCrJK6x/4WagslUToLs5o/
KtXC2VEIsRseh1nqaeBDi/e1NtniDdokZ5W8wkx1WH57hJXOCYqe0ZNNkCjNVRUX6Ksjg2F2Hool
AocnGWAiQO/YMR5BHC0q2R14O/JWqSt63UnExl9Y1Sk5MnBm8k11IYZMk3Ct5V5Vqi+e23imQrPp
jqDclx++bwjAf5GUCldHETQmFqW/kfDcs0DpJLkFRrWFgmpgtUGIrJex9FW34BedbucViFB+PDwx
zbwcE7/Jf94KDp29eUEoO0/Au/8MGS1RDdF2MtDK74k40/wrjm4mlJDtWMgzglN/WLiXgozdqXWF
DqsWsUuBYNr0LALh1y4KuvgZ9Gj4j5pEsoCRT/WQ+Dt0hB+U0L1KkjHdut+7Lui+SICMO3ou8XJJ
tIKK7b/z9eJxhc7WfhIkAu8OT1LRQJQmyMymrmdwhCnI/oftwUYcdj5nNDRBOZTOuDKCSyNs3K0q
Pg3+HGyBofUgNSufH45gE9K3u3Gy8XMo0P8PbNYX5MyHeXGgeOf3+cIymjPWfRI4zq3jD29o6194
VxiuegppgKfdO4qMPmd2+BQfxcCC49buzR9Xys9PjUD/WWASAT4G75/jzFhkFWPLwR+OiKpZ6n7R
xwfU2AeTlV8byGUiaQ1mWQTwApp1J7YJqPUpr3V6CEFHQuO3Wp0bSYBXpbddbLwb3tCdMeuH8dDW
A84hCVBM+7koy981ah3fHT0geFJh4p0zKsNszPGibpp2BEiDvmDn42kfCxTok3m2X3k4aWV4Wjxn
03nsDnpMFOjoPZiMXZKXquXlVgOrjzrdjonO99SxWF8qywCCseAUzR/CB6fdFPor7AmXPIgvgHg9
2pBN2VBraGdSwpkenRPKbp+hUPcn0BOWh7QDhjUJj70u3O3v8FO4+h0G9OkYi67DqI4g7hxxvAHh
ol0/dHgoT7LAyv8aM866N3U3FLXDU8l+Db/ccGBXuezi/9LFoX+fsqtoMlUFwo6oLbb5XG6qszN2
XTiwrutQwUJbFj3beEbVyHrAFu94W5KHCmhq8Sq4al4TsCuyHHJWF4HIrrPnkl12Con4FDb84JkY
HOkpAo2eCsaOHjwyiOVvja2DxHV31E2IQalh+y3tP4mq4rHzfH2/xVhE4xiq/l+KJLvYMSRQVO6N
VICrTp82u3MyqQk3c7tMD/o+QaxLovLfXujaGwGjHFq8ZZzN2a468a7dNiThdb6f1Uy8975hNQEI
ll3twqkoFUnL5r3+4lj8qaTjoHZUlRBQhuPcb4GbS31ChC0c6dmnZSms/GeC+ZfyNGXn6KLgwXee
tSj+XSrtzJvNWW/LMgPgn3sPJkEOrOBn0IrX6kEpg7L1LSJmcLTYVV5S/eN/1fEt83V1ofkqa5uX
wLq8rd7N6VE1AKDO8xMTiMAEdoBfX3NkGKGW5ovc+yG9XcBd4+QbiWVXsLRwD4+CQ8Qdx9ir6zZP
hdaNWrRU0IA8WSyO079jnrtrSp2vHoTUugzLfaPz+1vFbHBAOkJcz5hot38hjRsSRz/vvGCJ39MI
50GbwdrCdZbjSIuxKWlZn30XFzrMJP0NZd+UnfYcTaWtV7ir0nXx1ZRRKkIjh7HuWc6GEUtc90g6
YCsrocVa4WARGD5uxmGQqTeM7rX8q/1C2LtQqhPs4BcmO0fDQlJuIEVitSjx1qC3G/vI5KtiA8ZK
Fl8wDusDvhpZQC/m7cputZnpIvON755QxzCCJzn9blTWPvgBGkhgS8dFNhbFej5Dk7Zd4E08XBz6
edZ823yKfaXUSOeUJ1xe6cGJUDQUuUtJgBWfFZUYBkt021lR/FG1Jyq2fTMIVXd51hQTr+CuNzHN
U2dom6jsoVlYMvCt8L/IeqvLgZ73bdbpWFUtZq0TuEX58AGAVPy3Tssp5TwmXviGex02YT2+p9t5
/RpRYykwhyZ4MHEmju2Y0YOFWgVGmLoC5StLbDNp4CA8tV3/QBAIjM55KGu6cjhUY18MHEYtAVLI
DHyF0FYotsIBzGCUTR9C9VepX4x9CaHk/cU0A//tRk0+HIeBeN4PWzFf4FlVcIxPTNv3gqmnr+s7
OkeO7xmTcdczRvm4kwlanUr6/1Yah2VoKLiklu5C0tPR0788sHUXitfxiUT4zSaHqcc1vUfEkMuE
cYDnp0nGQ6OF3cdOpLea1WLSDt6KcJpsJ/vrzY3+mYetZnG/1UjjkSifvD+Dc4pyq0vTzDiovLgy
G3nxlOVDQ9x0XAoZItbt8ujpOvuv9XzeshjHfkzWUKtiMUPilo7uTIwVKQH+bbBWk5REgTpzzTP8
v+bBh+bDON+PIPWYvVPOZIscaQfVN8heIDiuQKxysJ0vRkP5SQK48+6bCKTZU1MS6D5y48OTLwPF
KDi7L/zA4uQWYk4F8z52Nald3pMNwnQnSWccSLWUffRgwCDjnIe3J3K6P8klSQ9tsJT/HWHKLan0
n96s4AOO9jVzKGXkFcfvPP1GU3YnVC2Jh7WWQhozsSbklJDQi5vh1cqYYNZcSR1U6gOk5UbLHwoW
pDniAgrKpaHL1kOZy3AscoNEnIbt/yvWYqKqCj8DEBSDfHrTlw1cf19pg/UKOXjW8Fz6EzdQixFO
y93qLnIRUQGifXg8gARQuE5mkg0NCvIb5Eeaupye0mzolF2hrPj6uCR27Bt1NqFvQoOSp53rIx2u
6zQenq0Q/KUccIXJXY0YoW/pet9ZwYvMbrNCpYb5FmgM+PBQPMjNHg4qGRvTtFr8itexL6STUKKa
HQK0zzdzqn8iY2gzIOYWBMjzyhAiobWyne3Y1F6T4/VN0ZIyC2X5xh8uX8oNgc1wEMx8VsGEO3OF
0GBqkZr4pGNkiu+YORdzp7U+pQVcmz+I3IO+dB9lKpthAfPQyLx8/ILjn1IByberQZnF/BRrsMaA
8fcDzBj4GehQEdzxEXoj+qRTW/S9qHRrOPsFDeKLDkzvgtDvBnc2Ir58Zod4IedNV4xejp2rItAW
PXP4T5SqvuvlpGzGd4f4tRmy4mCS/1a6B67Z3++VRH7PUpF91anS5fkRlTK7xzBWavS1+uGG77f3
cmrzbigU1A+wfcIX5P0okNEMgohWzaiIf+FqYb4Y7dr9DZ8PRyISijW9/Atgw5XzMD2Dn5CSODSa
+nnEKjJzgaiUHLoXj6RztsMNR9uktX6nZqmT6/6fh01AjzZoXJ9n46XHCsJkCAPObr03ZffchbpM
NZtdJdxqHbEfn+YMIG/IffAWk5awABcT1RkIPatD4/I9KsoSCgd0tvG5HOsfdo4hbbElxiIBG1dS
tDHYtzC4zL/PRMZAj7UKob0S6q4x+yJx6dRgemnMPqMKAJD/Y3TGKsScXOsFl/Jdd9R8JODpT4GA
ZQnqabRN0953Fimtkhawl+CnFF/wwevPrJygQEupZKAGinO7OcaDYJVbMUxSHBymj4xXeZQcS6xg
SuTds9RR1h8qkDLP7lyo+9X0nx9pvhQn4K+nLq9BW9z/Yz/ihfwDHrkcmIwbapezWNj7dF/S5mSa
PoW9CifIey5jV7XkGkdJCgIIVNJCmPllFTpifxgF1XmoaC8IWD86jWPqzU41m7FMstUYUhzjSMdU
PQBKTZEkLnNBkAtxqB7pP7zToDlU+v7xkqT5Mdez33H9hoaikdq+VcmoS81S3DfGoAR5p4UMIX3R
y2Hjfcrnt3WSzVUKWFn62/U5nA/cyR7HGqdPkmEUvCN1KciCpa2d66UEAPAnz2NsdNhliKb6tTgd
YFdFu/Mh/8nBfqxpHrO4X5nj2O56KorsC1TZ9plIwmHen+3s21hdlgnsSvLAINEAWgWZ01/IJsha
9hPP6rpo1omN4oL6351E9ShVIxDfqTUNUsVMgP1kE6oFfIsVAhewZ4JvMCSYiynXZkYPTGA8VpFL
XZcmOFx8CTSWxiwLDmhRKwmIjwW5sNV7mDsKOMZ30aGlS6JN6w63ADSZE/pW41fI/7PyFl/1E8Cn
HYh16k4NCJRADlea3/gMPIN/nRV0CxYr68kVYGvDzzP8dltak2koyQ/nVTqIMU0h+wJUQNPZXcro
79sYYdyGD4GirjUtnJAvBxtCcVCHbFJcbu4kHgUM0wXDYqagTqIaRYTYwkPsv1syPkHhlLaLbDhv
0InXpF9OmzETJ9gIKgSxhp5DRMPCRz44idafNussSTLLpXEDL8LdQv/S5Ic/qcR/EB9Y85m8fo6u
b4uNBZ7mXHc9+a0punVfBc/c39g4bPQ3dDVYZHmJq124P4BisE34tde+IosHAF1yfWp9p9dv6+oe
7SzGW4BIawH19FM+/YS+SMCbDSgqRUcrO3JWm8/9bF6CSOVBPUcknCoq4hXnc7fqPGcjvE8Wce8L
e+uAIKJu3R0IZDRVZqKdLLuxxQk+KQvekCCF+dMZlyRpgdj3EguXCxcVhvxktXfBJti3RktSHV6l
mVqnIk9ViYQBGnJPZxD+Gn/y/M8qRulwcRqUq6RqLZDpx94cCMSUFHFGL/2aAi+vUwADQIt47pp9
POz25vI93ZRUt2sL+UdaHxIR/mCyFtWQWTCifhq10muVZKcFNbfjQB8ihXCaqDvaYaeKZiEdI9EB
qG5M/4kwzBrn8p2I7V2fh8igrtNcPyulHdNQnRQdy8MRur0mi5VfHlT+oQdbkWqcxzyxF82/+BsZ
N7eLP1QpBdexJV3Xh7NTgmUL0MfxMsHKKKqT7O5sXcELDgncfKaV2WzoLBO+4cMomnfJzajQRHA6
9TZZwU6tCgnYvRKzR2bHarKuwxU1pCjzPJOP1T4mcthkztvPvMiIkeTJcZY0SH9rX687N5h+BCzY
Ji3ftKv1ssikqY/wOiv8PAHXKv4Y+5NquvbtZU+JC5UbHCNm25BUAThskhfp9aBZc0kv5W5hDcTj
gPRdz5h17LYAA5/AITyOW16gc7R903GnAblYvaZvM3dic8GcfMNLgOCXpQwX5mw2oeV9FXWPxK1R
M6es1zZzeMWNrSqPY/gDR+0yoP5cZ+VGGfoCSAb2O2eGvZSVI6WcMGm9gl5SWX+nNYnOfxQMn7ll
695UCTD/XWACDDkCVRs4aMJcoQIA5J7ISCu66D45w3Gas7lUXkjZwHfCvzhXLCXp4HiaVubR8drL
CH4tO7tlBiFv1qx4SW0JlxrJNWBM+qT3bRDssxOZISnIcOGTah567Lt0pe2D/gHKCbMZ06xbin/J
8hxP3wrFsI0phtTueUNlOy2K1KMQ3LHVj2qQor4yeRAPFnt0EueszQJSBdDWVxSk4I20xxv2jjvl
PF+tLO5R0ZUtV3hUnuqviNvjvcqLotE+Cfx4viQc/THdqueqQ330IJMvvhi4TCIJjhAsL7xP7Bu9
FduhcDNqAjsRyeu378frgjezJ/xMcMiFmT4qglC/FOk1KhVXivcCC9E9N2ufrH3rnS5cMQHsd9Mk
+jXYhwZpIywzogsLV50xpr/hnWt0CL9Dj59zfimp5YSlwF55o3dMckN7KxolgSKtk08W4IeKmEkk
o3x18fkEkpX4ls94bgXIXE5gH5nZxQeSZKrYM01MLH4gY/lYuyjep+FPhFvktzuRuPowAVOgfbJl
rjNR3dYBhzgIG8mE2kqutcK57c+8if+3illWkMWTJi7cZ+Q2P2/tX+B8OH7D2wAhZKu7O0hvodEC
gLWjHKjAC/SnkTChRxDmnWCfWlLMGm9wAllvyQ7LWK8MFyk7zTVMGFhX4ogAKK0uPQKUdXANraBp
MdjbjBkgnHWtTYTQdebptJrZbOQMOpMVFXdo9WcKE2n2zyejudegoO5113bO7ZI7LnvkqkobG10R
in3l5EfrfsNd6CL4QS/KacMnSvfXIpYkqZNbJOW4fmzhuzKKpP+3hlNQ02+IHrZcgxkka4NuO1Z6
xgAHCVy0adXgCQ5bDhRzejlHscme5gq5DQcU52p/OV36dk+ZLwUuMtOeyz4em9gmyb4Ma7ITmU0g
UEKL3IBDLPOGVCufzztg/9gQqUkBx2GjWJ1KFSG56qWQY73tGC1KGzqq5yB1N8Sn4X/WG+iJXhqu
LBLSUHJMHi/hcnxsZoF+q8A/cm+Y4qoJaRF8KNE4nzNLtslD00wGtlovkBwBmfKKHEtVWYLtKCZa
zNSMKDJ/wXohpaQrvig5jjOJ4jqfCsi71lO02mVIgB0nlpsvo5YMsG0Zzc1TrFNvh7FOkNIO0ygQ
56cD2Ppiiam+CGQjVuNTu+dY+1OGGADBTqi4AYpLSArSFXQi7cgm8BOavPOsGkXfD+2677w0J9F2
NLazRADrLinCOTvLoJVd2Ya1nImXKrqaDz/D46ft0f4lHr/geK2ACzVUouGnS/VXwRt84dR8Aze1
X5numFgWDNFFxDlPKVGstYeFD+qsGCuMeB3ew+IN82hcKYLzQJt7F2vU7/+KJXVl9BazZdXsmqlF
IKfHZlaDuGkx66CgrLae2XUdulJnrzOHLAs4nTBPj/c5FdVCnMzpSJeFSgrWq2Un3JK0UQe+JtjD
B6lGi+fM3NWEVnM+xTZEtT/b+VjaAQhAu1IoNfxULzIYjKOwLAxYdEaTAZuL0cWY983iko0C9Id5
ZxzdURwP0VWkshSysts3B0wL7Qmk/reA4ld3uTuIEk2zGj4vhJ2CZbhDX7e4QWcW+X0LrwGwcNAF
emTZFuDJ88jNTQFduq3Y6UDsVF8SqONG0eovZwjUUUEIumBQVYgatSQaKl3yONZX6PVerZfE3RyD
27ExHXgjQ5P5DxyVh/DeamYljgvH8rVZzelzYDuKvPkWS9/IIKa6sxiBPMSjI0MrB+BqX4cgn7Fc
+JOVOEP6kwjR2S3bjH+ohAXBrqHbnAlyq4JWLQeBMD2+zPlKSMDuBZiGJ60k36Y4agLOCt3zjKzI
VuSzrC/8Ki8Qj+aSzavFZFHEELBKSOjeMN45LATdsql/JFi0zSPmjhF7TgWDl0kSkneIs94xbkwj
V3gSnyaoEf6eohdJ34S+008pyDZ62goJ8K2+34YFRXImw96UQNndPmEltwnckkNr/1WRZYRDwXnr
h1hM78/3bFUgUFPHfdymUpiNf5m5W/Mi2scTA3efGWOrKZEMV/QJvS0GB5H/AvI1tNqXvX5P6KNv
/f08FQd4kin0v9gfNS62JDUyst2Tra13cizmWz3uP/D39Q15ykUTFCOC+CxXh++wQ3syf/UBOIit
oW48zhXaImFGrzmUDz3PutwOflzzCLHBsnQ+/3pVCvnVRkgpeYgvciRPZQzK5U8MF6QA0b+/P0Gq
WyDjSSGEBH4Xz8Te7tcmO+WqbHuASsLYP3hDzvzlDNcrLFAI/ZEnS6MzzrvkeZUjnjhvICyF6Q04
M7QcC25hhmDPJF2cJL0a5UKzMNqpPQJd2dweNNFBjUILouwBqk1NyCPs9mqTeysnlbl0I11r4tHQ
R63vIvukUglA/6hheUn08i1wAvIJXRryky5L10rDStXLMtEQR3WS3kfmDUqz6I2IAHm5F3Tepo99
vbXPmIhkAjHHYcxl/m5c/ERo1337jyyDr00IKjbGGH40hGWsNJRWRqkHwgI80FdofbQt/xIk45h9
Lshd9Tbdbjm4j3xqhsiZAumU5IYjWnED9GJ+X0MXsngXpejIUnxhHbdsNs/Tf6HHPUVXpzPZ1P12
kxl+MDGCndl1TKsiCkWIxlEaD8TzsmG9DJdhy7Oh2Bamj38P7ZVbGoyuKZmAdfCpka0YdoNUiAo9
+e6wYROnIT+qmM96GUCw6gFVmwyngl3vmforrHGtN2qbdM3QHXHSQxL1RqrFyL35BjVo+Isbmrek
qhfDdjeWzxHhvyWBziQurV10tzXOC9nzYRuuxUk/W2gd0gU3nGRF1JuIpjcNp+6rXDYl1e+jha4L
hXKhp1JV05m/YFt8XIJws4/+wa96CttcLx3oIUFiaInFWCB8vAu7CiuojIdfyswMhy1Ebs5qM5Hw
Gkb9dlSPu39s2Z4dwzqxtrKVcl11XYsfk5LmmVJgsQrL5lV2o4tx0PCOUrq8INoiWo7xcqkAvE1p
MXomCGTr50sktxBazFV6LBP2JWV2O9GNNJjENWxy1FmhajO7ABbsEQHeJmgNWOisxR3Mg0PyEp95
5YuiW54OMcCEIkSV0OLNXKXqqXsHliyw1bLN28mcMkkkYa8Nu7mKlna7EECBx32uGsaMsZsVflzd
9lbVU3iOX9J1iBGjZa2E+R7lmQRd7U2YiOz2fYrtf0Ncut7SWNRz9FlMGCHBO6Aoi9ACeuf1xemz
phcUqnQJv3EODeilyaJSmO0t0/ezR9L98WN9V48l/rdzreKqLV9pgRjbf7O0DzqVLOgIzPPAE8UO
iHGcc0xvROiyePlOT0p//PTqz1o9OAUwcr20HD4MYCzXUgHsEeFcWaC+/avsuCSQkJyKdSienOnl
paVybZNbfYp5WhGIAl+Qx+2tz3OZaXuuFlU7UgCo5lSxz0OKOZcPPK7EeHgEMnoh/AQ4zDpqlKyR
6+oCbB7gvKFwq0QGt33bc7AuR7dctHRK18JWGz8XX8cGqbARdHaoxPpvYT+hcnqr3PvI34vU1HGo
8oW0qOE6ZOQroftaJC5RrLETjEF+E72p8FOteVloC+6/dentyZ7u33XtmPjutTTsMeqY2pFpBGhT
x4xK8s/rrVdnEkCL2l6Qu5mWY7lza7dn4DVZzblyn6x7n+DNjM5lZMMg3dMQy7Eg2YCXlCL8uBIe
XH/2eayGt1eDLPk9RosuUCORKPVWNFHiMguBf04kC09cn2LQ+LX1yjnDC+5a2EEz/hmZpfmEKEVG
UYzvQKteg5lmigiuiE9e5WRH8aWKf8RGBBgNplSZfur/EIiYB5w0kc2nLlYQauD17PbLH/9wKQIC
al76Fb4lC2C+wy5T96bLbUxgW2QXKIO5ZH7YswfQOsa0K9H0QV7zB+0zeadDKUBrySpy+TV8nJdr
1aq2r7hfJI0yBn1jtPvV6QyasCtY/gV0njp54FvPSqxu0hQQx/MrWmT2JpGkCwUfOrvDxk7+GpCq
VUgl7lTTCJDmBuQKFArNgkeNq/ZqQL/0x0jUqtx57I9Y8ZcVbyqDPQTwMySuwsdvNQe5JnoD+Ilq
l3ta3NHEPUTx+d1N8UZcdukM5QKnXzdvFW6qz7gdFvXdSUAMFbaHKqxqhBjoiZ6QFNBIifqHHzOl
pSUf9osiSCuInhqlAEwz21hPwikUyWC+CXvOw3gD2w8tgV4BMq9Dm3u8sbv8lZJffOSCM+7fFqEN
Zs19g4gCjVyARPxv2ZH5ZIFSMglgm2EssYU+5VP9mgVNCQcv6sV6Ik98K4pfN590pkB7y8mTfvf0
knMZN3/qfhXNljjEvh5Kt9YJBDxOfqum6Q6jcsQSISdMyv/dBsA2nNm/lvJKKFroua2nJWWvhzIT
OUg4Q/SR6zhHVn8XMMS/qriuSn9+dDf2Xp59UqEbI0ksaQ7qiGupSpX60v4y3Df0fSqoYHXQ0wax
bP6fMcsxgt15x3LHSaXU2dwb1O8/kf53ZX/5o6rkbmix3YySvSdhFuc6NU0UW1YUP/jPqG9EIzwG
VAH5/idifvBgyVvDoQ6ALV1z25RL0XstLipfD8lZDNNkuWjGObz/D6bMn+4L8TqNpH0y3T6X8DUN
4rICRBtsRnezyKk9O8BHDNLsv1ifoAmdFfbcs5oXLU4m48DtiYWQ/PHXqBYngvjxn6kVHHYHGSwt
2EwD/wiK8doAyN/2QD1jXrPjtwRimK2+OCRtjjYmcHaWEDpKRsdx4k/ATyla+Jtmq0I2HOvu81fX
Uixn+yEPaJ/k7Cs7Q6IbsANNZAj2s/uT29SquFhotNpuVp8XrkcqyhicWNyKWeTCWS3Nv/UvRAh8
vTznY9yB4FYa37ccZg4EikHaQGQlAow6518VRib6u2gxgaUfcf02Z6k5ShZVJryXzS6D82aoGROt
yBvzLbngn598ov2nTczW2x05rfGPteHjic+q6CT7b1UtIMtvhZqWnuh9+UgPf7bGBdR44psCKmsW
bsqqBUiOQiZfIwDBAQ9z8h3rrm8fMtFyUZWN7xUL3W9HehjJRdVQWzukzVSnJo1A6fwWgPHEk0AX
nA1GUgNQ7lMXnh8f4xIEgeblLUlGWjJnxAnbMOOffr0ODpFdaHwOhVY3368nlJ/1sn2h0zspH1VW
93BvxR2EQAtGlTRqloWiQsuTaoMvArUI14sUhFYWAUruaN0ls5VRLobkAHCeNrhaZ9WxAphTxnJm
14+ehGR3aMHpF+ul2TT+1jPl/X9+C7kGHALRB+tntV5gHp+ahpqAsVu7nY1emTuq41oST+dtXT9j
ogx3yA60cjFO329+eDShihIAkFtWCabGkyTW5K07toyYdkIGZdWgjYEqCQ19HsIZ0QMJJgXAwANP
IWAh3WxVABqC6CY3MTs5sJ0FYZN76NJFQ3uuOlO7NMtd8e7WPu2bAH/OsYAMCfWe0ap+mUfXJP//
ezFSS876TMVsirIzUezP3WWLtebY3J9z5o3FIS6PBOXdGUPyMCQtKwu0FVrCYRZoLwQcSm0rJCO7
6VxVR4Ms4CMNAIu7llZ/kFQNX6nHZsXaLTvsNFbYZ6XSUDV04XUX8tsoJ8SifnkAMM6816IpfRsx
rJI1Qq5qIFMLUrFl0UhGf7MH0Vk2WIoR4y3hwytgTVvuWRVUMMs7Qw7LdhKq3JScWzYjQspbVSex
0HytPRGfwVUFFCPCNRwYx4dzajq3DyuUdkFMpnmzrzZw7FwYTrNKqBCbSSLx0GgWwPgsQ1IRaYmM
/D9c3GrjV5PKT0h2q1980yVpJzfxydGTQShTIgT+zFJd78NMJ3Fx4OPQn+xYic4PSoKkLV9Psjuo
gsjq0i2LAFaeJ4ExmGC3QdsJ1OMrzFKn5NuU2i+7jES3pKo/huh3fiAstAzeT15/h/BjAKZrqCtP
4mZHRJVc7e/83qY+ezTeEUNgSwU8Mca0REw9ZwkQ+epR065arrvKeRKFm4tEHzDKn7hjyCD7N2l+
JZ+YPZbOq4UNQCbPl7QECiTew504GQRk+l/x8vO2IfJNgQCJBHGK+sIY9XdYC3jPayjZv1T9gyLi
gDPNtCUJxmw/Ej4M150E15AZWdwg5CPVBRXMBMetLsiJm8vkgi4EqDDcB4SP4veNUVrq/mydTnFK
1gc3gLKeDtNlJ1PiF6PYRGEqLqDx5E9A0RLUBkzr50p/IaECjl4a/QtzC2sxMUv4bZJ9um+1fIdz
IEsHeBA/MOKNt/AZGa3PQlnAcR3BhGa1gMdXt6UAtFRcsEE4lthDDKT5wqr18QRBQjrmqdDl9qc9
5oA02ej1H6BJVJ5vvZBMXQF1FLPkoHwfJ1NHEX8lBbtldG1I88eWM6Aeu1bcVXrDdEp62VDgSbnN
HGc1Lrnp4rmrDrlGFZNz0EnbVIMAiZ0DyMxa0TLz3OAtrYNr3cN80Zht/1OOcfG8SqnT2NTBJU/1
1Pu+pksFbxvGfC/6E3fAHwMwUVgzdl8w45djCqmjptTVbzqkP3aFWPIco5T0FXfh/txEpIpb4LCn
if6q2+x77/nJAWWK766R2a0dLCNdGXveNcM84kC2TucRdq3Gedq8FnuHtxFWrYuPIUvS2C3TOAnF
UR531T2Sa8oQA6m28GiiQiKKwtarf1942tB1pcCkqWDoP93XySPk9Wa1P9BxzxTFYizxK8ZqFwfq
RfgaXIypvD2cvcx2Mrd2uqRFQ7CVRgjSdfJoaRVDzemrYtM+phtaNbM7boLGNM2P7Vo6N4p8EWZQ
cZNC0JylaNOpM69+ornHjTqB+ghrDOHNpS9QlQqoZ3n5T1pZAHFr5OGnpC7dFUm/+J3RcUDiwXjE
8bCckc1DSYifgnSxEkPLouqrD7PDULcYC6r8uro5O666Mz6Y//7byygN5UMN7kdZrtCjVCJTyCLE
qBAzgiip4TZGz+SBshHGCyCAR7Ug9aHXXXF4MYxOyCggz2+PDNHXl14Wc2lrySNfKVG1nHt1PT9T
lO92LdDnypjz94F/jdoodONe+Hyt9eGvjmrAbvlo4LsJWbpJTFzZ+hFLyx2a/KPiHmnToHx+o8TB
R8I2mJnzWTpCcxVgJCpfYvttUEZMn00nGviblwfbXzHGce1sMzZuEXvMfoEWAQ0Liv7ssyfCIgsK
/ly4yDu8O4Gd0m49Iemue8tHIH6hpjPR0vlZEqGW3fSFGbTWVhBN5wfgFZ1vHSsebgC90hybp5LQ
Ehpcdtbo+q+cjU2WsZ7mRcXNv3JkAYkJEniO4MTPQyUmqrxxgIF36N7UHCDuBaeijuYWV9vUDkTi
O8q6eHWvVkuU8BhQBhphXpxaONf22rgcGQdeIx5Lw3O5fPu7HI6mZjfjCgFC+3TEKCQg62TDgrrb
kwRTjnmzHCMkxArXr/R3YnWEbiBYHwFgQy769Fsizyd9wHvYVUY/GotSdPGPBMGmxrjTiPr19CGY
cIdKS31JATKLaDCoNN4lEOUkVcq39zNaMqvOaNFD9ysTt3erg6ZaLHGFBcc/bjNJwnTIR8JfzjMd
nxK+Ghf/WBRaop8VVnutqDzFfhZJTPcmHBZJSu5I1qy4MPlCc+YD7wlCHdLAT6BauTMUT2fSYoej
6T1eQf7BWbWGXhQWWxP+CujaTTQNeKQPdPfysaXNMlxMtGEftqe4ZQXqo9zC5IV8rxkKjkTuSVtE
iBEfhaMb1vZmqAHZSP6OZO2oI2QLFxjJ9zof20W1LMOagR5JoRN4D3bkaxRRbQbQjV2qL9Rj0cRQ
gX0Klg92pGkSIWfwKTlKccsaiYbvcWSQP3n30GoJ7yvpqumIXOFbdyDWxeXY25dNJblHBde1A5q8
7FRGFegqILrm8nSnelNAKIVu58H0Oaddp75iRK5wBz9VwnE7KB69201FUtG7acXy6P7allZOORdV
nVpiEK8eym4a2Cb1Nfl5ngvRW/TdRSv834m7i4GqA0C5k5GM2KsLe1fgyagkXk2CigapdtURc0zq
J6Z0s26+Qys9VuhenWi/3NQim1TuU/lwXjG+7UOzxadH0/AgUlRPGOltTXkrErBJYYifneQ1JNXb
yYjDV1bhcOizDXt7l7RhIqbgutHBLVa23vc8Jo0t/YEy2K7UsD41y8e1R6DQ6VAAwhqR2JJPaJlV
vforRJVUFq5oWoqef6HtFXPVqXijJiAYILLY5zF2BIRTKSWlf8dGSH541qD70Axn87cAQ+LorGET
1f1HJPHEgMEy4VB6MkEFw50VlUPcBv0uQeRENKU42MCiXSIVNsE0iZYGYjOHhRXsR5aeLO1ONo8X
MlQ+ky09mQwtBb1tk2SMusYmq2rB64BbNQ127tzTMFfs8QVC+bNXTiwpZsWsY5FB438ZWPCHGNWJ
D8ZfVQzmtiTcAlpjnfiMBdcZ535LvJp4yiicA+YF1TlUfkfVmluPdtTK5MPXSOjLWbheFm0JOTKc
1dQd3hXNj3SEXctxsoAyAanwEbQsb0dI2lAe2HJ+KPdzv4RmcS/+1dkhReSFZaOI5RYHxYcroHue
WH85SrP4KLRAqosYdgNnYYSZe8MRgYovik1iHsDC4NehnpcSOv2vAJVxSKy2PsfR8tRSuhO6JGAJ
jfjsaG5SIL4Dl3gByAw4ZilDUlLcdm+vxW8oXrIbs9ZNw+4s9ygk4X0n8VOiEBEWaR7lekzz+P32
sQeL2LZz1jurnUA+azTUVoRdPETossGRBUEC6xGijzf0zLFq8GZHyOC+520velvLL6dpiLHfhhk3
UHCgsOrslpF4rJLGV5LWKIoMZXhHQDcGJ5Wt6oMbD3HIF+gdh53BzI4e74lmqmhtlB8LoDEwf7xk
lL7BL+wRUzHfghguTIezkfYwjQi+3RbcI5L1RjMQktlvmJe462L1MrRWPpB2iruyuRH+BsZhfNZ+
sT9hbcnexi3Q2T3QY7cOmcHaHI6zNxyhIZoAMK3M02L4NU0YKn/20J4+aYku3QCrXx/dyvcEeOGS
wYbm3VkTA0cHic4IRN/JqOjJA1xsCAgISzR/cjfG2H/E5S0yYMVCZ2dkd4bLqc2IeSsdzWoGGmxz
6tPpXgIkeGon9EtACnWp/BTPBGCwDMdo9q5S/xdsmjGo7RXog9978pCAuf6ruw2HBrJ3DL4jE80I
UYxIJpGW0f6Ht5wH6C4rROpZO6G3ZbxWuSCjO5sEhhz79T95lMrnD2BFvmNBcHB0ekORsF4QorhZ
F92BTwdZXDJRTRv45iuqZmjpy0nAZGBs/fsYSXVE8vMbRIGlQu9vPJZhfrfkeG4Av5wETG/gTdhd
5GNytuy2yLIFLe8iHilhUhscoVctDRIEuRg/sTAchdr0Pm27XnxH7hHm+vZVrIDpjUwY5RS6OM//
Z0kCmQ6QLOTVBk8YVwDxnitJ1Lw+ihAjS4RdXIVAzpP/M+6hRXUQnL074ykmtplfSrPVT81/BYT3
GS1rNUUcKt3LxzUXEI+BJRP9SvImkVAWsmcCs+YrxXUVyiBqIcoHgdmztq37flT30lgiAdMBgw4L
fUe3C25OzuIqHca1hT0/O2P992Dihl8kQPYVXVE/2KufVcQg4QaDEESJOXhFy+Lp02ORGRhYAC8D
eAuCV4LkDWU91oPyzGoYjyTXfOvWLXfOPv9itopNnDf4nHmKQyMnFri/8mllV+MIU00ClZ+NfM8y
RjHHEOXl5apQ+fV/lLqp9WBuwVzYZ6VNpoHaXSEMYMpTPA3PnLklhD0OTtfKnAZ1NXBWtpS2F0cb
PXW/UEb/WwBSsPbdfOKdeS2444ql/n9TTKvJsaq+xU+k7eHKK3c6jxEQNH01OSXeCGZF6nHXecRG
XT7FskDPswy9yBizVCGsmWByQxn4RlKoDaRR9C5RYcRYS01gjUd5rE+Zs4GRVp7On3SB17d2T2Me
v7Wot18RRYcyvWQnITNFcTV0MqZtinlABuZCSW0ZUiGUxh853jQ0GuopClhegy+TzmQYtH9UCnu5
9JiSaUTklwCBODmFGQpW/dKiyqncoX2m38P8e21HRnq4keQlNn1VWbXtCDaMH6jH1EmVhoHzJfdm
oppF2i1a9AW+nB1LDpAivoiKejP/0sWaY5aww2D/gytUvLFZhST9TIGJ5zxodKiZdkTxJ0lwF7gS
W/LyBv+YNW4sSwZW374AK4eHoeXTUhKWup+AngJkz8F+CVda7bLFfMZ0qxl7juEP+LEeW64J+Q/E
TcKBPKNjMd3tXGEamZH0lWtpA6TkYbw2ppuCNbup1An9Hy/VVvvHDO0wXHm9iDPPlYHK6inNfI62
OD2ovazLuR7X+T6zqUMBZ0jy0UsMvAZuVLrZSxeKUHimi6l/5A6z/0SX9b4ZOBKh0AHK8AMPKbL1
YHQO3wK71vKntYQkFb7FK51Bwfb+tLvbtj/wSFwDFSkeDbt2r9igM2tYnuNGiSnDHufrwvciV5HQ
YRZFRFV1zmZH/ZD0PBOhWdMMaSJ2NFVyUygMG7GadwnM4tQqcGcwtqtmqLqp1lcCLZxNCcGF8X3F
cpYZsOOniVy2sWxSt4At4iikpvVwu+LVw1Su6T/l82l74GF7lO2N1dqZq9tsNirY3MfZwmqOGsJM
OiXSptVhCQ9fkzOCIMTzgmaHWMXMn8+i+CFdaHmZQT26WFGDEt6Z7taXUJVVKtuCHAteHLFQ9gMv
1YEVQYG68M5WET2s3oHmIQs4la9DISU4HWb15l/+HyODSx/Z3lqgTp57oNtypkJl0/ehMfd75+I4
J1ZdOsumVebkBGByy8pzX6zuEq3BrHWoadGHh2fUZ/U1mIKG/BvMVwsKDJppB2FYZUfSKFrsmOLK
fh1uA6FdVBS6sgbd53AitVBxdPI09IUw5kK1cANm+TUR1FEYMcKQTeulRX7zNOoFS56D/bjRV6wn
nX1JaGgbYXMZ68bcbvRPdpT5QcIpj0KTza3a4iswW9VOnskbA/jVzuYK2fQOXWjoundOJxuncZzz
1G54vE2rc8q0Wt0AbkyEWrKiUY9ZkckrSgwfQnZTBny2d/0Zx+qtDiwYk9pFSMBaqU9O9dbVZIw8
hWGuVNwuNdTPuTe2xIve1oBwlav9fgRGyh199Q4Na/Za1jfZWHSyTE+ROObb5ICpk/mf8QPYzXlk
/xH9sFWdvwc283F/1J+h6LMkgL75mdcGy7jZi8bevqWqc9I8C4N162B9kDVYoNfl2+xwdU/E55Ir
9dJiuczBKaUYKzG9C61fH8FaanEoV3ZfoA0GXazJfi9AR0y8ieKV1TWYhkreUCx9fcGXsQBo9wvN
tRFJjqtFMn2ZXN0+6OVnB2dPZ/CmAloqsKLbN1oyWGXN/2HGyXW8dsB1Wlpz7oZGBbExbLtTCzdT
aXUoc8G93smoI9iUMQPJIbyCfm/i+gexijXUquF77R7o4wCxduakJ8dLaup7El11DzCDJnmYte8f
WDJmpTemDLMoK5t91bPoQX+Syp0C6wU0vjorBo9XbyOP2UB7UysjDLv7hbrkxg9Da9+Ayao1b1B3
j43XdtcOk+9y7WRZbpUMv0JVfeKPjBvxtWkUmz0/9AMdzV5idQ2hcdDa927xJZy8Tp7EdpdEGx5Z
1ZSeRqQBgUtS7j8EMEpJmJNqJL+YweeS6WSGD8BsSBumxewMuTpCBVyB+UwWF0bnKmDRroyRzYpN
gSjUBXjGuEhR7iplAU/PPYZPXfLPjAXaKi8MZwP9uAJ3qOTdWW1FHtSCmdRXH1oAny1u2OZp9Pwy
GUU56/rQF9zP3rLv3Fkzoq3lpF+eGuQ3WhryTgm/nML8ygpjXDAp3XuvuIOz+5VX8zC4pxfnKitq
k/uuLZQEgZ3G8Mh+fZprRxvsEnG1CJ6bmWXwwS492XtLw1CEB7EMUr9h6kpmSZFu3aFrnkuQdrXg
59Hhfin0xTxFUYcz8ijqMP7lhuAlasY7OYv1/j0dUqRmq/9/FDdPn0JkoFuOLK6kRezHqq21RLQH
ol3K41Jc2Tdf/ZigSQkmqKumw9S4yNzvSj9lAjm1bggfzdY7YercArqtxe55PXQhZArz8kDdJPjG
F1AwoLd4+aqiCLUxvcQlV2XycBHkeq5iTkMDg35WUAriWV+c2MiH1JsMUag7YOFKlNhFBe/uQWR0
Ut7qRppDGuBv1UUO4h0VR+O5zUBcmnn91EFYd4ih+9gN4PBiblFMR1n7TWVfB7O4bU55aj5iJ2LU
UTpQhIpocULVesTqirmwMLOnUYpqJ5XJf8IRpJv+G/fcRLkT6WDobGjV02hAFyagPPS3GRg2sKrd
nf8PBiAKYw6aGcJ+x+WSljAhUg9LvuXJ21ztShM9FiMP8E+u7dVI9B7xls0XHWLvnF0t+EZHGXXi
BZlg/hnDaHclv5tKYJtX4DdPALepz1Gnfi3iYBtIU8ThyRV9VgX1P9TzUmmLqZtzbpXh7PmfOCJK
0dexPlPQlKbQeKctzFB4WUcOCPrMvY7P8VkOUq93ueftyJkFk/+s99hpCtopaYM6Z7ixahsejesW
Fji+GBvCVzSCwpPLcUn7JUXgfirklDGA4podi+WYfKscdMfF3j8rexmTXQyU5x/FG0RP+V6DfNgg
//8/dKjIhs+C9VmG2AC2RxFWk4zq0k3nuzE0K6OVEZ069wBurAIu65wgwKgqFdzovHI5TjLL1oWk
TZSKpL6tl+Mp3D//dQOC5BxSgYYrtQIHN09BLHh7sdVLtkYI7X4gaVq5L7R08GAs21PHmI2GDcGw
GepUeM7BHRyqQWyOuSPcwQmcC2xV+UfC3+7evdN+D7+afA2KNO/U+S066/YFSXK3lGAJXhTnmkOj
ez7M39fFcSohShCHJFglIVDx7UXPOU4sFraca/sMinJJSSgS0U0pFJ8U/Z8EJmZLhfl8cpy/Xqzy
oZhYf07NreM5h8SeIVLcy1HwVnsO4d8QtSHuM54WSz2VlbQqqNt6cfHJaZ1eiROZVuuUwp6lFeQW
VBirxmA0owRyGFsBPaXhbWL54mrdsCtTUentW9BbTjRZf8ByQSbifiRO87koVpiWwrOMy0vSE/2Z
F9SaUYMBUf90dnRZ84IFPrj8cLMXIbtxybQkrzX8zS8tr9PAsDh9vPe9Lt2rBqVn7OQaIaeeayvi
QngLu8Z9tLwtdhqGR/QO2ND7dE9Q5wDIt+YKMiSAkQZb3kRpvw3Y5olLKHvV0yYzXZB2z3CsrHR7
uqr+QvsNSitY4yjKgvs0gLyniswWm90xupKCGztUe+v52LMP4Quy9f75Y26k1liHWbdEAdowvxWt
drKYrAvAEYr17vvsLRf0OmVuSpX9/gJMdSfI8v2iQVptKs6rOU+5NRIxhJFYjfQV8mkuKLmvxNJs
Qz9QF/IpbVd2y1ov3CFY7p1AB1mgDa+u/QuYbcGCTjLViJALWbvxv1Kg2nSAMg1lR4Trbh8+eLlz
JKqqBIX93dQ8Wmga8AEW7jOdIapoDaxiaAPEHs2JqToHpTXkTdjOk6eIeNPDgd9cOXVrPLxZl/hb
63RBNiXdhyfZ6HUTcBL7qbleeOkaFYbI7l3pR180SO2WwmzeHbSfbSoj5KY8LHtyicIi+YUfSK2J
id9CkE/16VAz9hxhqyvOeff7xWlWepKKZZ4SidcsvujmHLV95plUhJdB+UoS6Vem59yKg6wSpZbF
H/uwa5br+pxheZQ3/p42X+K9gGYzBGRpY+tdHHVZ7ewPJHwN6R34Zhl6UuBVAnTGZ5GxwUK1m9oz
knsIKxU0oYDoaozhy0MY4/pVKZOod93IHuJMUmFj8J9C0YyQjVhkHnyG9VwEuX00Co0RBH4EHPkY
KIJ5P+Akqbfj531DKIK10BBw7peN1br6SKA+EDfSqdZ+ckMKtS1vHZul/Iwjj1B82suH9BJYdQWi
D0qZKaeeXnU991rW17ei7vjjABHLaORqSWgS3h0xq4GwVkSKARdu9/LyNE04FoqvIGyxXwRwmVe/
ChwdYLbUxXgAlRrd1C8Pg0KoYAzm66SzsQnkhSNgFSY7WkbW0tt4bLBKVy8GISj8kfRCh9DUZm+I
itI2kmv4Aw6kAsAworVdAwVYskS6G9l3gXqDdRDKuz435BlDTlcIkXDtk2E1BdwBGIAHzmcAds8C
cKAWyYVHgyCOzojY1FVVaQi0xOVRNDBfhGgkaqbS/STZGJNepcwUQVuzEavc1Yuhm8SuoxMXPSux
UQ2OG9vcPvyel4oOJZTmtv31xINCJb6VfpFBp2uvrH15PcpAtQAN8TmxUQKqFZy0spj9XrdfrgL2
Ju6dm4tPTCJufvKYcjgkVJeWT3PQikreCBiG39iezxGQgWgjeChPbrTCPcqQ3ashmyibThMYU0hp
5t3MhfP4W1Fqpr2NqsgYRQFd8C1wHlsvHC0UmIFZH2IY8cWbnOP49du8eT+M06rfV0STyM9UmNb5
JcNOWnqQFT9SSe10ZAQJ7oTz0rZbUUk92SXfbcipYYt7Mx8xsPikLRfTfQtTx9ygDrkBwhQJVnzp
dvlA36p/56JTEqcoVluQyjU9ErgsuyEFUuva4106Zqei4NjzBeKpjsTJCIV93cyE4tlM6+NcIPGH
/dqvTMyJmivasusuy48BWaKOhGp455Twba359zZOKMFiwNxk6wAhfzM2FCY0n8C4jYaLOnwFmv8e
01v+02e6917lyUwyXm3NcsLLZ5MGYDEqfzreQz4UUtaoNC/s3uQmgvcFM7LaKsN3faxn39nU/6xm
TZWLZ/bvnocopLGVVOrUv3IAwfirkxll3/DcPGpGTZh+1v7WqqVuCCZ2y+e9kDnzLef0jU6JQEeG
i8uWQfWXxBpA8Kpa3lnlOvjGwfcYR1dzHwt6vZlCTM2fv6dRuA9evc+tJucUBxbTsaqK3XhKzV19
rERRpbVNjGFNhXpbw+bSQ+4eI1sb9ROR9HwrORE6uqkRGOY7Y2Y/MIZCjHtfjsjlRf6ES1njUjO7
WyVH3K4ApvTEXbk9DrdDBJfGCrTNXODDAU0Wm2h2KPIKPcQIEyxS/baaL3BwKBD2gzqZ8clWSyOo
c482BdfgZpe80lnmaCG186Qezz5D/4qOHlionDJfyHzbS85mtuElaLd1CfgQVrD/VApcN/ak0TNu
N2TWthKZkUUqwd1yAtBOq23Dj696QapvK/UfEnITEuI+q+P1GfzAY/T177kS7ooGdyij/OeUOXks
rBsl2BECG34RV/q3y9x/p9xfbt/PNfIoOmjFnIPs+tT0pXm4u3WlFnV4BREjLmpbUO645PXRy0GX
v+KITaST4GZuacX1uzFv8k9aEJIhDbKdDxsDHew8nCrBVYhxmluq47YsoNttaJ1BbFZz4kJlQ5iw
ESKHsEEotOlOaTg0axfQGlSNc+T78gs1lHdt6x5RUjffsjvCWWIXiodE4KVtljhfKPNix5pv9bLV
ybGvUGICj6OVLr3960ZuENgJQYBwvzGmgX25Tjgw4/zbuECfm6U0R83C0Ze+E5R4+oa7W/srmYWa
MPPDlUSxGCDJfilwd5y6Oi0r6GonvcNjLOH5fd1NWoTcYfDBCdILQOF9gbmdGE4F8rCqMeibuROv
DmzkHKvhY3owoQGS6H9uTnI0DDSQYH2ZU/G5H0YRCOhkvbMtJFJbaS0NSRCfsqyQGjhjvw2FOr5n
GJESzyjjWe9n0VNR5LSPlSLrEc9H79F9zDqAKwGeBKfdZpTucqTJ+5a/iKnsVUsOzhF2288E2V3a
eDBjMOSjoyAnTwWCENrlvS7Qi0FcFVRrM+XFmkJ/wVGDLsT71ugbrwqag35B2cencjr6jIbJ3YqP
TrEGF/RTsouLx/WUULz1o62g+tvhIRL5Gbsm62bbfXd5E/7+rG2bWFN4NfPWvCeauiMmKphGLPhQ
ZIB7Gcbf3DmpY/578lwKRZ6FuY0haXzr9kZKMfvn2CHXS0gjNUm+X9XCYkSvRfxDHgALJrSeFGAR
0gYZrWZlT5tKmPb2iAevmEwo2D+gJQ8hhHWjmbHWkwSm2MqKy2PmCib5LR1MSm2RZ3rFTvNwgQTd
Ak1VXUFfSDlDzeMkSWLdyhZm56uijs+Mbc5o9Ob8uRXkESzMyW8Kk5vRvoC+SjDz+WSAqqD66ikk
B2Y86ygsdVTTlD4W35lIq5n7XE3YxA2usr3xclL/giKMBzTjKOrdSCaEeu8mnLNV1xPvOO7cHHUM
w/n0ZJuhrDjntXjOUusrLm1CaBc7saW1ueUj69QVBOE05FWnPe6e6d7o/sjMY1yJQR+giWhxM4lN
r4kxn+1h0c1COZ1cDeSKziFqCJkBLf8glew6vZ2QrnvvERFeCLHEATmb1wfTa7it+XOBFdxawiZF
t1sji2tnf52XwZ97mn9qXWySLDBpDp9Nhh7jgLb+IsJS73xvC71PBh3XIUsbyjoNm3kbEzjNUMOH
B6RVpOt1/cZYP9UZOn4bAC3gR1X5au5cgTV3KUpvRBZLtWfE/MPdUkFD8m8Y9aAI0NFAR2qE+dGQ
W667kAQ7DMJnGuLSB1dHrND+6hq98to5k1rak4UmF+UU9JdMnsID402rKokqb4BuUYP3Hzk52KP2
4KIEur9eaDgueJfSk1KPOch/lkon1aHMv6258HJCEB4Quw+whSrE9CkvjjwgqU+0zo9Bn2sO0CT7
1swCKxOZdfeLlejtnoYPfU6Z6Biw2g+M2otQcwBX7iLzCVrHZpBLivPpF14JLhDHpINsnBW+bU5O
lvbh6RGLpPR+SAZPxLODzu4qkHUPrK5gPLLyPGRqq/kA1MhGsbVCmlZKKYuGk4dGPAGIk+rS3CbX
VyrRzBZyoPi3V95QFnRAGaBMdlTL/yv5Ow0ZmJY/HWnOYjgv4cqseBdt/SUCpfrV8gDex985YWVi
PF4TFKScrw7ArNQXnBz++345esfdhGCFB7k4MAhPf9ySVP9G7KlR2IIsQLnRMSKRp7dGwxUk7xxF
nFRC5A+33wCKb6mNxY9x1MFqiuZcvxamc7FIpsqnzMO9PRzWP4kWYkD7TI1DnYYdvOqqCRTdNFbc
Hz/YY/CbW8ChClNeiNTX7jfdj2KTWL1gGhpwit5x/jLMb7oJ4xElmOqQ18SCOBCTKgKvUmt8x+IO
OCQv/Y2aFTk6XmWaxCNJKatR958nsDK2IeClsuRnMQVWTEhms+zZuJSLehek4eXNP9bvnZ4uKhiJ
8eRqm0a0b9NTW5AGCr0AHTeaSRO5yVuRhR6qdM95pfE/js9YrjRtrIIJCz3BYBx+2fummF373OJ0
UzNcWYJDpvRx3i5MWEpJyXbCspQwShI2ITAR/joKxN/KKEMt36r2nxuCQ2t9SNLKNxdIgt8S2XFy
FSvOi9m/sluWNSKIvYkQx18/H0wR1xWqEvCDovWrSVF0I17uoM4GbSMGhJUHB7MbpsOY4bpRcoN5
QfGDljrL1P/qlrEoayf9YdxppXGIA2sc3E/YWmFiLbElEQa/ROYuQUJYeQi+Wgd+qylY5+hZJUit
MljiTWHVAPe+wDOu+vDPV55Bv4uwVkegythzHzUIIBpa1IY8y2rO/0E4RgFybpCVWYp1qODnbGY0
bFPZIHBT/FQHt20Md2G8zNhSUfkszBohRbr0UE8UlvfzV7ipbGI2/sHTkmvHu09763z0CCEOr2kX
xZK2AFQ4AiuSzfwuykg4MOZ2xn7Py3Av52jrDbcjkPs2QEEHrG37ocJuW/DBV/ciPYa4Iuujtj6h
wROrZiKLlG31lAtY47u55GQg3yRm2gE/lF3C1WiFoKJMDdBg0SE1+tqBtFwhrVFJgyEtPR6ZxfqG
Jk2APjYKSxq5ayOXEbDu7dbriJuWnS7HmpK2KVvmMccyThpn1RCHRN7tDUd2YasydL6I1CkJPDvb
1mi8FAIt1sRpvMJUaVY8B5QgFcfzo/n6BaTxEMnfQ4y5ak8Xxdq0bIrvGB92CSkJcEz4tEsPOZOM
L/l8adT538zqL6LUv3jI+5RIfWzDHNXfEYc9NWCU+sBS2rjfNjurCmgfdhRb6jG1Ap7IJqHJSF0p
L8ooNbc4+XoaG15qN2cAeJycHb5PqKuxyECXIF+aOwLNalKhxSkZ1acD/1hAb5wjEJZESp+iZCxs
svcYOtRXtfpDPlQncu4TwAJlXZUn1phkvv75ocsGvWcDWK1rlUSPky667RiKZ/jFLK0eMLKmz1E9
4RBVa0vQNbPvjvLbBpDmyhOUKmb9HNa3lyy97AYAbwdGOg2ZtM2GY6JHis4+0C9+3lPLpz/qc6eP
M+eKCVDgQGv2Q8vmMsWDqSX0L/Ay4+a6MaBXyHdkKA7ifIX6KoJeyMUHkWKCigncznLUzOc1uLn3
Cc4qOkEMw4XbjYMcQiDFNOozq4K7MLskdTbItXy629QFUB24nTDEKCWJfRvPzq3C1gSEgUI2H7oh
G8VCxc/rmzTvtIkOn6pXgEcEJJgZwY1PG9/aPRlh8Q8HswIBx8zgLeWlaVRBwQns8seFzYCWGNa0
CSzVW1q+Td7P0dgMS9TncBdeJ0i38LEyTNY2z/quEg/7WNMsReTri+oLf9XgrIEHHDn4dt5Tipd5
mwKdwEDz9iTF8hfvbZkh7gKFqhozEmBVwBYE9jqqvDijA5ficd5A1LONMQOH7ExTpLZfa96fiwRO
CSpsVO2U+A6zbRBNvVJIjNuCZd7MzY2pZC5iXLHn1MHTNvsXYyb6xliJ33BeGVKah3p9VIjk9jDY
CqA6rGsCqQHrIy0TYooS1dVv60Wb0Fi23bpfjr219LKegftfCKcgHJJu6KRLklvh9R9aVqDaIZzc
Gozup4aZy6WsBI7C8r6rvTwXG6g9/cgU17lo3R7dj8ar7+Ib4jpXUx3RgWcx429hbHm8aFeB21Va
9Gf3fjlG22O0CPpPXSJRMag9E5Uw+jDpgrZ63I2KkRqc9qirUR9xCHXLd8q9SAZT8SSDWms8r5JY
kXdPBWs+NDZZ0gWCOg4ZAOTOX8RQBS6YAJX/RrvD1lKwjT1kIT+8h1MxgT8a26GWT1qIotUTLo9T
ZWyKnhvResza9tpJRA/kA/LXV9vN168DxJcfpEm/c6NGSTCOEo3qPUcvR5BKLt9olrvz70uMAG1K
JB31x47gVxsvhhUdFXyfbjksvtvUs+FZYi+QQEBDflzV6mDKJULR8hyhQUlQ7uPqMfqBkrPlKjsK
y1/+n0dR/SpaPhi34apvnK805MXOZvS8xlrXCWUzNMl3J20TgE8N2derQwRpxc9loSD7Q40X35rn
Iw2T+vSwPaWdkJYtJeYXQT7BrIJeYGbf8vrxiFkMXhbgPKy4Nx9aVkSP8N+8oBeWcPfzlOyhE7Mz
d9+EvWI5Y4G5MMZ4PGnVoS+dGjQzWeIoY9xl7ZwU4ALmT2zKwCsz59GIQ2Uf11A+mmD14E+omkOu
W37ESv8vz5UvUBM9RoUQ7VlfE7ATkzE675oPy1aQwnPZZ68JuWJJkQH8+hokZk74qWM/xCK3PcjZ
j4vNU7PDYfIO2IDKmghpZXUQ5SZXi2x9yXTGJlG6Km7hQ2Stg1XVBEagiWakebWUff6bWHGD4NBa
B80OsjxjK7Lvp3VNyjzYzoUMsyE6SRFLRYfUfrW4Fh7pXn+JUBgOLtIBg6bE5o7XgcDEEfupw2uU
6KDA4DtcvztIutOP48FyGrJzcO47fWkC8VbEoXrLrLqDqpkFcyxoUZLHNqOfgExqlVCmf521oXjv
G+J8fJSKOzfO1UunjDu5a7XFFcRAz/jw9FaJ8q3b/S6i+A1inhWD+f44HFhs+Uthvj2glnXa1VqO
+eS7cx64jjhaE3vCqFFReEV8taNmNFdyOCYjFDNn0O1PC3xs18lEGUryd451OgtmSv3xRlH+Tpzs
pXWkyRFjDBztQwIn7lxzmWSOB/T7xnDlWE7w3yy0tgOjZNGWlZFqdJ28o9Vij4X1t8iGHOWOokl7
Mh3/kZKJDS0UsfW10DVu36T33sLycL8IYk3lWr36qAvU5sJlDH24OpYxWM2IvyDak6GAC2GbjBL5
HoHyXGjrUFa9VJflF8F+eND5nJdaravN/C/9qVER5ABrVOhIUCZ9gzGlFK+SIeGLgNOPzokiaCaw
1NGfzZ+ifIBxTBsE7PZj/GTzvtY5MNs7BIep155f5DQFfj+uNRKDwTe7+4QEHTRE7s429DScV4Ce
JFGBzm8rxbPxp2RaRjuVl6tvJ27OwQdgRnCmdw8fCtDdd2EZ2bNSTtmXivjR1g0yGXj0Fp+CV08k
huvh/YO43u+5CLfifjHJP+Ot/c1vAYnod+ci21BWtAErz+9rYXWzdkRdnoaasMQ0eDD+8l8a7KsF
Lu1EXMeElzgoE/IT12F1Fzuw8Jx1Wf1bvEldkkm2ZamyVmEVwIilLzY4MDAM2xASlZeFo5O4znLJ
8GcgXRRTDCW68yvlG/bPBnbO3/4c6lLjfisJusz4GsHQtaqR0lFHpRJuOSSAjW+7UC//YjtQxcRd
wZHDLN9tMC1soVFVm/dQ9oTfn95AmHtPizXOMIZRgTocrppZJKv/pJAFN69VYosiL33VcX8o+70t
N9CpEmNV0a+CI/WIFzML3RtFRN0hHhO3MeXIm0DDbzh7JRjy9hiCh223w+3jf2TVxfYtzM8cOxGO
I4rK/pWa2inoa5ZighfESxG3ZIgleMSBRX3/COw/w9ad0qk5KWpR3nSP4Cd4fxLYC9dBs8bY3H5A
rM0sA0sx90jq92Vekdehm+/WSHp4Ud+3kydK1QlrkpT3eQWHcJpWUQSn5yUWzQXDDn3wxbRnzHik
li0U5CG/TNqSihaK5jwT3iOOBByi0DpJKooi0kVWTVBhC5fm9yf99QHF5O81BZIK67CH9WeJbA7M
QkVi47VSU+dthg4yW1mZkQBPp2SZ05SmKRprxgIhZL2+HKVOSvXsG0zGzfOfJ4721IQ9ZIBigeKd
hNY9bMj91b+m0lRjStPxIiMbD4JpKgjQZfuc78ffEjvTbKOeCVA8uK7RxK7pCvMM2Ok5TCooQDiA
+nYFB3FQnysiA+0kGyYujPfDttTS4I8f8bpPnzq6pmLGpSgimh7M3LSN8Jj6eMSNuTQYPuIWBpTI
hk98rJxf6hkqCRxFYGN9R6PWaQvJqC4cUoM1TXyd+OXm8lWWaNjQpGf50Bxp+UwhMWGIq9NUr6B2
Heqn4QwbrzFE1Bzz6LVQWelkM4uGjSXHMCfZM4Jv5P1pBYlRfwvQ8o/kar+R9EEubIgb42sVVmYH
7jhQCJ3sN+lKzpbGzOR4LyXftUJwjNSZzo2V9NDA5/5rU71UC5MmTYlX0zIQlXJYsGOTFTAbubQT
7eYJY4dQyNVqR9+zPFSBZX55G5g/9ixPFfHwGVbasBnAl6O+QkVPwr1Lt+CT1SwBOT2UZnihw7Jf
Pjv91ZNL2O0Eqsnvx/0gR4jSIyek+NBvF01fnQicrE5k8Mr8+47uYa7b+AV0TDevOw0C+XV0FyMZ
ajMfXJBtA1UIcWwMaESF7FawuhwhgjZLDt4kbF5Gt/BH0Oyi3jjrXaES3AXKqW0Lip9gDl+POB7n
RoyquxSGwGb4OLSE551QE5RNqy6adGVXgOuVjrh3i1ewu+UNnksbPNt2K5p8wF5sipmiNTV+PrY6
0NKovIBRWf20nvbMWC9SrrAWns6Me47+uuqy4XDlUfN/k6b5pHv+EIq6bIlSgmpAZFWrFU7WUfvI
PV3J3B6dj+BcEQoENOFdG5VKvkT17SDpgnJ7xz8yr0pnImk6FHSuXVYvIbtXC1adJchuQ8ifODtd
srVAB5Hb40CHmAoMcNCKyaxJ0WUeXt0/Tahie7LZB8lsXcHTEWJgyEFZZAkgW4pP9b57PTxoJUFn
a9ykQd8QUQ9v4VfaZjgfj3bm1RydOWLdyIU80f4LdVsxR4v4vPIZO/eU+bwE/3wccW9HrHfDWhDX
RldEsgaQxilg/KK/vaPwGVImZTGIxJQiBRAaFvZHih7FCLRJJgcbrcHL0f1HJctLSEw46pArD0NF
/+CrObVBECohMJZh3zER7pzPjia0sJ/5TkFX52qXHQDfSTevql8VXgDLqtKZ/+Z/h5taUKuhOoDS
vEQJgnCKpjiYj5YtdHZPFefzO0z2FRSSX0sgMJSLuzfQWgxiQnqQMuJiW6ni5NDBQZxvMdYd7HM6
sI1VqVlqi44DuP3wAMFSaVmnzOwwayBh0T51b7L6qt3Mlbw8k4j7VN80KvltR7aEjkCB29w/2n9e
W5DvrCvZv1EjG3zMPT8tyCieAZS+Pd2Ynub1vUGQEYDAVGBruvA8HavU9P8zhzSBaNSzb0tNPedB
yW08oOKaXkD15HCXKiyG5QY5TLE97QqEApUB9s4HEr3ESDxNAXjyh7YjZR8GhACHpe2YmoSWNVSg
FSxpg7PCbBIE3YFdC5yTaaob1/XL3eQUqmTCeKWc4vhUriwgXl7Pu4pKTdWE6TQu0Pgr6q8FHEHu
GrzrpCkMBaHRMyAalPyRw3uj/o+xIs9CVS+Sz4CYUfES4II/Uc159gxMPGwVhWht7lauWP4o29ko
PM1K8bDoaAPmKWVmgPCvVvkYyv4+O7l8+e0zUFKsLWREZrP+usltGRB2cjCCpPVgGdx+87IMpL0P
hs5jQSRQPGFhgV0tTdaOY/EG1pQ9nIIbcfs5bVC0XWy0Iza0x9vElNE77YY9gMPxzToDsyxuccoJ
/R82RFuCsKPgdKMNZY5rU2KEVIuDOWXU5IXegf3R5ho6wyEiboJBTXJtBgNqblf68fvqen7Bs6DD
K1gXGbppIuhJt8B/+zmc6K+YOaJQsDvmCifdCqF/nTnad7emGvyBrwueoCOfVmJE6w+R5w3qQJ86
NdUpGSQLPa/SdX3ZuYxyeTMavBdyFxOKUDzYBw1zeqr+aHjW3sd0GcQ+OUGFn7wHvmfkGaChC/8f
DQkcYamb1lOeH0ROzqxX4ZSXUqoq8tIBzcJlyBfrdW5iZz1Y+j2Sr7Dddjx4pbV2xWKV4VxFp4D/
g2rmmRx6HqtPSn79faJfbuFw1FsRpcMF7y46ChfNUK/sNt1jnlhmqjLoJuCtXLohk7uYsOSeGE4x
y+R7nyzqIOq97V8kvosHAel3o3DmGFUWzBqbXlBrRiYOJPQ+oK3xrKH21cv+7aEldlFuJXIJTrrT
pAlZcpJmsGYH1c1Ko1tjLSDUHNAoesNOH1WJncLdjY1LWbm2kUGkjZRwfgldUcewMUkl7aPhNDq1
yY7VyG2B1fNkfmj5WO32g1tTV7dlU3dhRUxo8umChiRaXwTdzzzctbIj5qqrFAVd3OjJm8Yq4GPC
RAWRc4SI0bLZk/iSsXDkFxELBP4tNDuEZUw30h+IhbBpggrEfgoVVTx6DQD6wq+HLbeJ50CtjpZK
IlmPk73k7amHp0wLOuwkYsYzu2IHBRNv4vAhgQvHHZ/5rqYuzXy+OfCxbOHC/OffQ/8AG3ew8TBZ
oYzkcozFePrusBhhSHC5FDjsA1Pr+eivitLij6AlbvRbIpZrYkJgsi5XTccT5wFa03Iu38MRCtUJ
w9j6EBFOwlQPbDTEbn6ixE9Bp2qIDpCrBOgYxqLM17qYfqpltABeG+DIGq0bpwlqMamyFsbLNKWP
vUXcvV9FabJ/Ny4not7liYjNbgm/JQPIa0hZisLHXROjHrH6d90845LEItgVU0S02nX8Wehofy2s
LbxwsgT6av+Hwqo4scanSjpajBJwtP6ZhFYT9/vY9RFFBvVY2panDuzP0b/C1H4T24pDyiob/4Cf
IWGtR/XhwatyhjDRakCfMFxdeOj6xCycVPrTLaJukDxs4gVS1GcOPiiTgysquISHTCntA3ieU9MU
BH4aD/WmBPUNM2ihjQtMoIGAKr8ORdjUiHxp4lYJSAR9NXJeNrqRTCkPW3AqMfU3JzKon4csQuE7
352qWoOcV/5ol9nrQBWMqvazqp1tq6amlIGW6Jzy7H8iStp9dgaZ3VyQjKcJeuQx5ndgDgQxktHV
CwTsGC6ipO5Av/MgwDXpy3dCqY0uwZJRZQAzOh3wlpG+GdLys/HwWjTyZzjtMw9T4lYZZmSJnuNj
3hXmVG9NxutrH4PGTSnXGGvcqYCLvzOHvTN+26m0v3E/6W4rklJlJHCJIX7ZuyGoFC1Z5AyCNsVu
TmvPti/MGhejkcbFCTX248F55IncZw4PeqXqqt9XEIXt4/iTXbOcvTvXt/oxW4Oi3C7SOEgXxXw0
pFI2VTaG6ZVImW6pqroxt7BgsSy10ZTXiAOMB6AxNhcqjYPcViSrCAkHf9s39Qstwl2qIRQwKgHy
DnqBnQIwDUISQBfaNozgdHVgxUxdlE1CAC/YgFfmRLkLmGx/ulmrZNzNOtC5FVTfSJlhTCv3Xnl5
7jujMRaXEU0TvinUdWhh/zN4ggm3JQMogGjZlO1as0unbS4LFCPyM2NkkShtN1W29U7qRxtgcBOF
ne45FOu+BLNQFKEY94Tsjwn6KXyPEUZ0y6LalL84Zmqv0OrMj1lXu7AJ/tvxnQcQFHez6JLegW+G
19By/vBvWbxOxrJcVXVrsETDoGN6/DeQMlP70q27Uj7Ps+iIY9mmd4jl2qUM25YSVquLn0JXvhjf
un9ILeNwvasvpEe9Q07jPMSlwMvO7mC0BQdAchuxQtkIX3t/jKa5DYVdrycaUSIz77bRAJbMSiRr
/Z16711kK5N+dWJsF5NmcmehgQnNLxofxjzbR70ABO8ze7Twe15vTtO1qf5THk0KQmajsjTu4rJy
UJOe7lZLDj2xs3TeqBzvWi6sVZC3nq2JDWTfdFPqyTyq7fynA9KLbsTbb30zwNCB/6so4F0ug7hz
KJj9P9uNMxnPMLPGhqhMQV66R9dCj0hAD7EXeZ9XYqFzFoAwcWDIceCQzz5K059O7gwmOSYxffvf
PvP8TUQ01najVxRu0ePMxZxdKXktcaYCCFD6Yo/CR4LCT1t0dfYfMPGCEs8bI1D5XDlufjagnUgY
+YomYXhFKAddOeTH3cd8OeGzalEVWZ5jzvDCuIyd2kWy+dm55LnowOPCkxNElnB7Y+Q/GK7se8Yl
6L5jujqe7rA/Ol6j+FhI7it+Zhbl9ZFqIpsjc11doNPffWhdOn9oNfHspGgTKJrY831tQgLztGgs
ny63QzUNuwL5RhVcNaDbW4x9a9wQauHTtAWjMFiJaVMrHbbCAvHRTDgDVlynaVvrBASuh1SX6Pvb
2zLf7xX3U+Zk7DS8VitXPYwTVOtkQh2l+Ey/qGqdWfUjAWq6sgPR8x+d/tBgPF3QdLi9yTTbHr9K
6q8RNclX7+7SGx87KlWvEd3+37xjtszcgMNo60/y4VHW20/ZC/+KLncgzpnjU3yMYjKvwuAEOHOn
FYzOVV22Xnp9bEjWUdp53t6mglf5CdX2G2Ncf31doLpdWm2zp7MzlAj7y91VWAfyV7Vo4rVyEGkx
dwUAT5OPUO1S/uNX1Aee3zoA42q/TmRaq6QEUOLt7xj8o+cRyNjMF2JqnJ7MfBhD9ZH930qx5sm0
yew8jCyhnG+JHjkPwImKriytfnUtExQHDo8PoJ/I6Qohg+A0nQ91HFLdBBYazJYTOtryCsJydjWb
TLkD/rFnUxDxH/Jj1ofEWyG6lz+OHHOuWHb6t2MSNYtVyOOvY3qZR+od/A9FeYnuRycyYvGA0AsS
VuYGOyKbchJRi+B/RrbPXkqouSfweK7f/6K6c1L6lFO/Lx6oWZzQktagfJCa1Ht3h4J7NNL6PZWy
Fe2/zDzwd6MTtUXBQlbGIl9ujMsfdkFCqKXQIt3/e/ARFNdLzwfz8M18nCxt7ASRWJfxfFMbOCQ4
r71Ry1eJsqKVRaTa1lp3dErfK/X8oBfEMWWg6UCbh5kBnAv9ofKrDLHSVNVjjkmHR24TzrBZ0aSG
HzpOFPnitJsI0LgkR/w4uiQ2rxZ+aRv91yZ+4/8746I5dbG/zfCqrScbO4nG9QLq5Mg+jQnu238Q
6171eyaU+dtlc/D+iwAQY7gJomBPWsJReWfAJGi5B6ZVqLP6JDbnfBpXvUh/YPoVqCZDSWoJRDI/
HW3lEsI/x/tMZwx0ymxKt8+X4nTwtgXzUpeHlI2LYIETm6pLS1dLG2/aQVR40R9cyUkggJZimxKx
Ca67zfBg+rv/HN5yYRHyvWLLWm9PRpMefzdzwAwMEEJukmcdR6R2JSTFR74RyByx861pWo2W8epr
HOol18AZ1T4famnkL+MEZMiAhFIgvDjjjgLo71lyDwmupFK9jZPQpL8atWYbOOdifmAh14Jy35Lt
pObLDRqvrIIMiZJJ4SU+HWsoDMpVqGjdrELlcsrMH09jyxPR2ywnH/Arr7Z7TcXcUtl117KwFu8Y
6QvqgPsbDFKvCylNYXfMWqSZK0Et/cJnx1q+u0QOPp4Wa3SsQ/vBxsAb2VrqyZsZtj35ksoD1RZf
AUOvZMQG3T/p95J1cGlTc4cbaZb6w3b+ndaw0lu7bJuB7tCqK1UBvejXsMVFG0A2pkPDYVbSl9H4
OF2hHrayCmLNsV3I3toJLO4tUJ9VXAPXGh+vp7jov6ingBMNQauy/U9qyjKCFTnSddwr8VOqHisH
BMqZKj1vuo00oyIuaACwpk4L3Pb1bHYYXPtS1xHnXXP85l6Mi92EpFy+j53gYze4i+naZpM8gk6V
UkpfTJktT4leSbYU8andO265KeNpGIR/eymWE3kkdWULOWS8/2QTYXUhgZ6DAqZhkl4G+V90E9Pl
fD+9KilxFMIrC4pUPkUZz4T2hYzk7db53E7atVgPPTmPpIdh9USL3sqEp9sdkxjLNAPzHBO5eyY2
DKeB7NvJKiQRBzb3zxMHxRXRdpa9rUuHOsIs0c8azcpyVL7Yy8nV6ePX2tx5Op8MqBsrk87bNOyw
buroF0aVq+Le2MRbSPLLhTbRq9Y4DgfvExS+bG/Q0/ml0cJrXEpuk/z3ehdxFkeWNRdgIQpWtr2c
3c/sklXAp+HuGb6J1BE938ehZiu1ne+CDK1pCGUni8YuRMsOkHSgcMT3SwLSmvja4dIZvG0Me781
+PcH7qJzC/adckcffU3AFfn4h1J9XzCa857T4PndJ5NAokzyst4jezDeOQIz121LlALvR36fjout
XBt8H3TDcuEwIq47ZcQhnpAoBI2BKrtSmkbZG8oRZMNoDlq3X6XivHr2rn4Jg4immg8ifU4QhfAr
pNGIrGbQxnGzrdpv7TjQYfLPzoA7oMpTReXYLk0lIKHMmAMw8Cg+UGb4TUrLmKmNFjov29HtpYFr
0n67Wtv8xq2YwCT0RVFmuGmDaTlV8Xm1TV70EX5pAhEu6RSXS3wwzMRzlxytArneiRqa9H3wXqsQ
eJ1PHUou6hDwrTvSCFWH4Xc+455hzLbOpAzlItxO1cIUVtGPtkql0NnXpD+wtm662TiGxXItMnRV
GJR0zrp0nLC42L9S4CM8PZYZsdlES7B59p9ZVymNqQs8CvUvz8k9fn/KQie5zhc7CfkmYgZLNZX+
6jUhOglUEbC7MwIZ6X3kw2ZTw4UPNnQJAS63VgTbifPlEY6ium3bPgb8Hi+KUkcrAcSGijHtG2X+
OppXwNwKJSr5Mc7/L7hyAqsaXgM+na5tr49BVbfardvtFVF0feZDJ2BYevyyG743FWM7bXU061Va
DwEoY1Qq8EoL+eGwjRogtt6kdP/9ZRE4HolnzAq4yad+9XCDn9ryIdidlLrWo2acG+nasDtkhz1n
fDSasDLJVkxC2hsjWePmNcRsFZZ9f2I76zQWyiymlmO7QvbyrheRU25Allw+2qbndVjMSrqadrCs
VbGlWlYcLwLFSzdzJvjWhaz4ExdN2O4k0rItdi7zDiKv/BKNl6WSIgBKIjOhU6SkRWG9kHSJ8Ss/
2Zi3eGluZtovWyLt/hD/pr5OcnJzYGhzaVh5bKTCCVNMhh19YTeSeu6rSBLrjeml2I8e/lEy8viL
IPGFs/lIzkviJ+Z3sftJ0GHhaiI7cjX2TrZA2Q62xORYEEgFIk+ZRJBPzK2icxmBCalONBcthT9d
YlCxQM7i8rXSOfwM+8f3z620R2FyMfIVGoWE1a1wGzKEzn+giBS35m1UKMtXIMH5sstpYPKZrPzo
X3TGUe3X3RIzfetFwuzTv8ChcRKwTHSRVXSBTSnblNxyGlBODF/0rQhp/fqSEfIi5LKMfgYgsamD
vD5Ut37oFkTO3pkIfkldPca2dQBOgR5lDHb5tp58AsjblvRPM5WlTR7Otw4aN3Vh/vwWFW6+T9g7
MBHI2ugN/uHvUWQ+wGnNi3Ps9UF2xMgzO3jP7ybyjcOlRAzMNYq3IA0kz9/Q66aluoldCLAmft/l
ukupYOfHuAhduxAMxBMsp3SBoOaR1Eb8DORYZkx8rNepMVXfcAFjL1AfFFtRmFdQrEgRM/rPd30c
TcVuY7SEs87xjxsCQChY8q5YvIRofJg+Rrja6JytVc5G166GQLOOcia4IRUvaO9V5GYr7bcaOpx5
Vy9nAMOvT5RS12N2Bb85fGWDsIYGyiavuaGiPzyb5RJsZXHFZQ3Ua5mHb0RPhEwS275nGWf+0/cH
086p1sR04CMqbLfVnrQl6p79vJMz1Pw3TbdDygYEG3cAEeen2Ns+/2Z+QWkAc8eHwp0nmvOL1jWS
AJtNtwXfZdZQMAoRgbP7NIWjx7cXOIEvkwp9AqRb5Ol/jAKb0nonQls0uFufhG/LB2VgfZSEhcu5
oECb5OMrINUEZVIV3mF/5hLfLF4f7CxN3KMNYmcrneVsj03Yxn+h99t50Ke7Z7IIjC7c46IkjVws
dEAe03z0+FtMT7JdWJoYym+I6GERvK6eVd/dGytsdeXy/E81J9cBHExgWYR+2Kk6p3Pbr08uAqc+
rv37rVmc9gQ/EgkEKJc5HEdxO/COxQ+8Mu7cqmHbNVKZvidT5m3FYaYDGhzk8+0du9C6Qql9oUlx
iVgiOf+nVGRlK7iQMSBKEQicTGgVpRvHQ4o2LbPTxKolT2+56p8yRGLmJ51NgOTwwXMc3LuZzwOk
0aZWgq9FhDMYEjXwy7XJtu9GpNvmjTYgg10WHwjIFQMF5uXxXZOD/pJXWqqn5oc3BjeUOAWapX7o
rbu/a1O2zKFlGhmIOpvPqsduFRKGh7u8Mr6oocdc7A16QV0A9elzdUGJhNCljt6uIlQIQcn9ThL8
mslTdgfSelV3VEbtj3zUiun6A4Z+wW3GltbNZIALMA3y4Va+4eFbE/nYhkDZLpC5fFfzGj8ciY31
Sz0i49+XoU35zoacSVVygWqiqzN9QwjBFRQ5JZEs6awMHm/3BsAqAAhifc0vOg8Q0frqfqjsXKFc
4EcadS4DsP/Uh27K72xdA5bmoflnmcQYhFqaiOc4XKQXCDwiofgBgxJnPdzoXGc5nISTBy4PHlaS
YdbvArjzt+n/mDeDMGvMw5KcSkUdRmFjfGnX6shdVz4/mHwZ/+E7CJKp+TAoYKSI7xkf8/LVd5Mk
A9QEt2EThu1BEARn+96RJ+gCDjqFO6gsacvX/b9q58a3M/0Qtgx/Di//H4NaK003f0Lyf7lKLc25
rd4j185qrzCkGuGeoSjXcsEx9+AAW143b9SiYuFg9Hrto6Xw/WFf6/ahIvipERGBXPeuDksvF5UF
Y10Fdg36yYYANmcDBUlBFWWgfUS+9Lj+1sg4l1wRqY5Wil7EUDQN2W1dAOaXeCC0wE50vjl2BzSk
N4Lw+SgW1tgGwZcc11gh19UFSZ5h+1yW3Nh5hCXLKEpExFmNBe02ttaENHRSs3grhohMOX5zvn0/
jFIh2MDMTDRuteKlHIsPcSRQ/Ye4mF+uXexAB9weisJsiNwR1RGv7JcysB4p4/tFnivtRhglvubQ
e6pbiTp41j/NYog4DiintURegUpszLv2o7kivsUv435+kNqYK1AIqphf0rby6jpc3CdYJ8Hzhrwx
e11dnvWpezPDxT34G423Ck1f2WIdCSP/wDH13b6Fn5kTZJpABd6JwPMo4c/mPZS9oEXQYZ2AmuNl
YwvQZo5RLkvBs3l2F+3mLENt2S5Fwj1T0JTuAzAlYXSXm1a0ofxTpqvELFkK4bi34EC1TBTUjrv5
EU6LvPJDhp1XYWC0kndKefMsOkXqXRj3ZazQApnI2BIGVTx7LryPBOOt+l/IYTwqet7lvEN6kgRG
6k31kFJoxUfOtvG0CQyxMXD2b2AJXicbT67xSwMFkRtC3YjI4CYEY8gDJ7RmmkunjGPBe6jm5keW
Cro2XZmvTRzczjC7LfDXaSuPKgQzqKEuG1YpzpC9PxGMPhK7Xx0/NlmXZGYQEvOh3NbSje+eGoEn
SJnJeZqiMsuxG5hTm/6tu9yOX8Ys1+9fxfSRTYzBNT//b/PHzjw1pxcUNnbRyRxJxx08cVGdagF1
SrtxgAkd+XoB/mqnBDTv4YExh6HYZLHPByXt8M3HJmkPTPUVM9JjVUe/pwQDQFaPFPVKcZfOVdXo
Jsjm8748+PIgKutr64MTZc/8QuSzBxVKKeCVZ4/j65cZnEPDmsqENIOSqoq58gSRy8y9lQt4JEVu
7cVrZYXEZIX72sLZSINPtzxizN6eKGfuQwdN0uQEiD25K02/dUSdErMrT1E/ORADjkAURLlHDpoc
g7eNnV+/I7aoEJdm9cuovT1sz/oR4sR7Qw76ttlfx/3krGYWAa6cXXrnaonNY2HTbBPR5Qi6MwmL
869irJZsv39UjKNZdZMa3zaftpW7i0ruPTVYMIpWU3yYJMIJ6UldA8oXspIXypGNUdX4FZIhXtXs
kzqqpn6YE163mEaWzWGhbo/9C6O4EBpI2+mqGEDRRf5W1fXleUKLjDp8MEhkJfhJ7vpZKCC7CiLx
8HqWAJFVbV5QaI2UXpptgb9TpDNBh8E9s93IvLsGcjhIxB/EDr4KBkxNegNE+JCx/Ww2pTXLv7A3
3NZugbpPfI2rp5OA9lw/GTwLUllTs1+PdEiJBFgLJWPzvJqSVHMCYqwN35OnYXWBIL0Apm0LNSDu
Ve50kS7EYYkAbFcf/Zgz2xv7qBBAMg5fWPVmHRLmobTAuEkpwQ7Ni0S4bq4cr7oTPUTqaUyW7rZU
RouEhs0eJn3HDhb2zn7Q1BGeP4SmT8Dg4qjYmyNT361D6+STk7DKS8532ASwzvXRtSk/ttYmlQyT
dingtu21mSXiJj5TNNFKM3TNSTbKp1mQGamBBLPH72PEFcTbFEXemAsmenIB89Whx0V2a79xF23a
ois4tccw1IJNTBpx7XbsrFGDBT3SQZbzA/x6uTUXrJTVaJ31nqbJZhhcgQzBMdxggrQ3qUYRX0q3
fjIuepBY2Js+L6r7IgVk/FvdXjIbjoUl1NnFackw3q+vZZGbI9lzLI72iBKmQE1VCX7TCwA2giNp
rSaSxlOOPR61g0/IC/BALh+exybqiiBHVRbWlHWU3YoMtL/jQIEe9vtlxntWmjiwiAY6ZVEVUpXy
ALCbfAJGj7IHoYrIRq3ba7ujA98XoXv46b9CQoSDH5fJ6qTlahltBa/dCpjG+fAd3voavpAxYEAn
C5SsjjaQHuDZToRQhSktGypAl2uhRByjSYYqhaGWJvZj27KKVdSiz0R7PvohL8NtpBeZgp6TeY4r
SyY9zN2JlNHXzep4i6AMfKETsytckxLqiCH0BNkXc4GFK9tI96SQJDZ1KA/qK/CWtHA4DaaN2rOh
pYytUXCSo00xiBWMqieHLA8VeFlb8tVDM5+oqolxh+7GGMErsejXe/MuOJtK4H8ljU3MowDTAZ/D
Dj12jm/BIkWxZ6NLTYa8wtAom4tewiSVttVglmO+1kTL7LkU9aSKTRfoHFGLpeDU0Dz/ui1CYLZe
seQYSeCTtpCGsDgUIH4gjmDFR+MDhKeP2daQPs7Rgc70lUkGu6cvf9qqL9yuL/2IcMiYpbRvqy2E
By9PlR8MGvMlGmPFCWXkvie3++IaPLtTKiBp+AOIJkWsXo3JZ9GQ1XnmT5h/YQPMcYhLhVNV900J
afe1FzmOLMNjlJr58j9fWJg1PxsYyic+iDc48Sl0wdYc6YkqY0y+DTIosMeKEtEBdxSnSMwdmjai
ELbGDFOXQ9mfD0M6a69BNoaUI2kJa6XcZIrSAWhb4MmJd3g8wKKZfZIZw3VMTAVvBopucHgF6qGo
Nirf2gXL/8J7QTx68g8f6kMOlPnRW1LY/q8bY/VIrgAcIYIqTCLta9OEjnlYB/Jo+NoFyUhwUlDY
F4n4FeF6FlHMxQqVZrn3Ok4tHtAUpaUqbzoO1J0BMkQHo1M4xJn128ZJTf8RpsY1zP8YvdJ512kd
L33ux0Ik+d5tSz6es5k1o6BewhYDemEW6mfV5tbjvtIFAJlIZkOm9eykgmqAlZh4dA7LlwWY8/zw
DgkBhWT6Zf45UjpPRUcG+6e+Js4Z5q4nQ6w4D+GaJTLlD38gF8K41crp+MaFQ7tMb83FxuZmugyJ
RkTSIxumbXGZhzeBXXfJWLCCo6hDstv6eebkafKeiZSFpa8Pp94C9MA4oBzRx6VXVsAqSIyKf5Jk
Np+BlOsDMofkP15H5rzNwFzb3TuwKoll9IvA2W95DeEyfYm7mHSCznoRAOg8xHAssi97e3GTJccv
CTnXjTzjbyU9mdK8wcwiXVKjuLDmJLn1GcXEhkpGqmXv9hDtoOlWe2WWlgHVFTX5wTYJGf9rpI21
f6Rmy9AK4ClN5LSer3ZyoSc2mzDIJl4rjKI3v3CgiMrIOml09oZMloBvEBOaE1k2Pcv/BRc8e11a
/C8kKj3JgS+N9CuTLnnkFxiyLHya1zF0jPkClPtx7B60yj5rIi8pXUjt20R8rLnDSys/SCxHfZpH
d7BAPkJvwAzwXNo8C9MHz/lUwnAENkFF7widB29XX8V2KXGzDq/fIHF8dN9RFfCM8hCC3u1zKpG2
ZbUVWpermwvgzCeH5PEk3HhTrns3vA0XKG13qyW/WiwXMrXBb/b0EyajcET/SAh+Kx6VUOiUV08v
MOzOqueYF4EUFXgdBPRNgnvSM0DzY0XJmQvcFI+Bqru1MF53DQ/ApPYgdscq4xKm+KAK0/PUFmBs
y1viw0BHff7QCvOPiZd19FjF26WvNGDhhIJSUvpKvcl/nwekwKU2DUQCiqg22GR5yoTaWsYPIpvR
pteXdzjqAuAriLGB32Kg2BdodcCn/4vhjPjENhZpj+8wiNJbwFTFE9M29NC9asvfU+nvfwuSDZKF
wYVySA+BqqjgnTBX6z8BpvvM83eJ9VUsy+NwqnssuuB7avqOhOmwmwit4KPme3jWgijcqcFOLyxw
mbbVK8uryycEvSGo3zdhzEdB+2ruQt6BjFEyw7BS8A7PnQEVOzizllrzR00axqA2zxzyCehhxrBG
SGATD3xJuQQ0FmsB8ZdzWFiad0V5wWEkDOjMGk5bjh10PHqoKJAOynYbpSMgvbnFs24YyJV54tW/
2w46RxTJnBAQ7rXHgEaVmul0t30xgad0O7MV1fTHCZSiKiBemBVYssuYk9lWzbwHxNXWfKEVicHv
E6YltSBcv4g7SYbpVPE6/ayzwqka+w3u/RPbHWF/1DPkYY39jJeQZ5MnUA65PVH7cqhiykXDmQWG
ofBq2zvY2UG1bko+YU72QHP/7DubigtPLXc9xuhnHdSXEOaAPTMxBqHezGdPHREYUbApUgiIcq4Q
7crANeRvGiMa3jVlWUQnhvgs1Hb9NZIr3QR+VXpMnBfqgC+FGFTZnsFir4JGLABwjJ2e7Cs4Co52
ttufSN4j6vl5C2MCi4rsvQgLp0j9hloso6hCbUSUXQvFmMQ1vqmNRNH1T+SCBzwWtWrVCgVye8Pm
VxH3dMZnw7bRrAuewpduHg9StHqcIq+FLEG6oTcxpgunlA/iBtlNAdwz1D9E/M0raJbJgmwjKiY4
jdf0QdvBC/KJ7expnwEHy03njlZFW3wnYYivCAuY6fXOPGqdSu4jrO+xcjOBxFuFmgck31Ql0rfE
wBg8BoE5UQgqKuIFhi+C5QUh4MwexOMGISBOEv3ebg9xyTvcR/77Npt9A6osfW1RMpZ8OpSxyFY7
8saNBk8tnH5m66zbdKMyoN2NeIFVM6Mj3XEOPvg8dW1iWowT69nxgDSkSAl9j3GpWQTpTCUHkwbf
W5A6a/mTF9aCPJK/t9DdgJYqdU89PQ+tHfFAbAsEuY24zfzSuwq+/JVj/6QW8VAGHhOFErz49zF+
KfKVtr1jdf3FxgsWvpNeTeuwKrbQ/KrpyqEhVcrqf0mBzC3PPAAGzKQh1kPShrr8BZ3aWpBTjofc
l8Z+gf4uKgjNEz3XGmHWf+B8FbVKT6UZAGU2CwBYq52mxCJW/5qm9NCUV7RKJKfP7kE8DrxAO93d
Tv+mqJcCQFlFOoE8QN8KumQeLWPaaGbK934eruXG5EOkZDFGOnj/SuMxUANuyZKg8CVEuZLrKtL2
s5jXC1dnRxErGw+GJqu2rD2VV8TnAPOZlnXbDufQaFiWB4P8s9YP7qp6K7ulzrR05JN9KTfHdrvd
arY1UCHUOcb1FnrlEozYGt6EGg9WqERrp1YY3NDccRTA51GZ7r4fLbfSayYHGchjt5sP2xNY32HU
vq2+o8GuuW6v3U5HPxEU8mmyIrRUhGJin9yjcjN1JdPfA8Byema5o7MwMqkOT3N6iee6Lik21kd4
/57orLYUMZk7XlL8KQ1oVqHxeRfnamkAvA1oigzyDA8gQ+QlR5QGkNPfOUoKy+UbMcrVZNCe2Tge
6rcaIKZc91tFwfo0XRmxLIIg8lW6+HR3iCpNxlTg3mL6gJbmCpTZTQ8wwbjIdWHHaUUrepvPtA/W
UQjoIytuAv9pRplpUaLYtb5m4cNj+Yo7DqXBS486GDYmyAi/kJ9BB93SNht+G/jAqc8GUVJk0p1T
0ZB7SjtRjEKbRHoF/+tlCTx3xzjHSvNIOWqKhcKHqW7JJ7lki9btFKF1znceKL/M5pipmFUvISEc
Y23nGxBKWJ7CcHr4DJ1kvcv5SLp9HHII0W+d5eyaXhL3RSIV8VxbVlsUaakud1w/lt243C96gwwm
WSJ2ej998wxXID0mycAFOgtuUn88y22ZcIw0eCLZQiWahL5cN6Xpyh4F8MqjF7hDXVys2OkSh/I1
9pV4FRNdK7ocbRIr78l/ztlVqRFlO4Sp9iJHPa8ssG9SsGTsFTCfc5OCpGgMAmnh+KDzcz1ixR5V
2F0Th5DUiS2ipcdL4MCbUOjpEIj45EVLsk6QKFFwXKJIAiQItlcntqWw1cMYEyqanReQB4V6yw7J
R5ohFKVD6WuVEbgZwm0XGNGnMqBNj9audyc0BtifZ9DG8p2fHOXq53eZSyipzXuIhbUmBk01YzQO
P6vBugIS9YFXe3MAtxmmX5VC5yLN1Fm8WB4YwsIma8lRyNVkvKSqzyJWxnZ/YJioq6nIrzLMyew3
1ObJLFLt7cNcigeDxFebaKv4yohS1W+sG3EZQkVWRo3WRWdFabOLUsNkvG6Cbxg2RRc2THuwxFHK
NII5bs7/LIY9SBZATfAt+Mq3FPJ2ymbJdF1PWT979HltgXGebczXZ5VA07nn1vuYD99pjPhvwdcf
ti5PYaIJA5+5NYbVm1/N5Xt62PfSZmH9qNKfJvGCjH7jstynytaTG8PhjwlwMaNlTqoxkXGXvKtX
4DG0fo8OJYjjRgGChPLoIvGVtsHF1yp8T04/UEh6K8yRCgqGkoZgiE6g4gWuPkDZs0wqxhvr6We8
iqsXS0iKiKnrIztu94f2DCEiCG+2r1qBWi//WDemRq9EqxhdjaftMx3IUImRjTiR0ZWixT0OhdUW
maU699UJ8RBKSf2Sx6M4eMQvrtCiynrX53Bcxj32Hayvt9Wt2yme4b4r1D0Ab0Z4rfTC2FwkSNtd
Phs1YEKn7v8MgZIB0iVtz9ofQj1aiHJbnqHddQtNCqzV7NoyQdG3TiiFnh3zL5lBt4ADvB87GOYz
NHQYVzI1U3yPPPQG1SBZNISy+41xYE9B2FNRwn8yWkpvtikI4yP9qRTH3AT3PPi5GqOPc3OQvXL7
Ug9UPhFaNyOVXedclvCUawXjUqUPi0f69d6JEzIWq4ops6wAcTV0Y0Irm6qjrK8x3JifMw9vWCRY
tcZen89HHhCFg/pRLvBJF0m+MxaLcua1+iIENuKSsTAkgdFIyXW50eWz6dMW1Aoxe7MS9BcBOShx
a6MxvYxu1dXd2ubWVy5gzzk6GJbw8CQUEpSot/4IIe4EPZBubRxn4Cj5GOv08c+R/dLjX5Q4q+1R
6KUSREqOWVMwSBowXk7C1O/mCqqxKLSR6JzPaJFvNLGbkf3hliAikMjSoJMsEd62smpmNpsLimku
jO6tD28+FPfQHr9P/Yljk3KIx4aM4BqfnddDQtDKXhHP2HOsxUJUgXZDWJPvBfK8sxoxA9vgrFWw
+1HBcns091KUOzDNA3UPzsPbTmzwcgKbqi+/MvtZytL03rQ2ifmsZtAlRFHs71zkThB7olJfDUJ8
qKvgC4/rQPrcNGdzY/vHdRIJuh23VB0Xp6Rfk7Z4PuO3fj9mo/yvlQ1E37ux4JOJ6qXwnIC9Lj1b
LpyQp3sMAE1l4X7NOutcFESFl/ToWSBjRp7jcNVyIe5X+p2/0wePcn5l99gGy6QO4RwAtkHmumE1
hZtFNmSQRGE5Y0fkRH5ej2uZIkDHTlCryUsj/mX9a7HJIN0dnE+YN0iZT91qICTJsCrrFc2qOoft
svzz2U5Dy2I7pvoJvsF794Q3m1l2jWKHT7nOa4Lvky01u0qwvhabrp4/aAYHvFNeGDCwvC2uTrsq
1N0iGwy5RDkhF1KqeHxGPsRA6K2nq3N3QsNAYVUyxv6sgXAItWS6bFUYgfsdlPltdDG5AhT0q6AP
MHl9mwWaT9cHD46eLFGJeqqrFOSS8gPTJTmjF9pkHAP0j22ox7G8E2+t8J/sdzKtbwNGMgkPLEpZ
qWxQEH1HFSNnJskdw+y9PIcVtuCkYMW6S8lPe5dz/iZuMHvyGznENpTbDhHc9GsnCvrSkg0afMNP
M51hQoakassowze8fShBrFvL/7rHAfoWPdsDdUBISJufYy3ONl/JQ48/vpPMFSqLwHIYKUocP95E
0Pz/OGKKcG+QgziEB9aUoIzI7MYpycgrpcrRpSreQJOsRnjBDx524TflN3e8gcg63PgC/OSly1GN
TkLYi1iauFkjx+06Nrt3Cqt6SZUGdxl9ZfaiAwh0qxHe9erAgArPdSxSAqNC5N5caSDCaL/8gD/r
NCdWIgaEEjbXhjUySpS/TozUyCo5NleWa1xt/u55zJZev+BK6qWkBjesJ0FbXUFNGgc4sajvXIQ6
vrm0clBgV08GFlSYEETPVePHD1diOi6HS4x/DNt1sJNgI2y+0se4ReDm56xg0pnolEjF2VqyKe1S
t9liql3YE1iRg+K7g9r9EVrD7p42hLvgXDWovs9bOYq4e7oHFgjxB1iKQzPqnD5SKNmfhe83Vq36
8CZHlrt5nwQy8EcDdvbok8yWEYyI+/D134/si/1EuFGj9oi020frIS+ZjfanhQGRmS4+lRMpwYyD
wQHziTOxRbSiNNWdZ1bBKzWOJBm/87dVjWgzDmeYH6CGqAQOd9o9gK+gA/w3UBhj70CRjpGc0ROn
YTV+Ux/27MoByrALeIGw/Yfkwr+RA6mZx/QK/6tXi4Dxg3OnYQ3lINObgpgZK9IuR40149uzA02d
7FkQYRgRsTqXbisH4FPUjEUoY/kFYo1RU7uKSM3cRWy7M+fgTM7pshpZeLamfhKajXKYNwC7F2gB
QHxCzG7S4BgBYCciAy3MQOwCZe9ggHiR7XGAwEMKa6B8Igl3UjPyCbtgM2gVniUBxvepALXh8ISR
8cn3AMl6jKAezsg+lvOfjv1orYQXs7ol67HFUAsXc6e3ZIRntv/MQbDQA2m8aTLPufpRxtdsrxUg
qmhoePtQUjqnV+L7MyZtcKcR4JbPlUXj/lSN6bl/RklbV3skwc4vJMqbaUrOZOFq3HnSI557rTvq
F0rcfWPKnUnDy+1gja2FGMYLcjvfpMPtU708PTH+xYURC4Do0ZxJmoNDpSl9AnEK/HumkuZJOxya
2+11oZcAdWwFj0eNG2X+0aYfnzH+RfDXvU7VOvycIUOqN3a95kpB9Xl/4ImWCW0jJTqw7uKZ/Bgj
jdEttZNBuf57slXZmIZcvRU4OiuhEhV+LwIru1M/XhiHbabMnmPjGiYzJ1FBITVrHUk6rJl4m92J
CZBd+3QBwwwL68RJC5kSHcaVmGoCo1B4nWBhmYHya9L8C7C+oQ1ExfGU2GtgYtszrLrzduN5C71Z
VaS+r8Lz2WxS3Kky8bz2qLpyuuZFcsdbFtejoQsPf7tZ4UuVLjNNuO4To3DZ/hJ/njA+AcGKkHn3
IJUIrwSymj1w32bFjm7p1ze5FY3/Rtv+8pOo3Wp9GsHIjGSGbiF98Noobn3PFTw+sRV/F7Nv/M9y
1itBbhpbgbIG3gKwjRoSjnhjXnQ7X7vRyP4mfUInk22ps/gg8paycK7FJZRLglnblAQSDGrZVd3q
pxmBYAbVKLRMIzoL/PtNHJEyjPdWilwj5Gg72jsnqIHLH6H/0sjSbVbvxt4VtfwtBAPOjogVUwff
UemDqjuqqEC4I4v/X7ghm0CA7yNfPVCW63iuHHe68hc6lTGZhY//zORm1cOLUzPmXJsYXuV98TZN
DuuWdbOclw75grGtCzzqduXQ5qiyDQNgo7chRaWaTdPx0vWDtj8irzI4s/Tq58IEJIK8AJZ4EJxz
wuXfH0jKObATOOZDvu3YAyI9P5j2K3QOrH8Ez/39a7RMWIH9RGX83yIFP9hwIn1se4Cc83tXC1Rs
jvToAjXWriRKjEAQ1ZkVEKTnjV8L4WRh0Wz8cmVMOBzKZfZvY9FY0rkhKkksmwJQZ4a/+tzVsQi9
7CVHmFW0T6I9sRH7z6FythWzme1Cupay/kitbvV6z9/AEi7IbgdH3jg7MSuebRbSTTVNVdoXgyGn
aGAcxvdJXtPe4WDzIoINEQhBUBkp4bhucbOxKvQPI/CPaB3ItIl6CFFx0ELo79ulQsHQYxyAvCU+
cMYLzTFixOaWxVgE5FCHGxDaFhgZ7Vh6YzpFPpmQtPlNrCyr5J5LH0VBFUw8w/RyStmLvgJsZar1
Rfd/hghG22jDJdJuh4dnxtbp2/XvCdNXyX6B10UwzoxlHx3iNG+m8MMAH6Vcj/PeEd7tFChrBTKt
FSza2/edRwlegY+yW3zOFBsb8NfV2EBi8b5hB6xJaFKhocSFwl8i6iPyEojQr9ctYzVWh6RuHtUh
QNVq+gl/i23l3qDrXHZartAQ2z6oK49ki6Gleo15RjR+oHGcTbvYpEFlV669gdL0P/kPub0oZi9b
bcDFffBXBE66KPGieLuLmFvmNa/6V7X03vS5WEncvjngcBOyFkznTe66yQaIJvLqsLXw8M9LhcRV
Z65cyz5EXkwJbgAul4s6TI0z9T5sv2RMwkesgAIEJ/dRhil4dayDXKUr6O4WcZFx0Yl7cO2VeMHv
zUJCW8YDkP07dfByRusAq9GVRXlMlhSX/qB2KwmatKch60fzW8vkUM3kE7ilSdn8Z68wZh9MVQaC
GeMeN5fbQ+oaWPF67vmB6/QJz6e0UGdBJoaEwqGpZlJtdoSh+BzcX4mRRiFj/mCJaiGumc2PZ6ft
N8IaGT5Wby+FeDTXIzwB4CnI27+XEphfh+yWuV6SWt/0zS8ULVgE7JiHlgGFwJoSkMsvzjg3M2Ri
AwsTWUpgzo8aRmKOzuITpsO21LbI3js9zEjpGHpCr4CXidVj9sSvEw0m9rmYAjXkayFT5ixDEms5
Gz3yxHb39gbIozaKFcksrb4q3GW8q18x2Wv8MLhMgQs8tgPR3uV/8lktttjMtQq9MGH0s6GPnaJw
fUG3MVG82VaVf7xglKc0p3KSlBxBgjxgLHAwlWw5jQXHoPJdLkgTogXlgmLj1n2XRMQkpXGbsxDu
MZ8q/ItBGNr08nvz+lD/SDYotJxWWTWuRZ8TyDFZc8hxlPBlXNJ36oiefp6DNgi/YmthUSqey+Us
DVBa90UzQ4KzV1VUvHesC8s3bh8ZighK5BJd9nbiet2UgGnymBmJQ3ehJhpIw86MJsSdyNYkxTpr
BXiUyUl1VuaxqYgOr9AjcyBqnp5D5btFw91yLItc8VNCfDcPeKeQZWv+enxv3UaGwcVdKKTAyAiP
BxUzt9+07ZeelLI28v0LxE9/13m1ntmck+rM12SSTgxIIhlu+YH+tG92Bl1BnJFRL7wWrQiQmT6g
ZBzUNVr6/O1KveohkbhgcjHdF/dY1NmtesGF1/WtqK9uCuXYiPEC5tvO15lcZjeDEFw4mzNT3zGY
4Ebv3dun8MDpSpDt08NdG7r1yaUMtOh9NQUMwFUmRVVUUmDbcCMiqX/ag7holZt59j9FgltWr353
ENu9jNRchYExuW07M58ZFNwio3M7HHMDngK39IT03VMvUsqln1McQzuuRTHB3wpcsr30JBdfZldv
7Lwj4sU/tYF7Q24J3OdJj/KJCyEi3B4vSYShMsyz1XmyVslm/2Rkf17rHQ5ryTOywmbX5RZTdn4f
ZrGZR0NtbGoL7VB9JoN2AINLfNd37PLAwCgPiDvWeJxnYJAjk7WVgjPGSdzzWTXyrpQf9wNwpedK
/DOEAHmRI4sjcn/eX2uXLPGBdcIWCkicdj4tcDHbN0PbdMgId82mVJ+gudHroTKDjFq/2fVfbIo+
7QfVntcDi5SZsr4Ax/S9uuPp2kMmDitTZbWl/kSMvXOShjUbnev9pZt5jGXYtBANE3KHWIb2DZvX
pqw1ftboyDIylqU3G9WJN67R3Il8nk06dPkOwQWpx2sJH/3LcO8OwBjQNhfxUTI6oSfOrv+HiR4y
ubo1Y8nippQfsJjTMrlyqIQlYA0Be0zZ26XqKcUSPupLayiqESo/38Nf/AkzOxlxXyg8ggZOOtFO
zAsNbZ//09a1br3mSE9vJAj5kNZGLukzWDGqbcKd+oeX7Se7TWFCrJuXpXb4+N2OVOClfTSFDeCp
E8SBuaH+VoczZyxWmu6IF9D3tQl1xbUrn6qEmM4Z6vCLW4e6No+TjojWqBg0sJV4I0ROacFJigva
LHnOwMAtfMmBcGIiQOd9u2inqI1zDZDaT8P+1/4/7gp0k0ktBMB6nnoCiQN8sx49/KTz7LxYadgQ
lIPGRZMH0sYrUh4pOqqWFzmK3WgOWVvY2AJnbzaCm6bwIcKU7MQaqUQMicHwq+Mdgd6Aw7saK93k
RH+9IECVAFuDnbmifYDjXWV38uS6vHlTRdMziRs7PQAuv50sXairAFnuLQq6CEeVpuLTeu45j7+u
oKDobNPdQV3meLBT9J9/wvKMxrRGS6ir1ueW5SrntLPU+OB2uIzsTnkhSJePV1vGoxct2fbrdyn2
AD9Vgpe0Evs64uDbA6FbHjMRI6BoUCUA3ktnUA52fAvtfZf8td/cjIA+XmxAerlhGAJTvYxxtRhS
qf57jMlhIVp16cde7TWxGYsy/gr2DAPfm4Zg+mw6ApIaUVAZwJ/UEv5Thj8MVh3+JyIV7NUKbv1W
RfXbfyptPdbGfg5Pv7HRf1xAwnD1iMSbj1czEOqZqJI1xiFbcJB3tLzxWicZmxL0GKZeQVcnRrHt
br6eHDvc3vS0THDILoqowSuOqizqKFMzYd7Rb+INOaj02fkL0Ry1llG0dwCnwtnpQYJ52r3jb5eN
eDgqwo+2E3UEMHoGXcn80mSIlKQID4EbXLQ2GDTQqbmZZagy2aaQegXMINB637yFqQfyoHJTWO5p
RyDJue15u5PZp0I1JaCL6tvWw4k6Ijp0E3VIq8VDWA0wHQymjQt/kdqiITtkz1Lu9Mi/XWBCzdyi
a5j+45Nd5wTS+tvPUXdytEVCslLkMXJ32LNgcP95Z1hpfDHaTbitT3eJfVwMWQS3r41a9snX9uns
PGI/9kt6GFFdyJm0o8IL+koKhTGkecQWk/4ig6ICHAWR6JBwUFGZ7fk299994ClrxIr6At1voU5p
1f+R9/+s3N22rUG1BjhezSfIkn7Fs9796DjdbLiJ6Ax4fseSn9Xk9KbxQDzk2o8oY1TDMqmvNCXo
4VhkztgUc8aL/v6pCy4MP84eG5pGuZ73TpmDr3FwMEajqOVwK+heFQTFsHnBpQkFrw84d3vVNC/x
u8XSMOTfLZcO7+Gh4HaAEtZtwJEDdD0SyU2tWExG+YXdry3c8wOcFRwEjIPIUCNdrxqrtC/DKWGS
mSJp+AI4E6cvPEgP41BU0m9d6UXTy1JyG4NhK+kgCfOD5CZAG3HBzMPzifq+JDhKvtvqND66Axqn
/NfZ4cKZxi9s653qAq5IF6M5oGFbrj7uLIRxmqws1RBU3h+2QcFQ75jFuN8mNNPLXw1QlNcG48U7
ylHvQEOpS4vTQFs2gJ5lImbDbKcWoAcltgWj68wpr8PpuRi57no1A27Q8eledfNhyxnHWEGAi6+C
1cm0lSTUxZ47JLk5gjyfy6+lslgKrCLbUF9WY5KftFPaQlPcHJ0jjxSeJIB2l8G+sUsqKgRZLOG5
R2d+TCKVSLatQ3uwc+NtB5Zh1IbcsFszycKhvu1R3VFnwVOII6sKGHrNe4lDJcu/Z2pdaku0r215
xQm+ZLKb4q1vyFlLEnMGHKAYfoBd8B23sVMnHnU4UOggCzqduQTDoyE6XWZYwR8wg+U+yy066AJ1
YSNiR1ypTrycQtsCASUKwLK9FBMjZ3NnFZPLQHXC/SYqA5a7YCyteMEWC7PsZ2KsSpCGOvliYcnK
6O80L1+boNDt91wGzDQIpozYGB0Mk/aueOD9E/AhoaU3ZzdR8j2B7qafWyf3M0bHtNpxLqB2qjVD
ZL83kctHog5rtOy4RXS9gvrcCXnvO7FoKK+Ayd+MPwzMxgrv7y7uSme/KhamxnEx1mOJS5JtS9wE
616WQW4WI9eUkSv+FF3yGeC3CmXXk7/dmVSiVCl4L6KF7XvCKfUJvA5Mchh4xds5Gnc7/zejDDvk
QAGGrJZ0dCiYtlLSxiKr8jNawRmBu+RksSRFh8tShjsA0Nk3bf0lT7m/4LUSmMd1BE0yuCXjw+20
Yh7dNEFIhUlCAuk+c0PK3x2N9fwvjA/rqaHBarv7kx/553g/k2tWpRMN+fYG2AdzA0Qqhn8Y5OU9
oy1RXqF2f1HVBj7eVy2mHIFDnM9MUHJWWtwmEdbf/tg3pehXWuuwrvL07q64l9DwAefWLEvQoL/n
4JuvkmCg7a/5qg4bMBRzbpBEhXea2M1v4va7ezUuovf/Qs3eXUpcVMEIzo2qmypdiNqKtH3Pk2Pj
UJbtnDLMC7Gs4/pEJBpPXG4T61ZTY4BMRJadbM889N5Mu/AgURmYX3Rs76FveTzi1gYZ4CVigRUt
3qokt3gl4IvtVCb4pbiguf8OeuIwEHlWcwpFkxqgtRUmPwNI2JjxLx4aiR5IDyZLhBVOwTLXsAVQ
xQAqGHO+ps0sIoyzNfCazK1CboGT84Gl5kBx5T1yASZdbUxZnlQLc9XPG3fT+O01q15JY31v8X2X
py6iptX/Cq9rK9mlFKiL9VeQOncxbGVTVYAVWsa+59wo1Xdlk8s/l1w2gtg2J98ZEbQ/fru+WkRK
1cYFqlGkapb7LOiO+OAjgEfLu8Qul/jmcRA5T001n8azOhxcqT0PmRTUm5hyzNDQzSgEZaN2WJd9
Gg2VTEqRhqfVmcx+WfgHyoJU5oxR/73EXskXj0jGqP2kKc68u6zVXapuQeTWGq4kOFoVM/gotkl4
NmwwXKNblZuNx8as4TavUtC0lCvraKF7U+s6grjdPoejBio7s6zji9uSvE4u2WjVGlBer/i11GiG
kKdKo5YV8HCc3DpF93+atq9q8tji6+jeDptx5rAGngZtwPSl72mqq0hPjv/eZt1w4xkLioxPlKG8
R/cOzN0IcG01fdKVCXa3t/Fwz9paThptTWkfNFwYWdZ91k5MPeFovTKf0zrAW01Bz2+Wig8RxFtp
W5goXZ37DbHzPbSPt7RQNLBmT2y9VIQ7OmTjMRPZ0U5aUastaVqHr1B7/HE0cef2CAWMD7MIalnd
jeh1QRCZqQeAys+gyvBUbkuODBe4/84AsgRXLiaOv9Mx0GfIgE/Vc5mPJbfco5QRzVqIP6Tiw6s1
Qe+kVSjoXvlPkeJQsDJeX5afHfHboPxqp6aMHm7+9o0S4skXWO1iU8VX04GG9PKezUHPOIDev3y6
WqZKNLipL51XoVzPYMpeTEvq7IDoNeYP7C2GfmC0IiuT80m0Vs0ZVPcepF4wiUSfkpLH/N1JanNy
6Q+2/EJYaefCrrSjxG3fFd77pLje1u9D8guCghz5jD5k7ussBLlf5WT3EMSxF9h/msBujpCHYsSL
JaOd5PBsyLpKGvb1tgP18ZX0/ImcnxUNABqCIPclCJW1nSOfNxry+xyPXsRdSrJJ3qPkO7Nbb5yB
EG4BbToOg8JJ/8FbN4H3Hmea5N30ft5HXZ+dK2qK3F7nqLYmudHpuMNhHPR77kj78GjwsucSu+GB
vAnpUoi9mZds9m1ifQXBuSevFXRO6Oz3yfaapmzSvvbsTfeLhpPJzmYXCrZFW+6Gp+rVVvmRNOpt
TNLFqFGKnkUCm5DbIKgbb5LxuvtL71z4aehE7X+yUZwdPcOyAi2qan+pR6I0MjzmpHPBCSlJxKYb
HzF7khQkT+w5711uEBIpgv8k22koIGXUVHMS9Lvpmf0BgcGD1U6mjslMW2EYPsT6xz7KahRis051
iTPwj4G7hySJbKlYF+KkvIft+pLdmeGgm4nfpIk83BI9kHBMkZelW8/5whG5M5efu6JS+A/hR2ZG
AfBjMxW1QzHqX7CRwzORWdW/wLnWEl2uIAx4cvDvw2psBgroaTtirW64gX3i7vbMYUK+lNcd3N5E
e1ox/Am9KGDw4M/kaeSNMAq60Ozmk6hR7j08kOUDzAS56335u9vBs34yJJJl9E9OgT0gj/NrPIaH
b2X4Mq7eTI8/OtU55EoRLE0POglSoBPmXHQdFVrVFvghFjIMBQV87DLyV0He88mS/aSK5M47Kwtu
+Me9hTeOpST6DLzAaYqGo0J+TPEpYFJHLpujENflxEpdg42Gcj5Q9KJ6aBl7A9T+v8gwP+hayg4O
iyYFp+h9q4i4MsIop7KMA1M9fSkRRVvW4WuCNQ7+8YLB4+u0DkXUPry5uAJQ1QcAjNnqRzfgjJlJ
XY3hSGG84QvF84JVm9VKsAArZVaW9rOyI0rWDgCggyrdpJyGquebvOoklfBTqSyBFoAf4BlTW7Ti
XmVk5sL0lAjpUgjOxWJ9PhOOcE5OG2bz85f3bJE3g2tBYIGyucJ9UwHYhK9jggO/GY2qyDlPFz+v
KUAM9SEuDT7XzxwBPz3NHnSziotOC0kyHsm4phjjXXFR0rmcpk8Nul79Bz72vrZVol4z5CYiY0PM
/7nCAhxXq32Ml+9heYHIr9Ykj2PfWndrkpfnYXVGn7PRKQLUDZ+6dNbmXdti2VMtr1yR5Qw7XAsL
Uc8DsQKbjDYcjqi+9IbvxFjanfkkZ3Gghga5kN+fV0ZF0jb2O6W4IRiZXaQlqsAI2ATeRExPMP+i
x1W3HaFPmehOPO8HzhFodYbsVOFm1eaXjjgbuuo/xOMucd4qRgFn/013DmJKZbzcGkMvgvnKWvBI
zuKJ9porifZ44NkBuvaWKJ8iVSCrBENZvmjl9yONyG2nK0MGiE5sCEQqLgIboZw4Cw7DevoB5Z6K
tU2nSGnMKMGI0hn5CSFFHsg36adSYNkKuw35jDdgwU5WvwXqUhaYBENWyWrQjQFUDCOhhPuFH/Z6
irblTV35nnTZSHr/5jA3NN+TrftJwlua2v15RKNbEdHH/Y274O1cit2LW4XcSg8Zua4phn2xBkgT
AdWhUvQoRMdD+26en9LcYq3ez44h3BVGLp0+rgNb7sFLtsIY71ZMReuNj22JDwrgPLWm+ANUQZCU
90IJmRnkjv7Tz3NRfTVvSVWopBkynb+IfLYQGhv+hfxhVzTbuRX3RI0pzLFkIfqY5iSJPZGaCYma
zJaPuuuNPptZ6e3NbU+x3YKdqPDeyraw+uXH3ScJOdrwfwxtUBzrwjw39R3ZAd5bclwc2pFxSf0K
OEdr1cdfg+ec1c8K8gcgi7RyOiKyBaE+zejHFn+FhGPX9zolIlHuNifFTf1dMbNe80GHzmgiRrPo
/h0F/BCDUxXOq7rxxeT4pvd61ZGxl+0NcVCWa3e6UUTgg/19IeYrxM52IotHEkIqMzKmORlsRIkT
57o1lrV3/4hfo7/85nLNwmMD/eTTyID1SOZ9Ak7pAEz3RRIMhWB+zPwk5WMNFnfZLJEU0g7d+KIe
m/T6spn0exKmWSCWgEHCF9INm2MhaDvV6ML6mmfzc4a18J/7UQAONtI2UZ8wymdYTa05ovBJw5Hc
+T3ZNtIbr8r7fHDyQlAlL7txKnjheZI52dY56RJWneqc7SnaUQy5X5brXvcjyhewvUhr26p/ArXe
+bbxfVwHzEBx0Q7u2VCQcaKRBhO+WdO+rGdW7EqBe2m/xbU7N2au70txvFjW8TY0BqyvhlnbQsAi
yW1bdTQft/dZP6wXIe7PScBFSUbkMqu3kiT2nkOLVjH2fSRwE96HTAXW+lb4n88ByVS2tc8rCQsb
qmLSCsnceVDO9uCzpdZP/7Ivig/n9Vbb/u/iYvvytTuzZMj+zhTuR7t+p4GBFHIsXHNAGMz3RF7Q
KQJUgMRVuLzK79OvZ5KCphGTFw6e4xPerXTUkJkwdQxKoo2THZybtdnM7nnvxfygtN7QTobtk5OM
qFmLgISZUJ5/OdASFKiJJjmLbvZLwHfkeY0TLxtQfVQQbtsxPh2A/LEemBsJGgYanzI7e1sD2y0m
F0fcXI7/AC/9I1G+X3YMs5CBO9TQT+Geehi708dgeV8rBtNt29jaIhmpPWwKfVvlojvXBW2HpTof
0Qhcozq9ydgpvc0VBSEjcsXQNKY3gcRcfFKn5gQhpbkmqmaHwKq0nzrVgJrJ7BrdjMqbyYwZooi4
dxiDq0LWN9oZyFLVR+UwQ7iXCDTGw1uoYkGA66PFOfPuzt7UEVWijEYpkOhT0LaYY2q2N7C7RRxG
muI+inm7avqnQq+wPOT9S/LFfSjwo8f7q0e2YD8A5hDXlKo8PoPe1DEe4AuaNy1pdb5Kx3wrL+Jl
RB/QTdr0zJHMmi446MLR1gdwDdCazuX97u0VESCNLSgQIVk9YTq0VW8K4j/ZBzPtiNpjk9xqOV5u
eKfB0JKt/9NTx/u90qMj4UTR8WTv03TJqV1inhEe/PNSEh08yh0yfLh+SDDSufxFUJq40bSWWlYB
Zy/IsHjC0/gQoMnJwVz1ZlivND2mHuvpCbPkrNXWoQiggJO7ErTkUkxtrzI8BTMW0iLYRvoacKaS
iwsB7jyvWbwRqVTi2pMdWm08DfxopH1qKEdjsB1SFow7ct/8wL3FL/0Y9xlqghidrRJ50k5D3PpY
TeKsKkpa3vq4rzxXIw5Vo4NpUFMdi3Ws6Omoa0Tm1APB+n2AH5uympEjfNnlzf2GsXscLYXwMJBp
WQfZUux0hezndzuocWxcg5aUSbpdq2xF+mBnWpExoDOOPbu2itory7lkS6knl4oK5SnPtBKK+voP
2u5ppiOxvg8LakyDKiIEyucK5Fzq36p8KO/QD5GUFhxQgF2IYmSqlERPkP84yxJpJ8C3kgtE3NXD
5mBv7CeDtxKfMzy4ZQ3IXk9Zwq/eiDnl4hRPZLR+VJLizZDLx+8iedBaNkY6BGIvAKDKf8mEWshd
WDO6t92nGaiUBeN9Xn/vYAft2BVKco7E/ll3+lQGnYzA3lP3Yp7/C+ndoT+W6nTZAGgrJ1z5ZtRg
DnW6ZhEEm+of3ZQ9VfsnmfyoTHMyvVzY+i2FMw/ONzPlOBNmJd4gJmCaoR6ln4L8CoKhUHLmJrKp
95LVTGyY92uYtueuxzKttV82wHjDBz/Upt7yGDpuUyYRZrsiPRjMK5zZC4+uW/hit8ETI3nsPMx1
uVPmdS6BNtJ1RzDUYlk4MkwyVg4tliUB1JxoTv2stA0/+XVasmlZAPSo0Wv+Yz9MU/zwa7gMAYB+
oXeXLH7SMou6dxTxAIhmGjZ9Mvf7Uzz1vHziuflJucGOVQ9iqVGrM/pcDawXPOrJQiCI02+yC1wO
/ZWP+8YXr3X5CWaPpiFnJDk7WtZJ/ytz3gvmd78LtIXrI+R82WcUUA7OpFNJ96CGh+avEIAzc/D0
CROOX6/5MVYWC6C7BTRUJALc1BWHNQmoOVcjfeYnANBDWE5GyPAmNhGxvHGZPxu1jceSPZCv3mqO
lyK+Vue7bdWjsk5JW8nu8Y3GWp7AasYWu5WZsVc4PrLtJy9iKzPSde2NqC5Db1hWsCzA/IpN3I4i
fdzT3WiGH5rYO4XxEC33d/afUfTkagxPnOYmg4uh3mNU6EDmVTDj+HXIbKPy9lzMUIurU+T7/o8t
Xfqe5J0fgvE7+54ZCoapmlxOA7do83fr6jkt7/CB7laKikyR0Cir7mLOFBmTH6qLggrNzS3lVALI
LyGG1xDKoWD4fMO3b2HvV7lcEJgiEQT148nqb/7CbDIJaVe37IAGCUGiFq3AGO1Abu5z8FMmBv5S
EbfReUVzciJfrs1V2VwLys2uRSYXe9D2kGsXlJ8d7JN/cJjJsen/sVEIzsA7WeJ7N0cfndnDJKWB
iwbMD4zc7bLtFgWb1z7TFiP7WteA5oe9jb4qv5jyGkxGwEefBLH/4/9ZXWolici8uHvFOui+MeFa
C2sH2GSr/lnNbaJ9pRMGlPQHOsANNFOdk6AMh2IMxUmI6TeI/mUKnGjdqQg/coDUI/Kh5LSNlytz
noQvErpCXoerB1GhICXJ0IQzmO7+SygT205gMe2y/ZfxS5FMrnpk7iMMur61dNmu7FHLc5EWveQS
YwcNrIfpFLiWuqcyUtyhHUgORa/BOOaPwTXNpXmd8uBD6YGCi8eypw9eDJ+VJI2orDEGSfi1Yhsy
GDWcJlwyTPyIXvTdxPHjPIbP5C4mqucAzfZuPqHLRWrJGb04A5HNqmnu3DEKUB3REUQPaf/OaMgX
QP1+dIg/1FSTtWhlXdX3+74zbskc+ugzbGca7Q6mY/MMQJ33ark1MLUO07L6WctSplugmc0qZZTc
xzj84OjgEXKIYPJEO+CONoEOwoOxsNdxBdIUQE/b/SDLz88m5TTjo6AyTvcGn0emKWrbd6MJRdhg
h4Xm+smENdcIUTfBsgD4O8j/5wWCNg5br33Yo4I2aLbtGqocXEu4l4mXqSGdw3LI+5xNSxTP/4WL
n4tqH5Soufmwr+r68LB5zXm1Gnt+URU4bfTrrXCNm7yuf6jOWhje1Et1Od79eIeLx5pNjzEcuJKl
DNPkFaIAyz5GYSlc0sdVIhnvAQtNHtD8kT/3U94khevqJQbc/QFm1d4QoevTtMLsOlYSVX7u2Fgs
kuDy/c4uBmH9m/L+00L30BTZh3d0yuSMK2LfHZSzf2oTwRyH0ajOdV/ny9pcNwSjBFnPiORCakKS
wcDDjO7EnkDxGgv27OY0S6n9PDlh9nGzbn7Aj44qZigtlJQHSKRCZ09FWQ0KprT/m9NT9OewITrV
ilnCBLJMWRMT8N1t1iT5UGrG3rzyfW2tPZa7dn+Z0TEHhm8G6Vbw3mwRUDvkx+3keWMYirwc/veD
ciu+20VInGMI1MWbnS9o0lSz9/V4+MMTgMGs4ElGYM+3gZSQNThBOmP4hzo+jTDNDeRcKH1umT51
BHMqJNc5U/utSJxquP2LGgCCJE0ng3MLdSU37Tcau/pAccq5vlDtuARbOg8WUEPRxzNri926gpzM
UicATIu+tJ5XayhO81x65LWYl0y3f5YqoRNPbOI5iu4LWG4i6OJuDncoUe9s7CV8SU73FHKCJ9DT
fozIO6NpjJdiTtfpJ4KpKhest8sLACFcOpR6JACU1THZWJCOaj+qSWK1LgyMeOUawsQ+pBLN6mut
SwqmTbaZLo6P+7c5/cA1KKern4FqCWHEJeMdwBU6G+TCli3bvaNteRuqRpGwBumkTWS+qgesZYyI
NqTGRw+L0/l9vSJwAGJzkQqfQOUpLctKbY69HTyRWvJ7okorstOJc9VKLjs3GteTEZWCADpESHx+
e/pbNF1aiFgB12i5O38IuKiI/fjhOAUwwq0dMGC7ntMkmrBM4EDJUR3DFPkCg5rCnyERya6oDfvk
M38KntKmAe8VXaKdg0L/HC+lF8EnXXTKJ5ihUmyo1wqbdKq+p1lKBx8tWozEce4gYpANhYhH69Q/
6KzYbk0mcX5/kxOuacZVlOUQM+fIkaU+f18sI7kGQRpL8k4CnHWsdVvQTBHEso7oUEjjgJ2J5Jri
cQ9NOkXxkt72WPsEqN81G+kJ9e4hQ9+rN085PCpfL1wNxizAHm2MRWXKK8Gcy7634BOSx0wS3MLq
auFiHgDqsYseMsXHGJG2zkRj3KX1bQEEn/tgbt+P9bgGZ8CrpFapY5XH4XRvNpizYqptYnOdt/0r
r78P5Khm/t5y56aaNS3HJl/FG22PLV/tIMnvW313Don1HMWrKSfbtfy6N0ILQqEOdvjnuex7H/7M
gwtVNJJiEv+RyyCumvtOVja2DIxiSjNZB1yH50oojRSkJHfpKMeYpif+c1xuFOeyU8b4ziLzaKDm
JiZd+mDpBS7Fvo/H0SGCk7UoR79X22LQEL2xcEDdMBfbx4NO5ZJaLCnIFI71193ROl92xSlQ4K1F
cW4RKor4O1IaSkjrVHcTcVK4+PQBuuTYQN9DOIEaEUW9oeGn5Rd5MSfRfifgGBTvqVhwq1IcJ9T5
Iu7S7+QvQdoSnG26L9oaQ60nXKNnOxwoT1x3aY9HmFXq/jkCQbdIkt2isRo1HXpRrJEvsH+t56/D
MN0b971Y9I15fdfsNjZhhzsmEV+VdLadJzvGZ9PMH/OvRJhcVJ6Bs+TOkb/24G4FCqG/4O2TXyBa
tYniKuRKxmokZ4un9RV+GDlx7D15HayoxmsugaqRp4oT/OCLj1PSW8xz8n15wnzhLDObmA9TcCJi
NbRr2Qt/9nlQ1qrE1lyB1X3DxLWBwBbMgN3UCXDh7upFz8OuuOfwrt+Twfj5aUi6eh1sYEjn2/pL
Pz/6l5uu6ERWMOyJpV21Zx03ufRZkDksgCa9GorPAMD3gAaowbeT0pYN3htIhJQIYwYjhn1fozaI
B94nB3AUJ0KbN5kNTBEMUzpxH+pOf6A6sQJXt4J/VMuCYINFaZYyOGcQkBmhJNYe8LBwo6cFcUfp
2QpuftHDptlBUr71Yj+MT8p3WOW6d7dht+/c0pevED8MSK5Ss7Ek5+q+QlLay+w87U5mFfPZZfuN
6/f0I8eaYMoTpjEs8LHXuCFqd/wMs7jGq2jdAs5+yPBZYABcQBCVqWakmb/1ANa69Yp/5jaoRQ8a
RztzPz5iCROLVuGd1gOhLctX/Nta+khsI2rG1c5vdzfl8bXhS2XPTe5cPPtVT0YtbzZIEu0apXgZ
C6M0A+PBrFEHFe4m8rFO5QXJ1bFMIWmlVVGTNpuevN/MynarQUzUAk9vCF+NyBGji4b3L6skBxQS
QQU4PT/P+U0LZeeueEcH36gP4Fq8L850MzN2+f5L9wni9WMpiRz9L8H4bL0dSRpK3AqvBeu1AcWU
GQSJ0LgoQyamVjLPCmxkozfLjW3OVdQ9jkYe+EVe5s/hdugBZt0zXFZiKSTnt5WoCI6bhFTouj9n
1rWQ7EpgwAyBQPXsqqdlKHgCc9Re3MtNbpJxRkSGN+F0s+Tul8TVu2klCrLqUNidLyrX9s6+fc1Z
LUNpYA5Cp+Olq2eaLTi5DW2IF8SRqYRdxQD63bRL1emNKM1bLjjxm66KyHFs1q67Pm4FGJyHfz5t
YVwJ1J0Zeg2s4F1SwphJLFzLwL2EwhYgXJXRxlkcJuh1YtEPms++/KAIkl6d3QxQiKR5xLI+odNf
cdI0AAjoEYJ+ICvfbUeF1dcUygiSLHY6B647z3UZ0LhbjMugZp+nbG1/L1iQqw/2dhFP0Hmun4uG
vGy2uXUfYRUqLdTQ0JQMc4d7itKQh2STGoOuDVfsa2Xl7JAs80LcbWfHpn24CnTMNtumc9ASE9lg
OGVsaDad3QzhUpGtHG2JwT2uM53mghLJ1T299UNVRmXKqrjgOFUc206pAWXlOu3PVQY6iOFhZHIO
UihsrsQUXiWpmp4YYybpCcpEEJBOnEPLr5cOEs0w+eW7+6Ia/leHKh9LsIfeu5vsJCXiZBZVH1Tl
/tVmt1o82Vdo/3aiDP4H+XXLO7zcsNG6lsdx9Uqmwz7m+vcTvKVaoCF6VUW3BRzmjgYLRPoyFGxq
ScjvRDYYJH3FMhWN4HEJfdNqZOrvOWY6YG64urxo5LTLmMTDtEssY9uIcT8EDg27ti7d8k0Cx3Gj
DrSH2HJkpeboyL0VH9uIQdC6nxn/puAuhsI/V0zTxkF4ra4EBu9ZV/rkNYvSkNSdIju5F2H7la1g
QjqWVZJuwRinw/lfk+0WxxPny8QO1NH+43tu84IX0EMJr21rxFsb1aJg2Iyykwg2/BqIur6pcJHK
OWcNIx1quVFxzOhuRGot3Qh4krpho9kyR4pMtdvWc3CDFWI44HbmdfhVIboPlyMAFtOwbYuDPvhX
+f55c2BZhor7VpMKWLcdW3Ocpy7anNj4ZbinUFuBVmB5fNMiu5uoP+nBhKwtixjpPx2A7WuAelEe
+632hO3fqIJwkE3pekn1JNCpGd/OGolkiuMfOgBMQ5K3UAqAT/sqfUfy/c4PBAHbPavk4XqbjxPe
81+sQ3DDdHrMX9lafZ22yLGoqSKdNbfDYVqHbNPHFzJGa9/VcQhKFKmutDOsaRvp21hzMKnuj65v
aWM+0JQo8eMZKC6WsobOdqUdc+GoMu4HeC8m3tmLi+Q0YsBdlMGhWWy6lFjGKH+Hj6LZXBIA34W3
bXX1SUodRs1MsT4rSbN2cerkFJG0SeOARjBqo4GrtfH1xXEBso+shilPgKvyxyWAdEs8nzPW+3zH
vtBq5JwaJdKDTK9SJhOtmQqKDyyfzumws7MGoJELgebRVAsV4uEKp9ECdQ76Ltu277KRQtn23qwl
+GKfk3FtI0n37xLw3SgvdvKZ28TxC8MsqgFD2WI0y3FeYhHaHEmAoi48H+8j4Z3xeEPiNwOeXjMf
9Tjv/ejWZcCqIbm0uynNnZOINPqkdrpmBswZXJMTUtjTK2AuALitISJKPxo1qAS22RZ/OZMDRDAE
kL4yjNyz/ShvM+xUl6Q9/v0eXIb2vuBYFfYMRzhvy8OQZN8P3uA/G+2sxJGhco2QTTN7MsIGTVCb
w7tuGQ5NE2gcle0pDyTCtv9L8MisMVMcWEyI7EcX5rmArcH8fyFWh3PVp/PNgIDWAbKeW6yVsVQD
W/Nd0F0ZJD3BSqR5DrVXKNB0t4vF966u7nxRWdtSIHj2IHvlRSm0NRGsRyZyS4fBAVU7JC1VjebB
xtG6wAkaPQkIRY7l+Igx/ismHKCbKdEmKQ7MCX+zHMzpmrDjgv7SJhgHC2j9x76EOVGJojK9nG6H
CO5S6EUBUX14ZdWEsS8v05FnDnF2b9Gr62GLtgF5wpaGR2N6IXmczW4swO/WUAc1JHIFkXBjwYcN
FMG7wG+GN1z3HhRKJkKgDy7ugVjB27MpFJT57+TXfyJur7aMOqJdK7qTVF3FU6FCPvD4r0HppgiN
h6PbdbWYJxZw8Kd+Yr9AYGxvcGReGNuNK9nha10pU11ReY/s0bFNrwgVOXIJpuCiJcdUaf93m0qA
UYchwFdGIY1auUMR1Kby/ZCKZaANKXT9cxvMfmqJEMFhWugXO7N1DtpWZ7oiObfugI2tkTWDF1zb
UaWtD0QR+dCOKfzx6XaW4gXHodoIiJxm0zEMtxa9byzObWaKTX2xDkQA4LjAngNreUIJ5LRvOJf8
/i3BQnd4Tv3ok2vP6ib5p5PhUs+34ClWE81Ytg5GOZ6V0a/8TY8136NwosKPROo4YQpANUChmKER
S9Xufl/DrUmMYPzhl+OJRA2FQv3prHHP1TGs/P5EJAcccwxYVvuy3BGNwMv7waVofy7jolt0LHOO
darUzvLzEfcNiXZ6PVjV5CCRFOQAx+k+lvnXC9w/G+m0L6ziygxUH5k+oE3bWuB7jK65aIurTQhG
ib0eJfMAx64MFwM1ifn/kFfcEN9krhHl+ys3MbClxn543QUeM7kvOfZ4o9mAWHt6LUsAz6+3fEO6
WcNKbTGMvYlsBjsy1vHee4wPV+XLCV5X5SEhysoL2wZ3ceHQOZ/AJg1O0JvuK6kGoNGVkNp19SIk
0a5oRO3rkKkl/rMqETR4s4R268/q7uElcSm4UJlfNipSt4IwAC/12njoaXzudepGe0vUtdn1Zgqj
HsNCK2/HJ+KXfLUpv3qAIqG4bx0QiAklprhl03ZJO90otDLClzptRIXFlAj2G8q7iq3sojXMiau4
7qlFAdiQRtxplk8MGDwX0t0MCCOdplDy5OPAtHShc+iJBjPAKN5OEdPkYMaBXol+mqtZOmLnyIXE
3PYWc2jNGxAx30q9DFqhIzxurLApXacHMAVE5Fu4i+V+p5Fusqfx0UVC2DSjBQ9WIL3jZMVHq7Y9
2q9Q1fvN1tCRJfbBCYpeSe1aIJwliPslSRIbc49laaexatTzrCmemmw0bX46/u2tibCt30ndY+wA
80X2hzecC3Fal59HeLClomwoX9xiqdCBOFSQzh+8yaquUo4yttcfdQZz8fhOjU+d8KVhVJZpcAOL
uzMjMdJEpeVkVOu9xFwrEHBE485en5ggOuCRT0NDqpb9WYty+M+fbwrJxEsQn+nIz2ftCQyHNmKv
RVRqPigLvOM2VXjC17FqWqWVTV37B2tBI3zxj3dlm8MO571SHVOyw55hV2vrnvKQA+JcfmPTeut/
C7wHqy9WLHGGDJcZJLM5F8O60c/17PAYDoIHO831hacsMOE5Fn/rzdvPrCsYv97RHUP2GwKdZvW8
KcLQ08GbRR5WRtiQQjUU7cCw6jGmrbU46IdcDy8/inkibKLcsOsg7umcvTCcwN6JK1xYiWDLoEcu
tEsw+1YCNqAdUYxATC7Q7MpTCz0cqSGZ4likt7K0NeUp91p3hABuDfn+GLGWyaO2l7MEnf/1f4yi
wsbSgbQWkFvjPGOFsCs8/006Q29QxvNWNKxMEpI/wR65VL8besVTWgFfaL5+bIGzIUyEi2Y+lcy5
Ct0JS7vhlkoxeuEspCrHk54KcOYJOW5Fsbu5EASYUE4NzCSafUbiUmLhO//715x3EZrfDU07Vw06
caSnvYHu+rczj66dp1hZvvVlbwuKbv/6OHC6RdPczzpxvIa1UYBFAd2eHjFKmrJPlCZU9+pms4lq
9P+1ooU0rErniIx/eSz5dft4MJtdgJ4v24JxJY8D09YYFsFnFySS8gfVjrOLVEeEBisdhZ4Kt5ft
E2D4LGOSFTsVpnO9xDm+GIL/he/k8M9NRK2Qny0OiSA2nEqsMFgdNxZaNwNmxBUNzcG71lRO/VEQ
5RVeZl+KGNdfuWGQUFUBIj0HX7PAFEWVK2qliWxg8ZAcO/vGfSlCOyDIaPj8PRqD2zOPkC1llfLq
buJiJJ72RUrdv43q3tra955BLNL+8Ff0lp6RQjJcik4C9OjbwCe4FwkUuwz9+RCur9174ls1y2TB
7JloK70KHwEvhYBpwLpf5iquBbMiuMSH+4z0eyAyfg9HrI9qFhkB1mfgO1cRHkI1GzttWsywE7tE
05w4SNl+CjuaASvfZCoVKaUGDKBGhpDJozRFT4WqTytXIB1rKaYuqSCHxO6qNNasx0Q5fYyxKOtf
pa2CIjfOWy0/UNHEEd2bLpSwibT4yCBAKnjjCR099Cg/h4wcbEZGc4KA/kD4x3NfuRgXrYXfnnGN
/wdKIoCIct1NWTzVDXqcjJq9H5wpHDpOObQ8hLtKpttZButjw/w5m3HcaIKih01FseKwN7rgx/ox
P7Q+pgnCGpy8hLKMaRw5fXWIvnUp86RuGQmmKh4B5v5hLEbFQ9fAqIjoeeSDoLOlg6ejhyNiZMY1
xiZkNydkXd15aZsf3iqLInvODDlLHa6AhDPwiBNmQiNp8gyo8/t/UoSf/LIBNBAejakSoqi+rFFK
aWqleQrUnXPddbbl8Mf5dgbyrncpDkDQEtzy3JwDKiavNA4Isb1n/8XGogFggkJVxOVcXu4rvHY1
UIkq34qxv5JvOLhEsBvwfisHIUA6IhONh0JdwrauOFhdF0iT0sdkL64+94ZZZCC87rVYTYlFRs7/
rvoplA4GIMHU9gG1qfepC2dOjjYNOvWs1B8sNcq9LBJW/6/+gx2l9e8dgW7gj2JANUhMhEucZrC5
iE30TqqSn6h2E9HCm6VDgwsCugRtDDKEY27cKjfMqphhsM7DEXBEcxjz5Onqij7cjtd23J9zI2lu
E7JoY96uC3SaU8wJtVeL2/PthCdzl0NrF40JUe76QjagPXd1eooZKRaPHBnQsGFPl2jJ/2/B1kae
BEbs/Jd0xEF6BCuAIzqJosMO02HZssdm8y/+Ge3kS+p4IsSpt9fiBhUAgxd+MnYs2Ew/IRZSlhKD
wn4AZlIa4w56Nk57wiMXhYx0Jvr2g2XLRtau0FZpFDjP434Jd48tM7uk49nC9uNYqpYteviNaBqR
D8VeiAONG3S3F3B/Nk8amkLRgUds+s7SelZlg7zmI0WxlvPw1alKKyw3HDYQVHRsr8Qi91B2CZf+
pegfi1oc9Z54NH4lG0RX5huNZF38BXgGgHhGfWUwGUo1d5Qic10ErhzylEbvhixCtUVEYAKbPpjT
nvb3MdJBlsT8e2gfFgaamezr3HLHfHyyDXlqkiBCLQcwCFb/kXlqRFxqiqzda+ULlLqv3awB5jg+
5IvtkJ2Q2kJLQ8aSD1s+QlrQkkz+hrh5LzRguuXfGkWXf0aVU7Ke9uXywvXXyor3PeSPaK9KQvca
d9MM2hfbZA6hPfuFGV7PpBIKKv+MHjuilmKjWzeq60P+xTTyPkmOcmv2PyTYY+N/SVmvjfgBwqRt
++0KTQ/dsnI2+wUtYoYGR4V4yjcmeTlr6mzd9KM519YHEx/Xx15MJ/p6sXJAtxg0DRJY8UpTbzsn
HAklx/8fDxzYSUg28PZIpjWfB/NaN6om6ksAti8090QUDqPKZ82cXeiW2nEqjUwQkiO3Q5QEk7Py
hPd7gn00weu+PkCC6A7z5iWYtgR3Vue8wRMC1VqcabjgWjutHlqhfOlot9LUBIaKsemFfHVL9BnF
si2oNjtUln69LQ/KH60TsakD7Yq5EpHD5xXKTVR5dxlweOeopEkjz9dvwre0lzMd8BAQmOFhvWpU
UexlzkgMolk3sYXpFWUs+H3y+hSgfV0bnzvBeR/pQI5I8HuNT49QotofYsd685N40i3SIGCnY7wf
fUSAsqYgGgnfsFDYxBi8yBoG4DJd9UaarCzpgDg/pzdKrgKRZ03JiLkm7ucFk3qZ07Fbma6ykRkp
n6lyZX4ca/W94XVkIM+o1jCulJwJyU9goawB1WdGrk+Z6oLUoxh/j4DhNVVgUyOSX2tTKlJQyu2I
MFLgPH5cnvB6LY+Rl2cinyYOMKFuEPxha4lLXBa9VGBCk8AsUnleFePmP7EBKXqL1Go2nond0Xn4
ss8Ce7hYYCawt5ryLaGjf3ie6mMw/KZopJhdg1HqCHIiRgsooSeosYPNaPiHLuCb16f6tTLItVdX
Rykh5Al6rC/1+joK9X1SPCv6MRLpoU6UXlhejMED4MiIfAtnJR0g/xVpj0pSpEMQJ/3EM9TtiCCh
civLdQRbifb+2Rx3UGnkMYg/A9tdAVTFza7hEwr15cBExVbUos9cOv+a67M7x72ktBcPN3K2Qi6V
o982AN6TFjxol54aqtswKV5xqL8qaRYVuTk+ltjC0li0E6yYB5LS42lwH2FdxTIw2c0uN9Zp8B5Q
J4ZUBIJWeXfJKs1tMn7rU/C0jxH5erqoBz78baa2fRqNMjxnz2houGxPhbfGcLWOQiSsE4haUaNp
FBO3mbnpV1YxhT3xZYTOT1z4S3MmGaBWczn4JNRHUE2Sp1q4QAnvkUFGnbyZQoJSnlVVzxzybh+P
g54R3vXRp2y4CNBTDxqfJsWYQlwHxzahSVpzd9bd48JtstUrHVOda4b4fbNQvZnYyknMQA4eBj5c
82tHAnaICUj7k0V5e2+i/kMg2MZNiQ7UaDmc1Xv1sUtJQp4n/hPqBNWcfqTU9qwtnFxxhbzHzAl5
/+4pqYzuF3oFF37ZnJ8fEJb4xZLKPEG6d1db+a/nTaym36OcKs7tr+O58bek2Rxm6dc2nqLxStY9
4ePLplsxBWWbFw6zU8mz4RTrni8sNnhARA+z3/zzYX9rMPBH03NTsGMseRl/63n3bbsn5gdANZys
6u6MSq3IVYgJI+TBPuq5zc/tjAxyL+xmUjcdz8aZgRj36Tz8mKtEvSOBQhQ2pE4qxUvX6TjRlL1q
8BrpvNBSDPT5rFzPf8oRaalplrxsyJIH28lMuEUuT5h2DL0hSY/yfIsQm9v1qcuTLqHlhS656col
KDXeefVDujfK1oMs9/9t9A6VVQHzcmsy8Xyn7pvm5Tjreh3attyK2MP/PyUYZ7THdOCDLvguWxZz
lG858PLz2thhapEBUdv67l8ElSv/SV1onMH6lNoTmX8kWIgRJ1ZLESf7bHjaQ0TScjStJWNcVS23
EBGULuH+RQNy2BcheoiTKmr7EH0wR19POq2yIyNtuiLiQqvJp8OClKeUlaObM4GxtMWXXzX13eZN
tpOiYtnV9ZQy9J6NYhTi/0AO6Ythh5AiW8cmPXHYc7qsenFEwrIqP4tHWRX/IuEVadLgi4g7H0Ct
mnbXnuHIi9Lp/NO3rmeexJbGxMLIAUggDaa7EOM3P0Qpxyb4Oz4agGtV0atrFm56zFMd61urghm0
u/8jbbuXoDlHBvN6mpWjT1jHYsCjGgNmGx2/kvkXRlKs1dsUUD1AJJdyfWaHqRjng4cTN8Q2A+2G
BVLiAQtyxgJ1lA/KJGTzS0ubOxUYKbI9FkG+Y42f5PdbtDo4+sSBqLEFsh72VgzVOyIpK1upY1tV
NLx3gQx0qwa2Hpx6/L1Oz9D6emRPjouwwBOMzcZH/TFZRpLy1c4rn4RocDHClS8YpGHgrZTbYqYj
VOxhzmCZIxeZkd3DYXFwzFDE3NR1gZoTq9sBmcUJwv1hQUGwymFidcpInxnqWTF17hzXFH95ld4Q
01F5TnwePP2FoI27GwbU0Y1ZEXD6uR5tDLZ3+T+gojVD6VDkU/e1J/kYCwbjvkNB7zNWidZMZ0zq
hnIQ7vyUE2SWgdLHvPjHgvXYm/+QdteDVHOMKqcYOuOzU+V1UQCmDMvdjon66OgLkYhsMwi+8D2s
7zAWa6K+4kttZMYE5vhtMbnRLFJ1kGTzthqKEQaIJX5kLqhI+kEqoPdn9E/XpsqqtzcyrfAPa8f/
VZTWQLB3tlJfO8Oc++ep03620pp0z42oHyDdMB7B6j/IW+1SihbZOswpJUvhpvWGD+KGbnYbjCAN
Rhg0/PzDP52LMSi9LVjG9D+NBEBlOumLMhfG8lH1OJGyr7X1bieqajc/v5e9+megcZo1CWsaAyZI
qUcnI2rXkVw2tz0V8ARVOPt7EGYMv8lCADOSahT+mJxTsDzFcH6E8Ozi1rpXkHkaQnfgR7yhkTq2
I5yQ/2H80vRLd3SxAPRK+tj5I77xtF1nNgnfyoAXl1aq+tQuaOvaWuSaGudLnTWx/x4yom75h/zL
QakqaI2Knh8T46z48tSv+WEhrXNrQc0vznVyn6JBltQ6YuTc8AGIEDrnmH8rnqh1pRdDl+9B9T3B
531nkjgQuMuHN4vOxUlFTfJ3L/L8KoRarM5I2zpMliVqbj6uGLfj7SK5s1kybHx273DtnBGVa4gn
7+prR3ukNkzPqBanABpz9vLfJosaUvLxDB6VZrsTisWQ01o5u34X8GwGSJMEtVP2T6Pqjw8clpKa
KSXqXGDcsE2NKpyBwLng+kGTSMRs+EFvKXFgjEeUsLRSv3HCrUEJcDOBhZgVt+YXE0AsW4RYOypG
lMWOr4X9ZAQl0GNEyEaQQZnm6EbRtktV1LBqNw1aD7oFDUY2kkILi0oiX+hETJmCvl+h2bGNKLC4
ZAOwwocYzjZLakuDNiENTu0WW6kfeBDaoJuHeCj+BCmFjmOGuvTeJdU5DDylfh4lwFLf637MyGSu
ZlF25+vz+ocgu5EjP8+DxNNUGopnmlZoosN7tfNS1W6iM6DlXpxp7SyLpKt52UNu0XyLLVAoxHeS
vfR8v43XYseeRUHGAwSuxj6qebup33m6UlC6fUHkgbQQUJEy8g6PmKBjHD8A2SNriIqQyfputEQG
q3hKlUJkYStccFGlzIDPZHgGh2+KxdbgbiLTmTQp2Qc4GiODtsC38SGGle3px6s1pW9lk9a/sTIb
r2pGIjm8c01M2l+E3XrJfdH/VC0iLAIGhJcX82c5VYnyONUkw5DyhP8TBj/MF1lkEbFJ2YuanEAd
asc+Pl5g0bbF6F6sGLgSST6snCjNR0Cvlq2tCJPurjHY/ns5zQj/9PLb0hVo11uMg9CVXPxU6JI7
Eh9/dJeCMNKfONKT8tBZyh8DfTQN93GLYMVMjjiBCxDRhg5F0XMZTKovWd1YieXOyn5YQ/exneUC
TPdFDyufXU6sLpKg0fkekjMwD1COX5o+DBkRDMXMWCKdcgV8EH5FamuATqCWJ3X1mIvpnRFEfWVJ
V5YRch7hP6th/I8ofSYePNCSfkQ+OkLUFOLD0+vROzLMcFguXi/VuKhCAlByc7+tU1BGyW5jpOSd
JTaifUSUkIu2GvgYSs9NC8V9vUKsj8JKyxw5XogMCUWwPLG8k2bopj7NQubLO1cDzV+fiwJZlVc7
2sSBt4G3RjJaGyLyfi+hbSy5PmighimIAUH7wMvk8e+/YRx8TsiIpFjOpMlCZpF2/vJ5dmkigfAk
BXbwWiciA86OJi4KY1kxh13wnscbQDrkL+WWGVlZVlxM6/+NwTiBwBDdfHGdrlNr9opN1deQSjEz
5Bi1TDxxRJWJKjAETvMNLKCrtYJfuQoh+lQpfuqrW4bOJwBnOu5aL03HTOvrELN3l4XzCJ83qtyK
NCnZ5LhrrrjFM40slSddqd/A2f3comN43klYeqCbgx3Djky4g6wE0Faokt/9B3J4i/x5DDLQ4iln
dL8Jri58b4WZakMjKjZjPGVUkkkhXHn/GfxtN9+PrpwIy7X3OmiNQDI+nmNYLU01+gjgq+azMK2u
O48tFceO6cNg884MtF9b48LHgcMuvW7z+x5VPtZ4d+WrylKgtYT8bVOWOLdOzCSi9Yv7wS11y4Sz
fj5lSrNbYEiLAUqFbP+XgJi+mngLUi/Qz24ovRg1esfZHmCxj8OD5lY1ttBCo2J8QWlgg/vxx3g/
QoStpK8v1zwqisqENtN00ZN7TJiiI53qfBdu/1Z9XOPlOdRKE9uF59P4bPiUZilie7pIbTT2tx4D
NH+U3tp7SYK76EYN0dKA/o1q+xE1TL75MBWKtSSDFY7hR1fhfQ58nuPpOqBG//iXiNVzxuqy/gqC
x/vSiasf20l85i+TngjrBmca5CGpbTH3871nmNle2kah/XsZbv2SgpKEPqGNI/PA9Hvk7U6qqPH1
OQFsWDaKhZCsjQ9D6M0FQsET52K5z82rajrVL9CxxXFnHA1n/pUJVWm0ijjiBbgh8y0L076c/FP5
XTNxt7NwJL1uaXDBJE1P/jJFbJVCVlWRg3q8H6ZoHQqWn1DCd9jYdVb08p9mxdCnZkXxFkMt2NNc
v+7iPzQXtVZuKjw2pEgcnVUAw8H5ldSDakCPh4JUZXrugX2IP1O0jHEQJMkx9oOdGiOqaqVBrS/m
kA3RrBww3X2dqULGYi/AMMkovdokEztfCCj9aEWKUQeejuH8ZUrnnEtw0eVnjv1nzK4L3VPOHTwZ
Qcaun2tcCVQYCeDgEFaUsj+0PH6z49Opc6ELVkHRfIFYZkYXhKJnk1sPJ1leyjMO8K7duliC2CQF
XirVlN4DZUsXpBcIk2u2Er3QXBLAzmirRlC2vzeJKJT43CiRqd+Wq6tIfNI9ZFi22nU5Cl9NFp2r
FZAoRMKTSab762hhzcRiEnStCEEWmGY9C7QN9Oko4HWu6OU8QCTynX8ingJxUtJcPAMw0Lx71xIh
xEDIrIADKnZt8I9xVm+GAc+v1MeidQHCdEUkXeKROt3ScJ4eqEYC5E7oVY9YbQS78OP3OyY44S06
jJbJZ24GSJcSh3N5fKNq/GUpYnfl6KdEv6sDvnbYlTxqgxngv/YahDu8lmVrfB9lChEO4TW3PNku
c3afb6ISWtGJ2CXvTvorEC9OmRfJSW3+fU5dPtDRenYc+KVW4INy8sZlSO2dAe59CeH7MAoqdqnu
xpxIouZzXWvVwNT/wPuX3PtD+LZuGzGKbnEE6BNqXGznLEV8deZ5iz6uUs6Ge7Vjbh/c6sstTScv
hbpy/rDKrJYnr0YLz/mISunSP8sgwiN0hNJUT0bE84YdFVsxF1YjeL7G3cW56xTTO1zrb9+Nf2bt
AyLW5vTTevi+gF0o5Mbsg64qKrAbYrOtCui1Orlgx+GGh1J+P2zNMlnuord6idml1ohRYT8V2MKo
u4k13EHTtSVpgaU+126LMy+eeQ0wLB2jtOlnQRwHeC7OF6bcX/8sJguqz0kJUd5HDLyPNGUVcbZx
F+QdQMSqx/gudckEhQD34JPRBLyPLmlPpQC4JzbeGFCdMblEhXRO+s+WXu66LIEkY+TLe7WFBr0V
eRoXBa+SO0NWMdslwlqFlXpeTp13ekDmfpBjPNp7TfeyuZqPCRbeGkQnuDqvwP+dHLH/tETJt3Zd
eCXotZIOOSFBqGWAycYxLOK2uBNmokENIZQ/fcXI6oRWgvlFIRTlF+mURAStKKmKucCZsqdOL/pa
7rSyeFprekjbwpRBjYLwoS2JsF1WS6WO67pBtSdI1JDlM7lwDUA9NAg9Iv29mnZytH53X9i8VWfO
veYRA1D8iu38FKAMzllL2i9Ytx5KtCEEPHoWS2QzWkJ0sTo06PNHQceTAMrqNtofOQn2Eea4spQj
f/A+ZVnTY8fveDCt9GAhf1D9teiEInwKobDh1M8OEE1d3dzVy+CIikytjKsN3zaRNleFYK3furMS
PWZrOBSRqnxxSPz2fJtf6iopRFoyadPlkhszPXExqoQjnd10rfXM1iKgdk+mUAgrXUpxRkhU9RWF
odn6sQtv2RR6Izwc9GjHvuSNXHXrPrFNCgEp/F8O/ZALNg289o7Q9SHHb97TUMfVW2JXm4CCj2H2
pOnADdw4GzPUxyO7NsyxJBV3pmYDyMpLki1WEB9kFzcZEM3hLwfSColPQVMWksNpqfSWEpVy5szZ
Z7qJYyxHchSONMYHtqNCWg9rNcniEevaM1cOcC1HLeJOExPN0h8OuiEYvqTLoaO7YVOkg4exzraQ
IUcHn+r9ua5DTbvaTxTZ1dlDXMKGtIQda17MId02jeqQTW2eJiBY5ItSpDeex1MJUh7R/IoDEbUm
i9SCi1px60zRpX8PZceqr5Sw5DpSDYzglDwJiMV3T3vS1Y0JwvOk6uSEgbc5fknxbNx34iIMI4d7
9pQ3J2s7imE/V1kPwD22pM9sRO5Fm9+8AO35kFeeQQaPvcXxuyfll/2J4wuS8VEPMIQVd0L55vsy
8Jquc/T0abOMw1I8hym4xi7vSN8DIm8NdO4xrJwqLIcWgokGIYJ1lndFSKKc8j42lb5oEyXThSDw
2oA+SkEI83p9e7s/HKNhNsMuLgGEfMoXwwo0zKRrLWUbobDBZmq/ZzXLlA62KOCgh59ecfo5TUfb
vj9SkC0kZuvVzULsx9+1ZYwCRcIOHXzdfb1fZV83cnpdT7OZt98b2IeVjeSKW6fePbZAxOGPcY8n
gEJiVxcYcIwYV0DfkuJFDEvW2Uuslw7VDfhPizNnZuSBhYv3ipelEAVH+zmVx0ydI4Nk1L7dGc9f
w/TN7K2GzLG3FNA5Z3oI0AC4R4ZKArWelY2/xW+41jfqqcY4r85BXLam/vVrL99TE8oNp2SvXsWY
SxbbxBtYB5+ZyL59E5vcAUfXcZ3Eb2oFWECgh5Ug6rs/OyFfipmcwtrZ7fYtPDCXie8hhdRgDYZQ
vuY9DoI0GqE2N5T0/k3M4dJcpUwlJNJ4JkZsn+GVqUTNIF6sI1RSPHs5TFjv7FB5oxmMSA8U4CCG
Du75sQYQUD2wA+vSEDk7V0iNaVAlq/XL6w5x3Qj9Dg+Mp1nXopCXglWno7vcqKPcKsACgiKFbKxP
Vz/aYHWXtKr5lSfJLSRMnx4Cw3cL2loIgG8Dr9bubR2luE001C5cdNSi2B96QdjhRyC3Ky0FV+wV
Pv+PMJTAWDF5Ia7DL67c9eS3S+/y5j94AEN5VXEer6Tro3VKM3aMjXDrOx4D+4v3FF+GlEdXbAi1
gqM2CR82BoOvGrOwC2NkTeAr/uiL01ffS2donLramnXX/BH8Ns62skB/fYecMdyAZN0W0Y0SN9Hy
0SWiT1wl1EokBIDPCqxgs4GhW4FXpmufs6UrIVQcxDjnNWoOzQ/+zsk29A/HstwlACc33J+kO3Wb
4h/mqHwX/P4RjMhD6KvhSHfhth39XrTQs7PZmNmKBZKCWqUBWuqybg5vCA09tXh4XwESZjJvLbYQ
4tswxdJPrDLMKGyYLlrKPmQjzRDFZYuvDkVLN/t9kOZN7ndj1DvKE8hfxXb2LuwnmueXRVwHKdD1
YRUrKYKQzI3H+Fm7DlqZz3xswVUeLU7XociVrh5zv9rvd4qcmYgeZvkogJ9jOiayVBqkZxAcd4Os
aoHFQxHFEih9lDOJ9cZI4+0CsLHHGK/xpEunEROD/xDzildUYRWu5+9V755fGMpFaEt4HplScy2n
IeEWFHYdLrURUTXKkwlcJ0UTZVn5aMREOj7xHJk89a/l0uvMOs3l1Xk6epe1Guj0im5n/Yz1k5/K
fAxhRqRQ9BywahegE9wUoz4/cabj9KM1TRZF/kPc5mGJE14SeqdOMrxHOytKQ7hNDv1YGrrQMWqp
JhM9zR+oSA5NihpBBZJ+uTs0cvbbzDRcuOf7vOwFuVysqMokZdct7scJpI9QtDVvJ4KW6Ius24MV
uZbBuUEN9gTUKsIefzXa5E7freVcriJfc9mjOOuDr8rfbuGJ7c8BgiNt1UVam9oskGTk7DcY5gvC
KRwcyMMD1nw/sRl3SVAIhrqHPwql4mc1lDuryjr7pf9jBfNpFUMMahWLZS4jbOtUU1wDsbivDAHE
anosrzm25NJteX4uwYvPRQELMhCmyp5phmnBOkVohDCRLU62l8NAHAX+x4cZDzVvlMe4PkeJgNd2
Mt3y2StFD76k7pqs4qKwqAXqYr8a315VuhglRBIFUUDd4MrjbDXAA0u+ilPiCsxsXVH/+2a1tRQG
JovUARBSxrSG0cCCLte5Jx97sbqiT/IxTp97OAbGOn6lVu+1DLYv18K4Rq6pHxFQ9L+D+ruFHcfq
rO+v3IA+mMmgslKQreSBmgGEZbkdKkygKE1NM/NGvcMonGUjIaay2bzYPcmKFCebfvWDCWvGZ65a
Rlm1qsqZ833lCpwAFNXrj9Q0iuX10Mm7ZUQnmo4tGnZ8tlx3fup9PJoveyf5AoqgQMXI65uXutdp
UWYHGicx5LmamSzcTPJhsC+PxCMJmBttSF0htBaz7ME19QJE66eOmudhdTSHwPttzQG+ewOWINE6
GL0jzdFNkG/y3y5595T3IXMdSbwo0RiUZT4eXAqmoGkbALBqbV8WIASX57BshUeap4J4jQ5Bim3R
1AaWOZMA2PrGSYPapdaB7/vD/d+Y92W5X/lUhfkolg4cm3fAc80BxgFI/fokmQoTGAXmeTl2lNVO
iHAo66/AhY/sN85Vu9/jN6p/QEMGViE+CM3vSmXzLMCklT1VyE+tdcPFvBn3kw76a6mvQSR49+Gj
+nXK48OVBzTZAIvP5q4Q30YcZMGQc9w6LoZIs20q6LpES4C/+acW6/mRzMmW3SWJIaswfMHkxQ8m
tX9SKZdrXRoVxQQs/lMod7z2ElATIBrKhDNLjFYA6tqSq1QQAm32BN3jwk85sxzLdxSr4XMiRWEu
PepbOWmdnF6tCOoJaxRrYcRZnHCRGIcJmyerecbqj8CaElLqbuldzBT47v3Uu3hvqHew5F39SXwr
poF0Nyx8UEmCMbizoAHm0F/vxQuuZ6EV6NzGGKT0gWOJjReoHa6QgaXA4wvR8FXTwWpYhkexhFJL
/lL2pelKA0KM41roMBEXKVwwUh7cTyGBJci0CME8VHDuD1+nHGB/wEGZyWXUv2jiTM3VLVeb8mTn
AkikI2xaX/6vBbbV1y/hniYV1JdiJWNa5+V0GJSeAEuy+8SlvysRJNd5IqMq0GFYjXgUk12TlszT
Bl45sfE4UkfOXG8xf8MaiuRde/wKrRq4ZTNK17T6LGowLNBZX/FtlvwjR7ZFj8KVATo6erpNfZbh
HfFLGeOcMHjqxGgMgymNs2QQCm0P0hw5eDHs3ZQ7NTwPMCpCXPKfzQuou6EsJ4MfZQbsb5kRrVbl
x7rVoIpS/MVP/B+cK2suINYhR6eqcvbZxaeGPBxlE3xnJ9tyuodS5QZLyAbo1IVzMZS4ykRyDlwS
PcnWccbEvykXH0PyUFNTgmxQKh3CGKTXsxx0r46n7K34ThNjksv9X5ofCJTPAyecQhtQV0l3WTBX
bm4Q2BDOqFibaKSSMuUV0Vnlfu6J5rsV57dHBjiqHtyPNVtOrfoL0dF/hoUe3vZqMUVBjmPIsmd8
iqiNyG6ldJ/eXCgNJan6yFSGuO3fUZnyrv5S725CRAa9PB7Bp0/ccI3US3ZI5WYR9AizCemAniRC
TDYh5+USyagzo+/3iRysaNKW4zaaq4I1P9Ep/wTG6OtDeyMalAD4yXl6+3Vg7kuC9iyZmzgwFuBv
k4qzoXRfJWnbwpR6I8z1RGzi8gRMnScUDPMXYkEA3NgCd0mQQ4TFuW+m8I1avt/ZBs/ddp1cNxIT
zBodogCJttmMClxvGM0uc9nz3GtyMYasTwldvD3OseAoZwe5GwMQYpUEiUC7fvftjzBTfYAPPyy7
chA11RotqWbiMSgHl4NIKhQscRajYLhCSlTE0F4xEqpeB3+QK67q2qDL36qelSngV2KrcTQ/mMBs
twObRppSSxny+x5SxHC2S3aRwOMz7kMzfBYdfrNyhkSwoEf7KmmNtSBIgWNgKBGMUX7W6yUhaI76
NhepHNXoamSivLhZKbYgAw3T5vbbAVbCpAuqG22w/GOHzfk708mCfIVE9G5pMlo6n1AhRXtPxDdt
FNItaUTq/mSEQfC5NRW5eTKvmZnRXm2WEFhoE4oeSGPFsmlx0rDjq2QYoXelaxtI1oQaWbaLb/GK
WmIOCs7oTfsckxJ8U+koy68VFXyn82gEoj1mTy9RhSItZiSPewP+0JOe+6JFqp7Ilp/GAJyLEJWx
7Ukw8C52pJIs114iuoD2rFg2WUszR/Bbk4jdUDKHMMPgoRH/9SXQvUQaXJFXLIaVwL8O4KkWY/bE
/mOzfRcclT1L0GckxoRJss8+XflwHNUr0YrKUDw1iHKEqVyLeryTb+jdfMzVeXbsrh0zIah65Lrq
C6QzK2X3rlDGXLz0aVPziDKXYDMY7ttOUIuWI5sP/lffas37dwItSfF3AItQF/cMe2p9qHz0Kzda
PwS93S5PwGB073ImWFTzdce42kTge6G4ZyFcb2j1qp5Thvg0kYqbUgH/YIYXZ6PGd/GHBtjSK+8D
XxFzdm6IVY647+IwPhhw01LVjvrLTtuKO0xVpNk5pgK4eS8Bw88KFumv9g5LyXPG2UqEIQ2u6n0J
mAE2Cdny1LT635XiluyG9t0qnBSEez+X1mNTAR8f6pE2sI9r8p8bjh7zoOgv7QQvHASHN1XCoprx
qGaimnlN4erB6/rRVZ5zPloEKm5hsMvw9Glq198Sji5ckNv5+Dqbg6Glx13XwdTU8Ow8nlwlQs9H
PM8nsHMYjSaeqTaN5mIzOdWs+kshLuV7lIPl1AQbX7fg+kv5k1dGEH9zUg9aJhq/NWGyI+IDt1qp
zWTNU/S6++R/t3i2Q+rjtxe/Lr+iETHZgEj39ypIsIku0lt3QWlIhsu+RvWs7qNw4gBE9v+lRVp8
4hnyq9c9SVkhq11fIUoMdRi6w5rwzuB0vYcugZpJqBHyIZfBAsPiep2G4LPUs82aGKIO3eDiTeLI
q8oHkaR8NLCo5oXu/ZMG2tNvI/YChw0KaHI8rK/L/LWs038siPhrcWqIie8/HAx5O/n5HKax+e1v
MQU+3hvWlzB35dHrZNFRQG1fu9bMxZRGJoYzJb5qGbUptKk5LRYi/yrNTT47/7ZdAzAYMOrlGIJH
kbkUB4DT3LYJgt7B54JI6PdOUzgJII9ViMwHP7W7yb5w8Bk8s68JXTK5LpDu8jS4TuLvCRmKyPus
aanMr9A1rsG8p9A6I78aHOQ0c8g6BntsiXZTD1H0igc+ZQdE1SBz4qjj3Oqu8+1w5E5aBPeZpIGQ
ZYAmhWMTboyGFuM2EZWTl5qllL+LfAog23nZ1HjRWuObLKW4tAy8N6BW+Wp25KDMb6Ckr5eb+QWb
mr3ap4Au8eEgoXM+21JiMaaf1ExoUrcLgecBshK171DKZvCXyGbau1XhRJpb4K4mz9vqaxofmykA
hceydChwYZ4taiTTRBa8h5XrhWHCuZJTU8lFWrxb/1rLC4w4eQLLT7iSiJHdGZVsS1Jgjpr9c0f2
f7BRCGWdkSWe3TdKFLrC9GOLsQeecJjfihDlNTsTZn1P6dUz2zA26dkSj2bVJCqabnr+hgIwBKqg
YZo8rF2V6vjyQPQPwlG/3C7Fx6ktzvNXeQsHGwOfTL88RHWYSHk6YBoSZi2zMvP6cPPctiiuGcv1
sI8BR6eIlur7BonXhv4C901s7iLRg1Fab+5liGS+MaXGg3WQlbNU1yBdW3/nBUbu4CF996dGLXwE
C6oDD30/7Vd9xyOQGZ5y+BPb02DDjrj7lLA8OGhMOy88i+jeRMKXuU0su9NvEY8wEAzwUQEaQ+9A
nj3f+DIpR0myjFUbk5GfUVpDLtwMKrmXuhPINhQh0maWovX1arRpjE3LldGULIMKpMw7DPicgcM4
SkTBp19cLyuIcSbJMvYW8oV12USvmvbQ8nO6JFtne8yxSPG2SIBUYXIWMSrjKRVbozbhJZ+lqoT6
JsOGSpEQlHnc36S8QWNxJ8/Yp5vHirkZ5ZFx6M8Sb6CXsn0A8g0BUa4SzR2SxphmI34nvhFLJOvB
NJ0vrHWlNcgzP2IgleO65p1OK0EaUpB0kPqUeVwPYHClUQxipnZW36kSMi+W62Wc0zG+AEfcRcR1
tAcSAE4RS8fhbJId6AtWoZaCRGBLQ5/eQjbXpv3/BsKVF8T1YXHhV8QYTYXLhOG/TjXLsWpRU2WB
h75i5rnuMmPfZWm5WGgDzW+tm5mxk1UR2H/qbuPqJ/hqgOEEGS39dj3vV3pQ6jIdEuUsCYELMtdk
gpC6FsFVFdNKcO6vuJYkYz2Cw0sRl/h6fpzeM1a656c0rpW/siq7cYxu5Aw330+rHvh8fuE+9bH3
A/DA7uroRHPIoZbRqGJzuRnRJLPfHF+IpAudibcCdEyiKuLuolKrBofGq/E/69xtbdiX+icIJQDn
qDqCh/mXkXctwlPe9LhpimYNVsyeyom/jFlBEZzXr+5K6RCVEKR/ekvCFPJREiK5rykhCX+RqJ+g
v417dmnBRgNwIrX42SzjH6b/4y4wPgUOvCj9LLObbpy0jmr4qVbcBv1f4Cs5SwOo4qwe10U+82ez
JCKK9WLQaza5O8Atu8b2+BYu3D/uoL9MZ+TpamvZQqJRHvFgLEi2ean+bhe1GCDIaPn8CAglq43+
S31DPUz42zjvsIGA77M2WBeQFEuCLZ2dxkP+GMMnsfxnzRH1C/gkDpa4Avbja55GgyjSaZ/FFr6l
2C2iQH6ePywCKtbvP02KRhF8130c9RoG0OByCJA4NWDPwEXk6tLi/fQoDJNvnj5kmixMRxdPo3nR
fpuPHknxOccQZGDUROKVNLNe7oDRSdfab6NRwsyAV4ySi+5QeUhKmxCZUXWN0vR0y2cCr346/yI5
tWLxbT6ByS7rESBrWGtLEXeKqYKoCaWYoEIPrjMHIlJHHUiVVLPuf97v+D+A/HAGBYR2l+K/qQZ6
HznhbuJgpX4mzHswT0+Y1fp5BSlQ8Cf7BkikEoyMT2uJhgfETSPsk16hjahJqeYT8Uh5+8sWH1Eq
RvkwT7r5t1R6uf4aR+M3QBLcyfMnNiTN7ZhR0RLn3uBgzteqbxfR16p7gU7RPoFAyCFjWEnO86Dp
VGZul9cfxwU0Kb4rAejE9FtgIMCDe1nYrrgZyDe7DwhFkYdrXyTOFsn+q2ruHaxz2Ug4EokovsEg
vHJBARRaUOLpaEbrr8HAUnzYrJLRm0qpprkLIp76OlE+iiPQkjMGf/CyeQ0/5SLkNu9T3hQ9x71y
y/B9lrhT2qnogzU2E9f0NDPjIroSASv9S2QvZzaKJ+eQCcexBFdOXE/W/8RJQZaCWjKMwm3sSbbj
uYllw29KkpXB7WcRxSLmLka0BChcLgjBQs/vlEXMq0CrjDal+rFdWJN7mSgTVG4sLIhdiXV7wV5w
OslpA9Kcc8ZyF3TsiTRduBkUrFF8MLHLtxhCZn9QzYjLXVrEGRj1pvxH9vW8VEhNh8bQfrE+LN2V
wRr8JUkEIF7rtgtQm9WiEr9hmnUMU5NbfrgP1iIpMD4yhzwwybPcUTlJGdpAko63aEuj8KqH8Zhu
1cmwkc2y8O6x2lEHTxWewW1k9dikzxre3z3vkg5MAmELnYQL+pEGkIbiUFslZEoQ90TrU0MsXjub
oQzgcexVFIgd4KHMYl5ruFDJnci4wWkLILWiLUxEwHEwVHn9UlE0I+Q5v6rYsyc8x/hrxCa7LSC0
qIvyPycGSEYLdnKTptXnpYcL99Gxgd/JEDcHNH1aS+q3MsVHzzY0x/0Rp0AUfYLWvpqrJYY5LDXs
WRK0u903qSSNxWhkXMWW1iU3d2RVNqlyksAMTDN90eVDiykaug+wA0cNLs6ee+UcrFkUm1YQg1CG
iy+i7eBuE78XnF4xPymvReJQQsfKKWc/7JYXzN1/oOUdZyePOy7tctdaXISh8zLGSr6M2weGB0rK
x9eerK6cyVD9X5ecv97qMKfPt85mnwsy5DLi4i6yn2yS6v2ynM6AH2N6+8ZnegMdtx+/MSrJOy5G
oF0eEpAI+CcV7DKiJ6r/SBbfnAHA8fiimWMtT0hYU0wCa5tSjpB6BcMQ0o3YNDcRgvYtnov+ndM6
utFPOT20YdFaeu5+dyI7w8IrYsdVI9CR/v+EZ0ogmUse7x15pVG9/CVN08i28oH3WqV25LUKN1MX
vusm5tcVd5A+mrv5J0BLSrqZtAdAV5FU8Pgz91Gyu95ip59fT5ZzWqZAuHh3CBcCb3G6ePxnn3Dy
ig9RDwyJVbQ7cwFmFUC4XFQ0ZMUKV8WfMK6dQhsOI7L1hoZrKa+PZlUBhB8ICgg1k6kvQJkZ5rvO
yZG6IosZv0mhqJJTYKb3cmfpX7NPbhKBMHAF34pcoR7Kkf3595Yo9+1PnR9P2M6UlYAloXJjjhhN
zzSPX3YLZmR/adIMEmNJy1kRNQww7UpOWETuenJaLzfHpwRi5RimtQPgJfuUqczTFgnhD73uTsKM
nEEBHpFEhn9AHNNUaG4mxQ4fSP25Irs1Off2TJuBuOuUaf4iqDmGK4PkoiG7h/3HlaVvakx8ilo8
cks16j+n5ecXEi9WSfo1TZDO1ovh6U5xz+/+6kHfRbXhs9qfdygG4DrW6Dk/Eaolt2kop7LoLfd5
yInenABkEeTLqQY65Z1X82itD0P5Ihwt+Z1waeVaulnbHynswrbKWwaGi+nyn+M980wYb4BU/ZMp
oLqZx+Ut6sUzv6CjjAHzMHVcG/ZPFtorhAYPWcXIBFlSIIghd9wVjv7fElvMLfbRYfzlkRqeUuHa
Xr0RLZAt9HbacPXfYe2iARPMOSXmzHtCfPyf++WolcT1nOmkpKDv4xJnMqCNz4DNrPxvk2gD716M
IG2iWHft/knjP0XC05pHpLcv9K6o8i3W2bXIXcqf+YZORCRPmHGo39Znu8gl7kA3uXm1Q+C9rfEc
JhPQEK3M4dgc3CRd37GkgUFiGWA2FAMy+S0Y1pMbazJ8VMc683G1P4i5IRwcsHgMQuWQ9xxLCGNC
J35t55XsRsIusDstf3LWyx4DfTuXZAMb+C0L5zl5Yjkjmktn9B3vgfQ5CjSPws2nh8e14eE2z8N6
vh8frWEUE3kKHpIix/FaW5Bx3nlieZl4MC0LKsJX9Qo+3PACjil6et37H1JZ+g5JwlpfFBHALvk2
lvqQQ5eJQtktdS5sy7OqaW/LEqYy3Z1DEecn3f8O2ZiNruKqvaHIa70tDKMda0ajXvp60RIhJ/Lm
zBNOACzQY/MlHKMdAdq9INgNifJ+Vge/MEvftMFEeOEvK49pCJ84l8nUXOFoyCvsqW+Afnrlrqp+
vyRUVNghrcUCPUaYi2sL3r+zIanqeMACzcdMoNiTWqkHW5Ps2twRE8lBpuLZQstN9vO/bJ8rreyD
89prJUGuA5l0FBNmCqhQCymNfx01JX+HSrxiQ+XmZqzVduvp1OTwPHFxR1MMu+W1vNhZ2lTyd+u5
/5/6+yfqngxAPWW05Q2Pohdko9H2X28Djk1qNjEtftSEnowsobWfOgtjF+4B/ZKIg2TsDfCJqypL
c6bOZtUD9HnktNZ4HQy0EUYA1pGVPkQzsR7n8tuhETcTPB2W652yd0txt11+hlYUlVHE3zMtuBwI
nOWyVYY0fyGopQAweThTeZqx1CigYEPfnWMYJ0zGswaVza1sp/uU52/JuWfvK6HQ+UB1l19texZn
oh3A/wprm0XlWedfUYPEtztE79mxEX0VswU+WOUMfHBsYHJs/NngeyHZOLKFO669tEMVkuBvo0Tn
ebdX2aV/1whMu6w6EQi7IF5NUcfqHB9SkYoXec4ZzNrErCPh+lwwK5oBnbYoO3k/11pASDjMfAJO
8uqt0Olo7YPJJPvqpfxRhQ8opnwE8mBEF/81Y36FtUlei01hBnoCDuGukq+vN5hj+nwkYpQmnCrT
eyD3RW/cNbYb9KomVwk3ySqdPVJtSZ/wBDcV2BzbZNTBTH4kUET+ICyQhHgtb1e11Otp4wDNtASd
+5XEcbHmR0l2LZoEuJihWdeD71EVhMV7Ukx0EAifN4ItMfP8nwvksH10DBKMqBWs/vCZkQss/QqR
9rPE7rg7Q+X2RFt28xGhSY7VTa9HBZwYO+PSwSYiCOvRZRHkfMSX+D75AkxBwJ40c7wM9CytZbU0
OcmUxWBMKzwEu6+zJYXVN0t/8xZtyrRi+6HPdg3XCk8hlO6ZhWBCCl8AnJ81URbny+vbAY7gnz4r
4io5epx4wC9cqez6KccNiQlgCFwmVWcEtgWfSUfxjl7bHeIdIai5WALRt1gCHg6igdxJzIyhTROK
MpvFf4AmdijGnQgvFcxRQODRKhq1TS2KZ52t1Z15DNFG+SzKxHxUAh1IHm9qrwBX1Kpu+vZgKs2j
zffrMkZC9UoJUMpqAol4zWTWuzGj/8rG80/T1GktDxeZWWzRgVGRMxeq2knIQDPjzoMN91O+xX+H
QrQOL6nNvLXVHiA35P0TYiEAjkV1VmhkwKBA4zoFP0H57oG36A5ub84XknS670+GQK5HCOA90bF9
jcrOr8EkASC59FPUZjxCl0hXdbpa9LUh/QYxzQHk4+MJ1Djhq6SHw95hHLp+8tiiarKyKiBMbQP0
l+vcKEv8kurwEzjyS16f4Ep6TJwusAm8qIpUgqkts983zu/EiJ3nW1itx3QAeFKvvmcmTYszVPfb
IYtbzKqxmvJ0ZGgzq22CQClrjH6eiPt7eUJ8sxKH5v8lKXE+e/+MKe1cXks9cGWR1DjEFbffi/zf
CCeyawop0wfu/0Ni5nP8ZaC9vlizB9+wfylKviI92WYiDvIXOCl8/LKih8iGtzdsPTJrwnN+hOft
gf3Buc+0+dCO5jcTSggcdqk7alRtPwjlSrVK9qOxAIumuzoBXarSHRtrmJOjCZpa84gYBV/Lo4sn
SkoscqbIjMcq9qfsOp3iHmNesPrJu6S4yKNnv4G/LDbthsQnaDYZr2it6avERlyGTxNSiM77Eslu
SNN2YMMkYkvWJ7/rWjfn/QFD1mufFmXaCPvhtLgw250qL+GTVWwVWX+idTW8OAj975IlVKEG9tj5
y2Tu6zYbNZVRyTa3SZSjkUGnH/JaYLzujWJjA34s3XHgIoA2VdDW7AylKgsTS6n8sFm+FOhn3Pu2
a4adYqxmESEqglF4TavXtIEeqv8k94GiWbWPJxaFGPKqdD5qSZftTQ+7ot884LDBOXW67HtsvqgV
5bbRKMIWITGC+UkKubugxbgbwciKueysmpDa3n5xYUi+Nq4ndLGVMWVVxZbqyMftLhK5lalNXTHY
eyb27Xi9gA5V71gRhzNdgnHXQPJ3MRXjfKwy9xUGWCylvdnuDk1x+GMHnzOsuD5ifvurj0gQqb53
ZpHgRRySR2B9ASd13pE6RtcZjBMNapHEAwhDpEO/E/Oc2X/vo9kGmxBT0sDRbTL5FvnEOdt1+98m
1DRSwSDgLjvGDuc0aOKHG8rUwHJjnGAoaVBcC98l1wIJu+WVJI9YgAKaZzsnDInQt46uS7AkUNtx
UHbRpcRsnhnsq0i6aNuKwUPSB4wmM7LOhELWYPh6OjyWqs+T5hYbAv3MnHVobJ98qGSHMwr7iwe+
JsxifLT1NMMIchnETBzNBFAHvZ0tCSYCMt+gWflcdFRmPgUf/X5k+6v/AyuL434VJRk94Q5A0jC0
f2Vva8RJUu0vEkZ9iZM826ZG5CFZ9R6Nb6BKXN22qmGJNhwg9yGJI5cPfQ08SRLgr1kEK4t2+v3Q
39SJHsn240CvBWScMElSqKtYwzF6Flt033SHESwt98VUsA73kjXCPucETfWWeIJCjGfgk/uqTH5r
D+wa82G5bjY4dKFNIp0D0weKYnEl+cXzAWQPQtuaFgWlegNhL38e8/DayVZEWsKwBWpy5n6EbbVg
iPJuhMr8EMesDrHfkIuu7T+RLMXu0IwrOtsnullDUvFd0OTRDLy22At8bpUgP+ov1QZQpIrlQJ5/
szTs5vVPigPnrZRU9TODFVVADkOajVHcmM/nrug0ByNlbqFzhu2kIgH/2U5AK8/T1XvwBXznm4YZ
x6gK+KKHk42y0MnKcECyKAqPSRxO1kls/YzxU1bhPysqp+rrAolXLlcpxYOBUO9H4dGciuWJe+cX
8sZlZuDqtRXyktbr5BC47Or5ynXbV3BbMPgk96GrM4RCUBXClHzznO4IOqMxuU9GXAP58GZTY1wp
OCOThoJL7pKvwtHVRnjFaa4kW5QbzwLDetd/rPzGmrWyBt8Taz0xD9nJ3kppb7r7MLQDTY8HX0Ty
4ekzlyY09YgnZyLgmLG48R+wQbINhHuwvyPtJRGcaKFEPwjy866Jvjrnk+toAzOwOjurZjH2DtEF
aMQL9IM4tJbjbepAgj5VSj7FLue8P9lYbng2l6l3fW0PFWonAUmubHt9gYTlxqbIO7jQzokvVvw+
Uh+FdiVwLqDFfpSHSA47ccMexrprQEbIiSGGJ/WYL13G7oMDg92YyPirEG1dnO3AdhYDZSc/rPmv
+2JfoOERlfoCeLmjTszPD+ESCleOifcZ2ONdgrhcJs/hhNcfAt4mixQZl08Vb9pxP+WE27fIdi5l
9EAPNcw5qaTBxnkgOtITJqa7wynOtODpDGTNssM0a2r1j6mmOU+bwIYt+X6l0r8msVCoNvGyDosW
+eU9ts+qAf8bHg/acQXVvN1vVcSed05J67fWMweVZj6gVjdh1PYP6SKwjEu7qqtURiYOfR6A82RK
3Zmn0UiK+nMDz+gwvgLN0yDOCJ1iWm0optCLYdUqV5cBc9NhtlECEuUvCLDGSugpTaJbSg26mal4
zkZq6AgQCrhlB7xFYVzg/HfbybFIcQJvR1zOJF23kPJd4XGcH59UsSXpDXL50aTSOtVVVug68H23
K49wCOhJqP23cbuYlDD+32TV+/JktRFa8H3426bQmv98+PJZqh3lEvBg+YiIRzFfx/3k99LN0za6
oe7mKssGglTHUhkB4pWHYSlJO3O1V9QMBJ82E/H3YIR/yA5LSebTodv129x9wFSeuArg6fuBstIb
LDmuCJn+taAhvXK9Z+N697dwzk5mfWOWr72JssHb5t5Hf8akxuP7KAAg27P9V5IjYqpUk5djbd0P
kIj/rSEZUt1CJMHJTsG/H5Bowifs0sEaszoh8gTDjhmQbabkRTs+zhS2tb/3KYEYHENnyU7JQ6al
d1nBCS9ZLJj0pE2tJzYb93jK6dape8K0SvK6gPRcFFKgDvClUeLws6Sa9USWLIa4SS2fGvnI5QeO
h3uQueFI0fQUDI8HXIQ9rpwrxNMw6tmZIStq2AeU6C6mIlMTZ6QIRW/BsNm/XbXq5j7X3Sf+wB64
TF6wAoHvBR3yY72kF/nQT4YD77mFbYSFYYmc4NAUwhjGEdibHjDdYQRaccLLsuEFuiapUCUTCACC
l5AQeAHGk3cwcPUHlhDzp9SPDO97xEORnLjW0Dfr1b2LnQKLJyath38/34cx5FZUocSNkyWAuWal
0t6YC2Fic93blB2+iezpRW/JHnKR0djmV33JC0s/QE3V1FD2upMqvLFMluQSk8IyrRi85YmAj7DN
c6M6ezqmm063BVwXhsqQ/PxO1fYaAzQRNwBrC9gDOYqs6ud80uTjN568EVQEGaNftHGVdAQ64s5Q
sU6006DHNEwc+SxaR2LnA6ZcFbFLcQtUeCSzFI6Eh9lNXGG7OJNfLucKgKWiNOm2FkD49OI8gaRz
uedBDJ1ZcBQeI9NtvaLO8TFgXw1KS+FWmuJymtKIpI1bo1gg+NieFSwbDpYsaS+H/F5J3WQPGiy1
e4cdR5xNPnDLd+77bBIC71dj6/FmHPytRfPjsZmKAH6eLtp2F80XrjSVOLGc1pZxjP3B/aDM8vwE
5IgHJBAH9NyQCqrcgN0/+5EcH1MQKhw+k3TElx15sQfMk6C6q/dX4q1/btJG/84TCaXzdkzQyfLU
LrXkjuaEbhB2Zga4+Exz+KvWCKuiko9CVp6szufvtmUFQpf6Iefq7uOr7HxbwgbrDGmtsxfZ5owf
KmuZtZmgk2YDstE8Bo1iOx0pAC3JjEY8qKXzIkiqNQ9W9aFXPQH+SLh5xaLXygzrU6kP+LaW1NEu
u2jOaNWk+3VcBE4rWoEUHpmM7mntWyvFTb2Nfce0FZ5ghShddTvINKWUAopNZzVuTlHLAZZXYu/y
lAnXpRGjkHkV36gf4qFRnbO4j4VqX1QbRS5zyZTOoAPgpLvoHq6bqK6kjjekG5xm1Jf2R6wCcM46
6KBKu47WqD75gVMGmyjkYnslX2kF9HqwPnTbBby+HBaq4OMzad6dMGbL8HNr4+Lh2/Xd8hsbO4uG
yBdT/ZH5p5ZA5GiLApNJwda+Fo0EMLL5P+dC9NdjwHbF/l3tp0TCIkD6LpVdSaAUqbkGNO8o87PY
xcY6jmwBNM4HqdSuULC8nLpG/xdFVjTu/PbvUY42Bro3qXQh2YZIcaJcP0IdEtTLvNVbOpnNsuXA
Oa/ltLqtSlSRGg3lX7bSAvxsEIAWSMz9ir0azjOLeQOpz3OxTy1Z9VxpcqQDQD/UFaXBmJYRAeHJ
vQ+mUIgnEa1I55AReiF758f1gbSGk7G4LUWlVd7FwT9DF8mKdtwCGXY6u+w77c0WNQP3m5xc1Crd
NOCBOUkaazpkQnxOet5p3zHJ0R3T0wIR0mHh72LMuVVZ25OhTL98Kv59IgwR/Q3McsbRZiQs9AVQ
YwvX9Y5O4k8pY2TDRXsETnkv1w6L2WZlxZYjg6jYSbDVq2l26e/x+zz90zMpTNjyQY26Vu7QNJyZ
k5IS8eE5r6GAWlVDsmlS1xEI+eOqfxzFxcqflyVkGQT29x1SqUzHVyZB7AOO8llC0CvrBFeXwsZV
Bzvc/v+jRHHh5RdZ2lrT9DXUMfup7E5zX8cNRVjhkMLaAMtiX87UQ1CA8mFWA38r2VoeTuLCpIGO
rMCxbEEgaIgiY5SGoaNXCi91qMGaWLd+Fn2CIcRc9bRp0Yy4GWYMeWcQXQM0j1m2xGqHRhRIp+Kh
sTDOVFX9gA69xaADGC1W2fm72hFAW4QJd8e+tzmTO/yyL9Dc4qS5VbldagXZlKbHxFwAfxJgdZ0w
lnAjhEIo2eYk/8XzD3TNXVzRMndT85h0RVjHPIX7V3TmKJJTMU9581x+OLpYo8xZHS7i0RUww4jL
vmgSbmCG5vKDpaPaLbiAKaKp8sfp7GctZ749r/5RZ8c1+/lQtZJGYoZJWboQLw0nGhfV8FgebNr6
ey4eGc8UXMc9ZsWwbpYs/MX5OlGdba0OBRuzpACXgAyZFtcgtM2VEeF+HlWE8ZTLepQIhHMTEPp1
W1F+zZMKgIsCsPYOf+lZS0+dZ8PB/uKhggpR7VGRLgLRqZqcdxRHY/HavcxJXlkf1IFf/Hw9qm8r
ADaBfvBvt+ogrCwbqinPAlLQfHnp4RMEJZcSM77dP6nVQfJ/VdM+WxBC7f84SRxAtBwOaCySQyP6
VixPgc+6jwguegrrDn5eTP0mSi6+qGcBGqFr9CbooXZMc9LViBxYFvvuMPjv0OtWyznqbpQXJhKd
Be1uE/Ya3j+vWtof2BO0Xm5nQGY7sFX5g+zKaXeV1yuLtZP88alKuA//bFu0SezKgJ6OhXJuXrBc
N5y+c8Ij8GAYEsx2HvpR62sP1PnmEIy4ZB7p/xWKNKpIbZDaoiLfgeMAqk56gFBywSkxzeY4r6cS
sRxZYjIZMdGpW0Qa+l6BjRKaXAIhR7m98klb2fiik+St7IQbKjCqjiRd5JRVoW3Jjm6QPEbYm83m
fktNUeCmSj26+VpHtDWnJe9N1d82tIrx56hddmkQnSIDPqEt/LhTIvS77EuUsKCV8+9gEpuuBvu/
OHGLkLVPA1km3Gqdez/HTo5flBhwZtaMHa7eu/3IhFbskpsZ7dSCfxBSNJqB+vah/48Djhvvt9EE
Xrowpu+cp276MI1frh+MSLumV3CVs6oXteR29+gZ96/BQORZSxbMTW4Um0HvR3LzMmlLI5ERZ3rI
g3/sW2AMQ+U/oqJa6962wMOpdjIsZdm81iUbVrbdz+BT4czzbgRbLfR/vPOIDvoE5XZLI1ZWscSi
iCwO0cny2UKowkAVCpdnckPFR6YfaHWMusInWyEWkvH2gvJT0ZfJLO8V2QIcz5zeR+LH7I1h/FTK
vBG/2YHT25yjrOaYpyVyWsu4HgszCwd6VtjeH84Xr/b73kg/WPu//N0vZyt4iK1q3twMXOOUVi4T
rh79dcWHzKfBg1LVUcNVYbQgLVJr9ofZT6dXEZaGiw6A+Iugpm3i+pzvtOZeOsudOuNhFWX2RA6O
4wzKFmCDI/KMObbIkCIBCPB+jt4kJM34uqnIvOMdzlckAeDVnZjjxDdvLcvj69hHzQrp5PXl0WiA
VVu1Wbj3NHcpvuh7uxH2A3HgOyBlRvomE63k0LvbWKdRI4ruJcF8rseJxhO9TkmuxOo+HjEfbmVv
1uwHJGPgRoIj5vvzWo9K/jafK9kOMgjPsaAYxnrG9FTj5f+INSWlE1BSmKQOXm5f/cgxRVLSp/CO
AfUpZU9nEYRSFjuAYJcFKMC6W9fIKoP3yeplISQA7ShOt3fWC51D28LnLE0WRKIYRsyr75+cJX6g
PNAtzkZ14t3X0/vD+pLkUhZ+h3a5HxkQ1zcSGuRuxswgHLZdY6+JE0TLfQF4khKB6VoY7OtKigoJ
yF5LfNdAqVI5icC87u+anQBfpu3XcMjve0UpokXwQ6Zdd8YFVihZE+gtKHcfp/wr6MZ3FtUYE1YA
WGQHdKQw7nEh252i633k0PE3psLhnrZsnPh5yvvcBLnzMZcRZ9gkCDVmQXDqsXEP2qO3NgUeGsFT
Sw7zUvftUDoIjUEtuI1JHvCCXDvTaYl4+V8X3LodaOJZAZQFKSdq9H5qh+8lkqAmm6vKi0O/Cear
fFGFLjGXcz2u+mQOVb5oXmhq/E9YNZrZ8u+q9TUaWSLK/328ckwdWH04PRdRzZ5neDrM1vTrSDH1
SWtz7wGTBHUOvuvms78GEt17hsqbC9JIualwFLq4l908WskmQPSJ3SKHOPbUqsgpgsCA5nwZDMzX
K1H8oGGl81s96Mt+FSHXutcSh6yPcYijQQ98jdMYNduDOpmkPz84wfDo5VQNnksX2pZdHp9LW3d8
dpRRYeLoZpBlQ0nhIUEZDH9925fSzuOitOfIitPRy1drYLtLR3PBbC1QvHjBLDYp9D44vDa6SfXy
jJMv2zI/zNezzmCXvfgOXd75fhwPdVgaPSBwH7ETwmoMdQAKVWV7gYq2YdcCPTTVwgALDM6yjDcX
kWodN8vp+8VyOlUzOnA2DccWopS3RWYu1MT+GAQnxZSZmgjEizrS6yuXMdPE4YLsAXK6j26PyLkl
giKxXhSWDmlWXAhewh1V1pqY+MOkYMzc/nwU3NGZxwBK5gN8shdoHotfBTdQXRMb3xj8yoEPQouN
Rf8qfhfkSb7Dn4RO0Hadnx439+YRLwrDSsvR3JmO7yEjDVgro6LNA50mA2Y6Gwiphd2knMGVbvBs
mWY0oTCejAzn/S0rgirJjdwN6pFWpRC5fTv2PicX7imbgZxQuQhXfeLdlEQqKoW8o2ekmoBuEb0E
LDepEwHSueIlvlNGUeyKnsvUrZ5XkEkD9j8HyDBw+8WihiYw+Q/fTQAk2D8wlFLSKt5iK9bDI6Lo
iOArQrTJFs2VRCPcFXZkmxHV5aNCfGjmbIao5oBwxATX9tbVdmAYzMDOFZo/2yxPAweZCtjbqpxS
8qt4DYgBSpLVMt+3GEq+nM+j1Y5ZGp9491z5pDokIk+df1o4CF58fHQYpSaC/iJv4vYLLvUd+QdT
utsQKfNvbiHLaxneeUmeY1foxn5aKAEUCWpDk8N0yVg+a1dGftm8bit3QFJDth0e/ecPLm6XCSEY
Ef8+O6P4UZOpXTMWKwqwJYE3KBkUsYFjs6WMAcbA6jAJp3rkghz5dWR+Y60Qvi2bDXqsu6do5XSM
yx5HjdorwBbg30HMW/ZcPwqEreK9YPUmfDcz5aPcBNcjrxLLp4rAN03oQ+Cg/8s52pw4FVkmhYaN
LlA4DoY49/qncl3Di4o4O3BPxPQhB90rACEJihIXFB7rDC5COBrl9V/i+1o4HEQr3U3Jt3c0MBgg
f+yXmhbIKUUOFxxA3LbE17Zs50+YPRSbi/h1fZl6NkqcP7sJ3l9iiYDrs2iCil0jLd7OlyaoYIdN
LIM5wOHD50KPJOSg9N2U87bQil3pZjY+kWGJytvfm96pUJ00lTKBxe5+NLMTPRymg2K4kE06OfTb
RJLEDU6AUjaJROiALC35ZxHLqy96gjNgcdsUEK2EtLVB/B3DogscLaSMnomB/QGg231Upmn+SHLI
SsjDhach7x0cL0j8KfnXrhsU8an5GO4dX7dNX7EQpeI+2TrNFK9I4v0P6vNby1losw4cRaUJxFP2
107q2yOlj511gHHLuH+aeW+6yXSTzmRJ5iyYVSBctBdT6zkx9NMn9EDkTrNe00p8gvl6Y6dz5OaX
pTfWW7cpcFlASzJpEGRrsuZS2vjsCl9cB7iD1Gbl9a0Okf+eNTEyz9wFVrPBvejU1i4E0k8pHsv0
6l9W+RF6qEo5jCItb4i15YC6N8NYeKyJska4QT24Ke8ocPmt6xoxUbFYbSmXUOkyrDs2p9yDTWkI
5apOil9roP+WW5jVrQ6pPK3OeJXbez6zaM4vTlobs7hSt0oTDMK1geF7/Pv86m/PRQOMvV61zeb5
6k18H2bz4fxGkXa+bhiaZHy9bbDVKTr3jsFiKM3hLPOKvldeul0nbh6JBSrE7+bQCrFNGC+7eJbr
HDUXJ+QXfcIbxpYBg2oZBKbwkTaRJDXDYdgGQQp4lV04P/acr8YRA1m2Dej4ybF3t9XZQDvZn+O+
h5+Hr3SgDQ5G68vctu5yoqsfAH4fnRvwt7060Q22GO3bI3OQhEZp1wu4RosvkGf7pGvRqPON40a/
EYJx8zEdMWbGJaLs/1AGo5yUB+3wmyaF6NgnccB2rtzk4xjkX3519Sgy8CzJcQeJzSaAQIvMn6OB
mfBLeteNUk+bmfJsjpZY/wmgZJ8EGFTnDlmF6yNfqIHOBt+C309cZYNPimVFsXZR45OBAO5Babny
EwWl3FIAYCYaFIXyZq8IsDCIiL2QS6cKMas4Cxa2A1blDcwrEWq16D69fE+3TWDixeMAZhfQNVEn
tmIqJDXBqPKxPurm1dLy0GvWy4OZxc1Y55iB35eb80eeYSFRFFo8In7yvw3sLbbl5n8UKzpDGkpV
rIFAr170Tx4gOJJzQvxmcNDmuLqR6/NVNC4Qfa5Bs9YAd/5JfOcpIKKJ+pATOvR2RML63/q+771J
gL8WqEeHSHAcaSf1Ns5ZALe28yWendltIbkM/dXXWwUzAIU32rHTVKLtMJJxMP+gK2E142o7lBdB
f4fclGU2HL5ckW8luqn37o+M7HHYDHa/G4wFCFrjyVAlmKBvlSDS/RQMZl3d2CNnVAsCp/ju/f48
2CiL8j8aXL1ShpLhgx2iuxK4/6rRkk+y2Q5JjGYZmRFDpvsekQZArWIJ/b746C0iQgn6OEv1GPPg
vykDUbuArn2UejDhgQfpxEveBN3aAGZogJ++JNkOs9BZmPGcqBVnDty7gRACkno32crLvl8oiUzK
EsTUN6FhnQSzMpxLcRDRJWGp7DQQpUp6JiCcKbLHDfW4ASGNjWMhHBPOMFE4Nv0OCIqPyozajbuY
iMTMaukTI3TUP5umq7V9kc2tTkCJKfnCWOq2j07ZnCS2KXXcSoomNDriWepHuUiaGpfs3D7I3QVi
McTsV3Vzb2h3TVnCptWhVGdYeb9Ikcts8Og84XH4BfOC2RE6DfBZRS3CCp9W97iNlUnn65d1snlD
trhPKifl3ILPcUMgPChewQycJe9cmumed447RP1ndNHoNTp84MzW/Y5JhsQYF8PuSaRL+D/qRZYi
HSquw+B5nwye3WPB4R+ugXXP9DlcY2hF0yXtdzWwclY/kCzkPbPFElAm5+k4ralR9uHJp0EpXvaY
z1HmdTrh5MKwJ7Un5VqdaczryE64UAwHqXvJ45c1ZvUYQmV2DblLdPYPOiPgVxrJLa+osNcSSGbm
ZpMWqt9UP1N0LAEZQzvYX0J6gFEOl7H1y9cplsP6b0vCikvolZ8Hc40jPteQge6kuedShMXqQAav
IZsbWUYpahOmFbOjoIfmo2+6qZql2Gj00VmYD+8PspUV2hwic7sGARp06P/PT6rKrfrPwls8yhBr
1hmvlMF+xkRGkPC6hV6o9nzjba+ITY7NkRokZb2K0SDTSccmNAY9u3YP3lc6QXdERBm2DbdmHhRq
vRLQYheA/k5vUlz9qo2iUWlgFYyOrBdr/H8VDHy8rq/+tfznZX8IUBDlYfxNC2DHhPaBynomGelN
ov4ONP9B/NfAghM3Z/htIAbfA7rw47PEBCqb9A0EV86rFpeULbvLYbZGxxsYGyR5HOwRfJIDZtcZ
Qz0/yF73yQQYSW/wmE4MnT17qbe4rXBbJlcm8wbqmACxylpoQY+Tu/8vyKhndBjtx5XSBiQAiq2r
JKnmZPxCqwmC/uG+IrJLUOEDuhLBuXMI19gRM2RaBTaKWV8aM92A1VDePzCo/MYccwaEiKrnHsdi
cmObHD6WvIGOANR0eZKv5rJWZ3sjB+yTbd3X57G9VLPJ734qsPVQSIxKnTUXe6WM3RCraVNFi8d9
1PF+bm5zjHcsc68uYBM1haiuE2sCCw550ZoMytRsybdISnYMolqKDfSxUvgSzvQPP7O+PrKWASsf
hWhfK0ebvRiKWd1u7J843AYphya3VvUvk/vq3wYav/+UDGX5W/HXTlmJDc2eCbezjYJ3xWWq6zbA
gYtZfuhQnDvsro4Z+ZMwv34KaViI2Av8st9z6Za/DjenaWlJO0Zzd6Wx6pVbVyJwbs5TvkBgmKQ4
y6r18EIzOJylb+TybCjJR9zeCAsqwygunPcs9bM2nbhGy0q5AEHiJ1zq/7SJubOmVk4Mj3mL6fp3
A+KVu9JS2N+TRuIx61LCgvTvEhh8XAYO/w2Tigcg3udgl496jgZv7KbyfrH3mtr3z8G5vGBEj2gZ
ux03+aSe8bz5YSu2goqECfHDkkrLVMT0HstkNDRi7SWIbrD/fViX6HqK/RBl1i4RPYE41PveUGx2
KJCQi3wQxwuRD+fV81lvGGY1okzFOrhsuXHL5NMDliUTSU0G6QNIzFSRvytZyfy0aIlMEWvCLksY
K96DqFKE4EbOpRdlcHE7em3YxBKqFOzdP7XADR+SR/9XjnEtGDPC6UFTWMplsy2OiHhG7xwPlEJL
PP5Y0rPM0SMnCbC2u9/o63vNEjwxaX783YEeofCc5u2m8soUFx51hCSJrzBNOGHSHuLps5xETg0S
g51Pi96cJYfXRYsh7yopSj7Ey5gLomPTj0eWvw7EadVjXdyKmjTIMiHnQ9tedCWwXyHXUIEI4XoA
X9K8PhxON/lWEq6SDlcOgUiuknCkREocT8Q/P0dWKpVCwHv8E7BUxxw4NjMhGYVq4bG+ZC106dBi
lrSp/0NhVrsEPtKgeP6Vkugg8Rg/ZzdPyBxSTYuM3qt+ZCsTeLJS3IG+FC8IHhte3AyAbGsuLxuQ
bNJ6oJfxzyIHZhAc8Z8sIqAbvD61mTxOVCi0M47EKy3T8cgMlLQUU+HWRDCTQNQElcSGw9b4HbUf
TW1OvcD1krrBfuB2HCu32kdcr5Onw+Zd1DBfKTWi/Fjup8AAGfmNN7JHuDZ/ldEbV0lr7NVIbRSe
Fvcp9ixOrTdMRZ8g+4EKyy3cP6GOltnlueU9VV9/xvn4je+EHnjdOOutySDOiyeJN7oilsSEf8dZ
4yoxrQET6Cl4QlVrzqwUFW9QObHQFDEkt4X3Dteu9stfa3+Uo+CPYEKu35vTkkk9pl0H0tOmsX4F
KGt4kkEGt25LbyMD8M2gxXWDja8PSHdI5FmLC5xHXvUB7Tb/TCMtlEQJtv1l19f/ZHG6+s20Dbl9
3XV8pLhZXA1+waZGVXRocZrxnqnX4qnhMavd64wAsYLHbSND5R9p/OUnrrlbUae3GFfAp65LGsYG
1lDwDQNcdKjTvG560cZuAVPaSuevNsCPU48U5OYHY6R6+Dsi3e/iz7CTpkIy//+/QTpJoOMElOct
6yS2Ad8X1CcLRvWglS+Iy7jR6KqwBl7UiuhjNRhw9OtEWCJKs8B3scT0X30PdsZa48sOFoixPCu+
TIbO1sd9PEDwg1kag8/XnKBHzGYk3HkMok5bnjvnjmTFAFxECBxlqEmJDdmdyvg/cUOSh8TeICzQ
2DV/9XhsBOrKbid94PDj3HVUyDVpYsW+FFrawUVTdM7aEln/3LLK2nGXvJ1Ajf4NOZqg4gCjAht0
IkT9fL6cKW9paYFAG9t6Me67m16YouoGFnTYfze5g/87bUk2e+Ig8yg0TFdH1LwVXmkBkIpgGdRC
ALGyKFUX66+i5umMQ0tv5A9do+gGMt7m7yoP2Kluq5r/2vSxXUpOwVr+iOrkN7ZKqmgbS1kAsZ+O
u7sDen02lz/QJmxYpuznvqyJn4FBhPEv0z+tATOI2A/0eukmNyGqM8XepZgLya7+tofmHYJyrhVu
ennvIBwfwl+JHfEe0yxEKPDJegEX3vwoobr7GfI8auxoKuFZdsUD1gYaSHZQO/OXbd4/r0iG9t7W
afcZoEltjKSsI47y6sMHu5AFuELRMQ4qvNUxA5E8JvFG/n1RWxQ8WQI0kifEqKPa9D5NgPLG36BV
3ZuAfuF1+JSPvd2ciVhzu57IzOqSKfO/+UPLXaH10TGFdQLOPzY7fmu/W5QIp8t3s+yjDRxP+3Pr
AqTZLkuGR7n2qlyYHwOnmmGKzkCYWW8NN/io8jeF51xJRO68VS93dAzKkPpwEOJTHRb0rkiuN01w
omNOIfFoelsbTT/zq8CkmOmMbl/jFAnpNxM2Q5VQL0dlkHCamjdzsqE6NoX5zL3xF+zoK4Xp3XuZ
2mTvQkecPZLrch0anM0lE8yHE5HpR66BrrpfblJ1rlvybBzr2hRKXBZMVDMZZ9C4dkqEG2lAxi7Z
UmTWxVHrud3BcBYUp1qdA8NyH+fvWUbv+afXRLTaR43E2MhIpPTNGJDErNasGh4QwY3I1kivEdmB
T+/d4SuKr0TzUsX9UDlywNyQevzXt7hw2ZWNd93o7MioWOzARfaBBNJwIA2pcNcEdpBcbdNMbvjz
19ZKcANuV9Fc0sMVhuIvxuoXrbeN/XkNzRGpyK9/78Z9SvPuTlhxFBYUffF8wp6kiV8jPCM2NwYP
biMDXV7O3yn/tMiNPdZyyDPbKCoZ5vfic5E0ji0kNBlPmf28+kDrGdSfYVwbjwVVQEi5wDrgtsWf
pSnkjqiobzWK0gID/vWgPYt92wtmmvwjqiq3pVRyNmCb6B6TY+m9QqNOiVE+dUnPSH8royuPsb7o
b2UxqAYyMnzGlBat4tfwPaDbsk/JR1JrXakImaKPXp8waIZl5lc23K4Ktme8ITn0bncybTLlXd6l
ey2TSIEHS6yeREWXqGUh09aSbkezQLxhfh8aJdS+8QGymryAelL2bVC9I1PMVVcaSCkLOAybG/WE
8w23oh4w8JgOggGAh2PJ7IA2yjKVJAdY4FdZjImoRbrVzNs3crr5bgkcwx5M1aopa5VXB0npwCNt
ByAaDe+oTNPCc9CLl/A6T/sgvYVZ7m6+UbDiwfzlF4/JJkmYS3v9Jh7Kq2VjKD4D9ttDQiA1n5Fj
cZSB0bOhm+wehPj8c2sKWs6d0ktEftkWtUzYpoz+RmRzBYvbOsuKa+sxs4SfIbt5Az6E571ZRhbS
RrMdDEjFP9eFkTHvEHB5EG6BHJ/MVBKYjvxstOxOEyKqw8oO44zCmvXZk4Mqkkoztjd0Xe50igwb
7kcM2m8xIipUCcYKJw5XlQIYMmTHHEWQeNZR3KiSiH6ElKbkPh3oDilHeED94htsxMSNF8cSbhaZ
ZwtCn4rjGH0zFHV/A7/DLCko7ku/va8LlDTVqVsx2HgISxMKqJTFrhlWavqn9MS11jN1pDIXavgJ
xfumgQXtUsrzqRv3cMxFCHOLZwNQwu1vCsYt0/G/TzzURxkvzQPQnrQrEDuP54kzLuaj+YDjwLA6
cDaAKMq9ftcNUmd3ZVisFFrvHC1VRNPzR8WGRZu+SoFzkZZb2N3wb+MuEYWFS4RyAFghakSIRBFg
KA5EQgvNcG6Ffw2IPE9yuT1V7HLsTpf31j17L2p1Xp7UaaSzl0TbLiPdEIOjjw6vviH4uuRGo9wk
ZjCPGsXxIz8TcG+mzp5Ap7QCd/vh1TrRjLGwBsFPSsTcFGzhIeD8oesYaygAF3GLMr+u6YZ6zsr2
s5T4xKY0uzkn818QnFWHROQBEGtTYRS4IY/UY72IhfJ+Qqpis7UBMmfQWlNQe/a3RbjStX/fUCuA
2QpmcQ+gwY/dQi8Tz3eNjDddT0NHEhVglEZayWFUd1dBCfhaeYmKjggdkQuCDytGLtLdRo5TcoWU
AUoehqfwAI41++XDxZKs3E7cX471Ptg8hi9MvyRhIMD3yfu0rIfpgNs1dM/YUrjCTRJ3+kof46Zl
wL2hvP+aIbtC9nALJtQx4IoJc4vdeA7h2A1a7m7UFAi02oHGCOtTEF8HgWhTgTc2lQMJNrfoBLuW
rYNkJwvPKOBxhsKiTMFgY0jzYp5aoNQQZr/1ywgBP3+4bOrCojMboIP7N7CbcIfgSgkb1SsxXVlq
PIy9rDcP02TiqtJ0H/RuD1EBgG2vEybSUzj3Cx04Mkq5ooJmLPBv8P+RVcovWb/TtAxIwwbE8HzF
9Ibb7e4Mv9CbbaJz625oJ7iVrt35LHYFtxFhb6H9o5xy0rBSOUeOQJqC1ygR/Ct4A2tXUuaCzPmw
rcNgU+k4hlPNPvfN6uO9ZxHWyTNSMbW5BAJ+tuLm/xhhYL5y/SOg77X0EawkX4SNsUNH8qatA1Ka
B00cWq8kYwJd1dgZ007EDguv3KO1L2ypj07nhMLnHG+tpo8s8Q8i/uV1Zym9WO507i18EMZfB82u
PkJorteWYrmqEfY/SVsagDWZMEN/r5nj6jHTUEuYWrAeuY3d5rbtV64rUukDtbz1a6Padf3TrL/G
vRof5ZLjLor6NInfiFPCoIWXw52kJ/zBQfhE/elwUxZShmT1Jq/O7ek0G0iuLAV+/gyBq0lorRSy
fRxJFMIqjbNldjZ5yxfRYwQQXTLydYVzMHVKX5J4PprVg6AND+4b6nATgSB9BKF7wqXfyxXWbUe5
YUEY1OZzvqCrSeDiFJP5H+81DKyFLxx9a5zCu5qCBTCQn6o6bKtWKuHiiGPijhpA6JVpI1xiKtn/
XiWXaVJbguCunwDpuhWHDtkxN/EQnQ6pc8vzQh2fqoF63Ct9P/binskYkohfBFNE7VXwBecTHDPW
km6XNA2IGOZcK88cYhdktowP/5E1gsNsa5mX2xke4nJNkah0Za8Rgi+jHgj6uLd194cQmUXWwyaw
6T+imggB9+C22CSnsPs142AwILKq1jHk3uXDDqlQVqkM1gK2m0DbLhOZFsI721xULuI8H/hKUavU
UDfK7c5NW98bJE1evyXO0jfdUWGS1VKARDwMFyDpS/L/RNYugOhGby9AAXwkNxybcsO2bU043N3M
1tMb9w95dODlQD+P+Te4RuR+6ywFw7Bl2p1bP5XpMWKndpkS/MhQjOX65VUOpWPciSSHTyVklfvr
fQ9wttgFQ23N2Tw79oneqy/5OGbKvwuuEoYbZXdnoNj4E4n84upuKHVmLgx93XIvN/zWzvCqVxwW
ujcHOb3Stwmua86+fo3dSdU3RW0241npBUlJYgAhkgmP4jQkk8cOATwSCaRunZBY+9GbMobeV03h
SZUzhnxa8vPHxwCngawuMbhKreqcMKfeeb8Pa6Zui0kRKnpWMGUbso4N9v6nV7eAELzDvtiXO8aT
5xIUHhtpWXg4M4fr+29hQf8lgit3O1Sbn6JFO5iCxsAWYqHI1Z69h68fTbUjZEjAAFW/rB2w3G4U
KGl5LMg9zHaV9Zoibr3+E7anvK87NwVQAY3WH5O9rfR+czUFcVTEr6fg/ozWxvSo5imvHxK19rKY
boWelF2vOraWSnw9eqNmizdKXojDaD0Lo5E464qxT7NTG+0K05GyL+640NsrPd8ap9G/V3a63oji
xqhvzwOVzr+EbvG7of9ss75PuX2DfAKkk6uZMRrhP8Ykpb3lUGhtWMTQJo8toGVKORZv2vw9I+7D
N+lafeWndv1IkPrikjmFnL5sHORTvly7y2hh27ot6vvZ/vozrCohV186tqIRQwqwaDGzePX7SEvu
THtbo8leXoG0+9biZ3dL8SL8TGiAsYGfaiScyG99uv7D55qjXdF0DIGqjdUANs2tom1IseyHW3Af
m7qrBqtHEqS1vCsPdaxkReku/NS2Rkut6xDgX0cU99mIFn8efhK62ry6+d8hlzRDHhw90m7FuJ95
rpXOWJrGjtVV3s6zzSJ4iDzokh9KkX6IsQHNcsFMbWbXlo2i7c2WhxzTRGKwm4D1MF2yV/9aotjn
fD/HAQaCvwGdYFCkcdHVV/4C9f5WE0Ru0+iMaGmcYn/Uk9SooT9QV9yFiAxXrmZ3nreIY/3RFCoy
NEWKrgqlgEP033r5QAlZOiuTfX9P4Fa3hzMMhGnncgyg8ZPAl0szFMZBRWJvbtnKQuKW1VKvh/g2
GLM6yRTYDcnnkzmD5JYVk//C36JGEQH1Q20teLe4+FRlLLo8kNnSPVlaGm7V4gSCjpuTrXV1DRup
aGU4pmsozhnO71DMcFEe3TDONKa59jEJEeoTZ0Znt15yP5R34VnDwMIk++fPYQ1W+QWt1Su2D9iu
6+nfXHgyx1gkfwbv2hGiKT9qyiC+dcuUuHhZXSXrLAj8Dk3UymTzoPINYECYLKZTgLAonuwgMdZs
ZctCXGF7j0qzMPbJaREEGBsBDROfQyY8B3mvb+CY9ubJo8+LBkze/b3gTAu0pVG/PcPEBkT/oYZR
7Q99vDv//3Ke+dhnyXzQ59ShPGFP/fEvaAuIC9CpcR3Uk4eS6qdIfeDE9wAx62hFoAerdFQnnoPB
WPWVS1qFUBej4z0u+n8g4ivUITVGmGD5frw6m2yeZ/EWYhhleIlh1mUxdkPW6bSmvQ3vkJnqSsZK
rFYjcwX8jNK8P5CgaTRMU2IQH5Qin/G2HvGzDLOMZYL9rfhv11P0jrA33bSUPncloXlmvv3ib7uX
symCrFPbWoY6bDzhz2Z+ge6Mz8PFI/cHV1HRIBsP8LVk6lPVxQQ/oQQBfhOlk0gEoajRFPCB7ijq
CrPdjir/YVYPD6ZRrqIxltEyj1m8B4DvsMQfOYimVSa7AxlWvA6HnmHsGCyaEEKYu17PnY4qsZjU
1yasHjLaU8n3EJCSa5Kv8J1Ajke1rzQ8xv4Zsv5SLqPmI7tkc/rp41/UkD3W9p/RYUBSPh2Erd+x
3J7fJDGOdxR8HuMP81pz5gu6adxzk9MD7EhvVMy231FpMHrEC9rIRWGHu/IkkeeQ1ms/tKmV1lar
fZ+61qt8uXLH32vYv/FXAhYh5FAcL8SCxdUqEK0R4+nyHt1lXeYIGik+CVSVFceFnGKXtYdXnhEv
ARkoXJ5iqUuZR+eFqHmj5FcBY5OYeqXQr4QhsHSuxh5JIeH2/R2/A/+g8LD7NN+psFqJYVyRQd5K
H8cb3c+zd4Dy1q6+jlURxbJ9EMIPEyBVvYFjOWVG9kyWP/qIe0dCpL8wQAaz9WlBsEOGybk6Msgs
ZeymimuhS1LBilRaaxvKrL7R7N1Dq9fkPGErFBnSRd4EwKaCvSHT1AVs3vgiKQtIRBO7r1rwoR7c
2XBDzIGLsaPKs/HcXB/mk+uhUBfeAW1fJ91l7pc/aK+2ZH8XzuzvAwoGi10p36LdZwO0RhnX5D8z
swWs0tnJU9hu6Ye1KQVx2k27+n822b/AL18mN8hlv1sx+6R15pqVOFOZrLvhHP3JrkD2Tb+IMtZr
6+tp4LcZnUuDIZjsa3AvPxFmDlJgpSecur5auqf3uR51OHMINcoPPjgoOhzfEJJL9eC1oCufMqQz
YtJxxG6PEUJLmRPpUxZpS97Mv8Pi8+FI8nd5hSIxy8JfLfhGPk1c1C4BmFNwMSVK1buv5cSwWoDo
VZ4qWDLYQuZBvTYp0JEnuGIfsUEoD3yn8Xb6Trhyxow3EjYi7TDKUC0f7N5H5kQzdcuXpDbAZJaC
HII98SXbjLkH7IvMOh9Xn9yXGByHKvCgrk1TWU9sy5Zi8nEs1C/9oGsRJlBBuL+vXvFt8Zn/e4zk
Q8J4kp3bL+Li6OGGZLRpGRcTR6pOcAd70pKW7yK7qhpqPJnp2mh3vJtDDb9kjLd1YCxm0gpmvmWt
W3elzfOXqqpdcn7v1xdcfGjWJb3kSnMUbaDd935RsfWvh1cBYmG32jSTZaLQT0erV4iGfc2nEieM
g2Txw8E8IVqspCDzkPbmySndbo7X0U/hQu1G2olAYn7WscJRxv54Fd40qvVmbNkqcUC+fUPQInLx
w0NXB7otN5I3+Z6vPYJKKigUnaO9W7yaheRVsHXwKwauuNsto2FHNaBfUE3MHFZCEzct8VcwA0aP
ubejXIs5AHqdnRBBRMSWM/1ZKLxxczAhddQaujFU/A6MAwHeJLa64rV4eDSzftt2UOYoRg1TICeB
gOw7feTHoLEXEU3qyndvHzP3jIwowvQ/WFlpoBH7GpD0yjlfhX8N+lnHbtek/BHd6TWRC2/941Lv
uNKMpB/I34nJuCOEkKquCjDcAch6vhet6U0sF3BvUl921wxcjXyUBY9gYX3NW935bhINKizc9ib+
j0Nkn6VQUwMeM94GwmFyqNTNxhEiQhyPQjmnXZdHH35J65Riq/4n+wjrfRykZNbip1v3L4bFk4pk
7sRO5saLLQv1S1KjUoCj2tODNDgKv7v9U6I3c799s5ZIXJYZgBD9qE2uJ+2JrW3H9+dUU4IKRbJt
mKQUmNtgpYLdt1rxDTUoagHJF2N/JV02QtbTOG/RWSH0MJZbJRi5SCi6KEhlO8hE3seQ0b7c/MjW
avvYnh7MJIgqRx4mQZ1ddwC7coN4MiLno+8mrCXk8YjkHrSJnR5m0vNb8HI0TiNpZPJzBBKOegWH
78rs4XIrT6WhZn3yWdnRAa5lUMI69eSJKsDLeBWE54JoZJqsxSyQPeq1/txNiY75cjpQk2ACQPOn
f+hgl0Mm5Mm+At+KrNhntVslrgshFEujMIBEeAkGpLAMxDZ0zJ4HyxegsoO7RX025vDIIEcB6Ygb
UeOLTBrgeO4twP/trELIzCdqut1H2o+PgqGDFCw7xuVlstDac/H78Y3OOoqMM+zHFvWZ/JRGlo22
ue0HOKmGBcaUy+XuPzu0m9iTjT4yTuYfXeo3V12VmcoILlU+DW12broZz+XP41zD+mtEEivuIWKW
TDlrQGAmlMI2wnyY3EswfhT/VhwwCN6f13vDA3Y7Khxic5bKMteavFDf+EzT8v3/NcpDPpb4NDtl
0m3o9BT2kI3uZqhLPiVcD+fs7vJyaK4TIq7kVH7DQuExYEBEXgfzkqa4t6U41spZ78FqtZAfZ8OU
QrIcMb4a0z1Nijbl1JowHz1fWDANdQR1LEdLfXgpKd5pqDIYoRLhhXOYCX8/VVOzxeD/vPNVI1Yo
o/JYgtwqd3Ti2+sx4S0FObOIPzs6pkJHBqf6c7XTojd04DIrFLc/WgoJOKT0T3oO/jsf1LKFRpK+
IB3goS9hw7Qyn0bFPDTqwPlcekDGi1LaHdTPuNmwwRISDdwnlnTjga9T/dxY7teVgmlc+otMXRfm
GC2hNK8n8Ij34xuwmSQRnj2mdHQItBXx43s6CHJL3eS7vdYRYzMHfpjI272IgJ8fTFL86+xnUCQO
NZC6IUUrAuDJbUjVaZ1jX2Z74hWhrJ6d31aFnJM+q+jLCX5kNPVxUaNqsSSq7YlkusKn5eGlFIGZ
i8BllD/3ECcKCWZA4NyuFCP/EcAn2DUu1P+VdQNGQ5WHAMJRQ8f9HFN5Z8GDDwPCdpKZ4pOEqFY9
9vYCMN7MmtFIObh2mG119b84OcArVPLVBD6086kqzlMQsPscKT9AkPyRZiHoAGeOxxlnoCRp/oEz
6Dv8IaqG1JiHit2doz0BMxGWURnt4vWzY4I+8PSisb1rOn5WIirT+Xct5aAcApZ416yEzDcgxSL2
DEIwbbCOzW7ivAzxhPVBgPaxLVEE4xV68h3LGxtbaK9KPpcfKYBzEIREgDWnrsDE1iWV2bC6dqFU
nhrPSl7JgPo1OvplkosHgQD1Qvw1Cl/24V2XmNOEk62wrBbqbe+UKgflmlOZEU1POW3y2oi6NGou
kuBQCv3M9WQz3gPeStejqMWPZyIFyeqm9il9unz33dty8eXlQkIPT5KvLtu4lqaPm5Fpa9GeVcpx
xLEmvqJ6NTQLhW/NAa9Y27FyqYa5spaVn9xHjRKpmI2o5WHCDHgfGIurPv1XzixsIwqKYopfwg+N
iAyI/D32LfavEhy4OPTYuPajtPdhoWWhkw8u52lGz+OUnC3yHhvo6wqmWrOaI/2CWFaa3XIajpii
Kon5K2T9eXBTvzI2eW4dZWN5MLwtX+bl1nhN88CMuVUxGc3rumYZZB1J0adeDFKPS8Wj1VHHtWtd
EPff2mNAMHyOlqKS9vD6RcDiUTJP176z03sv6ldvEOaNfpoFfKttmXeI4jKs7wMqXH7IKskoQnva
o6ANqU9oHyavC3sMqzcAIRkyArNX95sX8qwYlJLIvusJ1recWQ2pTyeFFKsP8mpIjLEeDGBIKLDy
iqbD1zDsk+YklsnZiwEQ8+IH/J27Tk42EJ+n0ptgPzjlz3Ld/YhliPc602/IhYwDPc+Gk8/y7hKf
/2xtXLAheeapJ30TX3ssSvdcnn7j7bhOuQcsZVxMDd6XAuqf9Sm9hI09uCtMEwjYE3cIwYsP3JgC
dDfOnuf9EiylKB8uXST71lvsuJKpX0vMsuPplOjkxpPUVHbfhTKlckHMmyNGq8d3p7VWg11UYseY
uV4t8ZjbwCgtPYS+rZAzhBpfSdFi2LtZAdJ9CNiK6Sq7kQxfSLlT9SljLBkQjZOqyvBBW2PUpiSi
6vAsGA7T5nKKorKzpnJ19CsN/z6sPzEjF7t88K3gdqtuCW3MjrPPcMcF2yBVBCTect7R0yf6NTVA
vWKztNn0I1SVxp3Io2L2oAi20ckGQjxZmLHtPLF6JL99gbIZ+wirq/nzp1vftYH9WIZz9AJS2p4C
KuZcFqJoW4jezNQCs2Heyfp2GsW2A8HmoyUiHsoNICoxwC+9RCR8rH7fB/eCKVn4qRFxMd4GTMOB
zUVPFh+2cj8zEvdSRnNn/fT3K/6Zi3e6HCFY1O9AiVV/uvQxai3dc/Jd9SacxiDFQUWlm2pbWHER
GfewJbbZHHha0l2/VpQy+CjOBNdK3aCI/LugmNxn/dQl57aT/nto3R4CuxutogvHWUfCH0BqzU4O
nbOILDUMylGizYtWEaekNu105Z2xRs51zSs3MlkZxiH6LiOXn9atPr10AmMMmITMUwZzhL9IPU8L
rUwkdyTL22FDjF/dm2KFgjAHsiTmzJIpxFXuDMO89KzwScdXdO1qDrquD98GjCzFqO5CfUHudN5Q
6gu8ebZmdMvJ+u6IYavi7RdvmyMBuXj4AFg2HBDhwfBNWn2RmvOoqrm4iB/TKukCfY92phMBFE9Z
VQyFD/W0f+KvdK0HrbFXIpA/u6FL44yj6Ces5IzbC3/kQlAS27KNd6rBNSAs8zSbzsuzTF7nppPk
pVik7j+NY1a2MfW686BbvQV8fsfxjAq71oeWJBTAR1CrajzGgkPrFdUM9jrG4be+TbJ0j008PGCt
OXY1cbFU/KkIUgQ5YyQ/BXWktpeLQ7tmML7+sFbXQQ/YuPpAYcMF28RLd9eJhC4V0pweRqCuGaQ8
35EEk9ZkjBJ/445hgPnGUEZhDanjwrbnDBzdXAXvjrb9Q4EHCHx/hMWVLXtjIFwd9UDrBI3btr3f
S/EMnwoCe2+wVHKzSU80y9s06aLuMUXVqPVIId+iDqACWgEGC90+8hxdG5WrIbnmYMh/+bM3nkSg
ohdaE14lXgr9yHdVrdo1AgGZq+bVsXs8sFoT0UxyNHqsYippZYki0O8xOmwTpzBcVOiAP1cOGEJW
VSQudcXN/1dsHGrER1n+THh7r8S3be4MEL4FQwXYW34KYNjJru+I8orDqnHspFe/GeinWXE9N1lG
9WWa7efDwdIMITzuamHT8HhYMAkiKccUdPgcXQXjU5D7nF92mLd3cLD3E4Agun1/RQpLRZwUCJnY
C4OlvvcK59LglTLg1NvJHrUBTJMcsGZGge0z1AtDtcDMiqRerkpsByn/Vhf4BjY0r/F1a2utdowz
kwhFAz9OmUPoU1PAAdj20dGFpPtTmyIiMTRi8Rj4e24dTmyApgCXBwkx1JszqkWVmLwx2fTPvZ4v
p4t7zja2UxtMtUB4C18CWYCRD7ZbXsvIqydqTkxpvQ1GcY3DN6djAjuWL5go1yWYVpy+Vif/4s36
HTju6OE5DmyfprxNTEVCl0ST1H1l6F0PxAwsCijTZSwKczTyz9zsAHfINhCXJzW8uejBZkQRG1iu
DlD6EHjDs/58XPAwjPbG1QxwyNLOMokvD8NbjKRGeQpejiYRw5yxK0fH9JHJj9qP2CTVlBYbRNhq
zv+tDwRDIdE7RCPVteUyUT18DhKLPiQuyr3wbVFzn3d+cr6VQunqRxvrxv9xgunMFxRwZSilxFso
JmL9gpQt7pbqXaUmvmRI4jS0aeypERkKt8kIYTivDkfoPmJW+diELq2qEZloGq4xU+t08hDbeSqr
0W4hRdWB8fbUakjEvqzwcLH/otO4rVlw3gMqIByRBS2BGWJnUdylHDOw84h+vtGJt+QGpaI83B3n
RvQ3dAH0+u99Zv+3Sn20nInkzgIfYZYn163yKUKiNMVKbB3kAOSi7fWZ8mIqDcYsgRwRN7xhhtgn
hWVsDrOf8UM67AR7vJuhYWfUDwHXgjOlBgx88lGbf9vglBH0PG30mmNgjPYOwLXQxPToHOaS5a3r
UxjOuwP984AK0kd18BR+vyRApiFG1e1hmNXLjBgX3mQspomMzO/rzpVHtfp1HZJdu3xOKTLSatdq
4ePvfHU/2pVePhdmK+Y7RVpPJroW73ROIWxdKKX21+gMnugIZQHFWqF9b+n5ts1vkztI1lX4Xgk7
GjQ5c5Wdj6JOOZX4FMPdrVxDS2ZSgok3MPCiuAku2SLCKoDqcxOMY/xWCJIeXQ6rCqlTdEOGU6e8
Hg9x82AEiq5oez/uCsbhSU3p9OarRqFttHlrm3A8KfAlBAvBsYfP5RdbIFmrL2/cO0DZz5NMV7LH
zGdnGYhtmtLvw0P7P+jdzSpuyga1/rK1eYmEqteOBQv2rtglkADhBK/INmpTo41aismGMkS2A80A
TtRnn2zzawzsm++yYcVCVHv2M81YRFuFoTXBEKGLWZln5L1cX7UkoF7XesHkSVchOSg8ExlSFz3V
EjLfuhSAALapA+ZG3vAwAZbMoAxBgsBbVSKTDjM3+5q9MWHqL4PGYahxOuEgw6orFbeV65lNEhOb
1vFOXEqjoZkyyWSs6eocWyZrWmNJQRUXwwBGT4zxPQBqYeEa6lY2k93tNMnWdrJr3VP6+xd9Lph7
AnqpjJ03fcnAB9Yw2Xj45kXM90aBBhIsjki5JtVvnwWI8WAndRHO/OB1xcqWUip4RhKPlP0gan+J
ZvpUOUBpGrEpfQJVQCFpTDniwU+3CVhuRQIFdw/M9NxDTBEv+P1NxHEWBE49PLqMzKo8Jx0ambFR
atYlg/Twh676A400Im9B8UUqCzSVD7R/TS+BCE8DlCIWBwvxUblfVQJuP2WBjAICaUGS1cQYf7O7
7rvS6ymbN5H63OE78qZsJ/ly3cbi6rl9O28uz47RejXDOBQd5Zj6V/t5o+/ZHfo7VNn9Qq1axym1
7awgFl9kCJiqcCzEgkQ/Uz0VcA+58QnwSZxpmWr3aByeMX6fh0aC3RW2M4VWn7ZOK05eQyPZNMul
8BRRmAyLJu2Z02oO5dRgkxCGe/V8riHJCa9bzmHJEDV8iA+GXNyK8siX5yf+3sNvF21Ie1iaHnnC
/3fPy7uD5SImahkJgEgwGuVXMvGxqjjNCJn9lejYW6jIGQ3S5Tdo6ZIe9728/J+mw8vl8bzjL7cM
KlVpLZaUgYIxCmGwV1ikcnMeyyr3ENukzL9RfU3O57vZEouXOKm7DAkZHhVoAIHXap9fNRpBS8pc
LVcyvqomKAKUCQ9spXpXrJ1TDwx0hKvAYM0S+xPDLkFUD2VIiv7Xq3N8QqwNm00PB6QimShmqwgZ
AcVYiZjEL7sRIt5gm1OQJwXKdcbNQ0gRkUpan1MgYfX1qvGpSgjd5U0OkBOJKUl4QiQB1a1LOuki
+/Swey2jtA5ZqGDEOJwhkjr4CEnsm0ppIZJzPoF+R/wlmGoA1ivvcMoZt4DuGzrycr0nms66nXCR
dY1dfPad3O9VDDG1BLz8OeSLGB+3z0UplJCzMGGpMfTY3bgoBO86UHisVOFggFe7rwVXkcHCoK17
gTEpT067g0clEqeNVWVu9kUPQd4O+AYwKwqCQdaIW0jpBZwPbwV6cNHxzhVhEikFaAwk5M3gtMSD
023hKjgeyIhYC8Q4jS55Ykw6DHRjrwhlPawmrlSP6DqYGdpT+EsytOpUQt7G2nLlg6vYXmH4Y9HX
ffQuNF7u4qu7hvB5W4sdBGthYzUoMZVnOCzPoNCepDHgmy6iQf3dvf0UPQRwRXnFYhHRM+t0kZDW
ijsyc6Rx5WeQCKu738bz2Idlk4v4/QJAuB6oJg97/DcY+8rmUQQTZRXWJ1O8pU3+3fnTEYuHxRju
YqR5ckC2ac47Hfl/aUo5zXVYmKj68eYgAnIAByEk8d80NGkDMGYAXsPpPoQwTcC0tRw2kR+COiI5
E+owkrfXjuQLJjjcJTasCk6JYpY9MKc6ebjUUCNJUK4sc94VrG5x/bmKRXN+fIkAgLevltfFrgTS
SFhHWMlulzxbIPZfOinOx9PXh+I1cJYqQ2TbkNq/Ww44OxsZw0GGllodC34WFDnhej5c+6S95Cj9
3RTCQ967L7HquN/m0dAQ60FwOFykLwfqvjtozvc5jIvV8Qy9V5xrm0xYoeD93C6iqAu2F+n5hqiC
DrndxDduZmN3WJTlCj18628VML/yOPLRIzwJiAPAsyYcS5fm34zg1Z1QvyP9NSmdub5gUNCEb15z
J0z49oLTaGgi926QT4JpvtmNru1OlRHPqIQDTwaFOl3QYmwkWLU//+wnaMkyGoy3sjucN1WTD7MO
lGWtfSpNnyX3Gg9CDf+CnqtxKo9GTz9yvtJprQeqKi1fa0l0uhFa3yhpYlwgn/5QVw1T/yHS/EDI
g3eEuLzYFqO2+4D/Wgg0LArUmX+qs8tzAnYqWhXMk0gIWB3IkO5qQsntvd4zI0KGEaCPN/J5acHr
zcx5Mvl1RJWUG5f35DBv+5qdu0JEq1QAGnGjfMAioIbDd7XJ/Ksz3DvqxIuoDG+GzUc73skM5UJq
VlwAlk/OCIsGOWYS8hXrdFGWlIGaDWKc/hZQC591tq3C5aLvaR0w7Tek/2lbZHhTQrKdwqrA0liD
4ytyMvXMzS4WhkwocF4B187tyIg0dAEBUBYMm9dEul41rf2oTtStRaDNTogAIZ6iM9MMQtMpYyhz
PaqkHAB7uYr6fcMeXgNbdzV+4Yt+WPK6FhSBOpKfUWDajhuJk64+7ywrwLK72ldIsxrsg0fM5EK3
4fCQNwNejgBxG4HWkVjAxYqWlKarJcPKSi3C8N9B4I65+NNEziR5DV3u8An3drBrRRrLT3QDreG5
0SM6szBJqp0uvvP8QMgCwArBPIU5n0ApkZEqhD+PXggsHfjfj1JgW7MRGm2bc1LV4UpxALUE6Peq
pudhORgilScaIVpJkk5ySWSg49riZe2iFSfv5ODtmEBrH4nq89bnMPuTHMO0+yXCBWDHWp35l8bd
FOPCgazDjfIxrPhrLgkmrsXRsWHtXowdyQNLYejoOUEBSjWf4i3rCYpM/dmUPnK22YgFLzj9Qtld
eUlJk5APiFUKHYRFUS7XGRGvR1+RDhxNRCLI8rZugXxGQTe2xwWYxni5Xv7Bc3pvtBI5KpuazpZc
+/U0r+ikmtyes91bGUExcnA40aq1493vdZdMlcajyH+k/YV3t89SHmbsOQ1SLZSiiAYz9IBg1GJn
vgkDTRQtzkoyYqWsBpO8dlGDsgT6WLRVgg5TQgbsQvIM5U5ixADHuE1o3F9yZa3Th6owpyank303
SDiiZ4jU54yG1zB/8n3a43FPKg0a6RvwveJS5FY5IwFzilfZUKudyri0KcQnA6YBdnwTElb2PD3c
D3FcQAjzgFsABgUEz8l/ngIeUbvw+dtkyk/jHgargN7YLhFHx4Cdx5bLfC0uVKw2FyTd2+Y9775Z
B+xBHZMfkZWch0oWfN6U10lLmiMWDH0N58/MtFpysiDUvdMuUwRbJj0QRoZk6boQR7AYxXcC5HpH
mBI2Tg1AE/pF/UXXUE3JOOH/bzzNwzH/2L02TJGdXL5Lu47HRRJoHcxEe2qQkuP2jop1KgKMJjkR
zkAQMQt2PFB2jig5zUDT4s6/c24Aih6pfBayu9NF/Q4OIV4U0EsWACSzk7yZfX++V/X3EPhVIK6q
q2i7skSe5TYDJgeTidGcD6bibQhZ3V1vIepxnnoMV0KUbkss9gDJFddmsfzHJmCb9UhTLdEP8UVN
ZBVYzMSHRuXmzq3vQnN8yiuLmJg9oVHWBMpKGvJdN8uzlcoHga6gIKqBuT1z9mWw2oE1PneZx3Ne
W6YtSbIhY2jdusQjJgjOQmViuq1GGwd/F+/xSScfPhOWzYkIfEMehVC9GxFzjifwfxDnFL6opVux
uOaBKw8mpgG7di+60sDA4sDZiaocBziYVel5Zw7xAMLGDzhOp0c1Ftw95xhHFCDjOgCF8mHHnfxO
fGER/xTk98azqUwBFdkPw4xJjXK1Ps+/XEfu0KAlJZO9SSBeg6SA1jtVbzs+jNFBSsncXdUm1Y25
ukqG142MWzW1rwEZEL201Dy8Y9qBNtNi1WrS/v6DihdE+rhPEJmncm62L6zQYLHZRuAqhJxcAuWM
7bvu7crmj8XpnV2qH9GoX+VqKvgZfNHIx4ntUg4hdRHZlzLKD/NBsLiQfxrFJowWGc48wJ/cLM9C
kqnwUDYd1MnAzI0QHHvAbYdZ7yxYjkUQcFRLYbhPmSXrlnq2J7kOKrhTte6LVPJoljuTaQZIhssP
GxhMbzuBSY3xrD8wKm5axptrM1AfT2tTMUvJp1NOgGAPNlHvDLS5xU7Lz5vlKB6E0AwWacps5tzD
WvXUFNWJFkPgzwYsBWDJcC3+Q0ocr2YNbHahczI0WWZ8M7stiqx50j3S0BXjO6K0TIEgNd/LBy+t
KkooqB7yINt5ZHKuUZTx6BKQ0QVaCEA7rdrOnsdqc4z6sZ4/ozNbslHOwJcgFD1HqVob3j86Lwre
iJ4gMCUvKIvJT00gE9Co7qbtq0yECQ8k/rKWRR+k+z36HLmemwYpQwch4B4vZjAiFSlgTY2ubGz5
ucVMAMSaY6wOHMe9JSv2jtxavKnHP8eFGB0n3buqCxQysNxqM0H/IRGok5Cx0Tpb400PpxVixJNj
1Qg2V4veAuTwr7IOK0wpA5a8u4Jyy+KRh03aPTYGAKBOrku1wfgA/cAi/Q05b/yV+8jW+hU2lYx5
svp1TMCEiuuTnCeN4lbJGdnk/tIXzSKZ6fzcp9x0HvIMlPaMu06VtOo72PfNiVSdGHMxB6bnn6Vg
mbxM34R7v1+PsvCDmaSgJ0L9mVWMME7+p8s1AO6/TT7+5JOJ8AXK6ctILeIl+Zi6JMuaZCAeSqVl
Hb8yru5MCvRSsmghdCQKKRQK1VHPFpkyGWZWfLn+i0b+Hyf3Zp604TM56tyIxqCKqjpY3aLBVzvx
7ZYvGji79rupMObwcMFChUQ5J98H4zWwZm+xTNCiNeZnncO5mcvPmrETSj+x8N7DHGxBfCDODUk/
oEr8OqiZGBHpbp2ZrOAVCQU+qKfJqCkSPv65QtJrGtqRabCKhz7nEl4drCyFLteiNw1/6csiiwrC
UeqIdJXXhc5YxzAqzT+TJw9O7Axih1yEGgC9WZmwAp1//gONkfs9Iww+GIAgXadf7XUVTkZZWA5N
g9aEvS7i3Ed1RWZCrFonLqMvbf0/DvgLCqaQbMj3m7eZ/l9UwGbTF3F1Nr1K3kwADkkFWzB4b8f1
tn7xqGVB/g17uRGsJ7ZtixevT7WoaFn/Mppv+DN0qGIEWmTENILYyVH8/rqWPCrLd5GT1rw4Gqza
wfzfWmPVX2903f9zItZXj0gqdBBRpDtvJSNhfjoVxF/qsyYX29YXbDKKrdzhvD9SUU6PACF+lLp4
xq/cXvuP2gzcU4diRmNxFfXCMMOcakJFFs5cP95pX9mYC1X39Syrdv/SKK4h1DvL2PshCg8SopZ+
/NIsG3cVgSQhXkWwkmdBFV9LU8QiQttbQxf8UA0SO0tttLMoabJNmyhDJR/Wfh08FVdLyvegkZ3C
Jy25CxMfgilqhZcX6lISr2CXYEhuGgWe9IUoQ7u/9K6VHAYcmWW8En494fuoWgk0l+2zTrLU2eha
D8uebdEa4u6MbGmRcQ8FhSYJDRKhg8gc55fbuoOPKO3TmF1W+OC3ZxyOTI8UOdzRE3AJgQt8RLRe
V7wewk7+xfAnlwixmy9LP+NOZfpzLR8W9+JPpNk+jC1dZdrz7xUs6oJfusozC1hRQVaqRrDHsfuD
oy5baaO/lyD51dEEmoGvlXCXEKqQQFFjYTxtg19D/KBrhdQ8r4bFkbRwL28OQBGtuKxhOiA1Swic
zR6fRlLepKpXNXVzrIjtOwI8LgJsbopKbS4Eh5Ohvg0pVSsxsiSMsnNslVMh5a3XOhAmNQUydfxQ
EZT0+6wt6FWxgcL84XOQtFJXldd4ZVA9gKHnvxiLh5QjMCyuuiewscAI+SCzkRMWlA5YMNy9AU4T
p9sQMlf0jvPYnOxzUZ1gdsePK/eHjV9YD/470VXj1j4fpie/Q8vZme6veIDbCZDgaTDGquu8Slov
TS+dkR5Ah3EjlC0CT+qUEGrQBq2PlU/Spzynxb7nSIqzug1ZwDV5AtqgtdQvAuSaY5rbAkFSWqdA
u8wJhIpfWe7KZDy98U4wXDWL9hdq6JJ4vYDv+B7fCZY3LMCZntfqquj6NL2fMND6HORjnNGUyfLP
wHJe4Ud1ZROY08j1oM34J4co8B+WxigWgXvOvBpGdqXhnzqx3adVC6Oy9N5aIbKiEkeQZ6UjPB8v
wM295IZ8vxks4le4TppCbG1jCQmgNgdQK38cv/4tCIVczOgcDPgrjYIqJW2wgGavKhhPFInk0eEq
LBvNr6KPWkRoxqhAvAqQW+rcrxdcpVxRMzRqWjwZyiFoAsGBl9gH8Qo1zIzkYAs3THn/3z/Aalf4
b8EDgTAxfj5KTGs6iZhy2iU39hyEgS/pnT1jPqM8O9wx7MPgbZOXBsqEyLfoCx3c1i5qE2d8sY+T
leOkVn3qTCnGZlho10xEyN6NqNfta3ktMlf3alwSJlr+om9lqg8aBuzfjRqa6UbKEPwAZ4gkYcQt
8HPfIqEz85qkRRVI9mfSENAUZuhJZydAoqL5b9nmNDwa4CaXgcqjFjI1yPNIPP21MFAjcCE0ePHC
T9eqbsnuhXMNfh9iC+fQrD5iqZwmFuuqK4qP/Z/V4rKHHqHfQ3fPJSD2wZocBb/azfB/BoBBPuWm
jvSCDszk0M2ECAs2Krob5YI+U6aBKrVSwEKGj7aRJej5O2N2Akv1evO20cMcMDYGacbsERCmZ+fB
2GChPQcdtw3Ev/ox4XHwWXtV+OPpoqKcX4GML2XimzPsxB+1oBbnZHzTIaZ57GPqVfGKQy9zktT8
u5wtutlL3DpT8cz7fqH/Pd+ZbCqKTR3OFNWoG75c7XGHf/znNWzaLGuR3pMiKBxGf0RYqpSQiJkQ
xqb5BnXeiLcukn8KnNi2FOa5ZOK7nP5JkYXQruwlVeiVEjuZHMfQ/9q0GEHii0wlDxjZYJAeOrjg
GDVCMyFFGVJeO/sQdPOTml82qzdncs9X5HdOGMSMt+d5GnM9zl18mxgUQ7+HtnmlAWMZ9gkb9WFn
1aKRlypHN9VDiFq1KTLQ3FxyGrVVEdEQ665jlaQc8TMzGeiZT5Ov+ZokxShP2h4bPhxcQ0a3/uhe
nRd4rwDToK3pA9wS5/QUFu0JWVYqXW/MnWFdk+hSLB5FN4mEECPyhKwS7EhNe8bI0d2gzcxsZhqm
nIPj6BaqMCoaVt24xfoAGxlg57qfi3QNa3/ewhnArQmo4ZVPguKJ1kmRW7czCtuSvhPyL6fdwXg+
UnlfNNa9+wVaHh+QoeNY5KOgQvwE9GSAjbn4ygljFxXrYmL5IOmNcjEIKD7yk/dUfFKFUJZ0YeZr
78u3mqZn4aYZUTqHKHjvvzoYoAVL/WHQNyKyBNky8tjXQf4Zb5mFnLuPin3WXYV1vLWw0b8OPs7f
sT/2oczz1+kAabQojqjPm6AC35v40oKuB1t1oOw5gk3hMn5ce/7mcESN0IWZdts0RDilJnUx+SF6
pRMdD31E5aTnzP9liYAbFNzxJQWcqgIZoddA7x+QuA4Xfd3KZbwYFnCVqIZCa0hMShq9jT8K5HM5
FCaLuYjypa7CRzgm/Us8ExIoxxkn9hPsyEpeT4H+Gs6N77R2Ai0OW5u8VjC3orGwZAFx5wEJLycE
EKNiNmWNOJdadK5SgySkSj8xwHlVtAhkxojuNONoAVtyY9cXYSyHN2a9G/2oPcNjkUPT0pb41sxb
1stRtKnWPS2eqeYBlUZWC2AgOOzy45FHPTJNhLOqoOueakePDGAY1b2wdnCUTx2zulFgvJ5j1z8W
l4lh2DChj2w1sIVYw8JQ2NAax4+HgbA6g75BSIc648u4U/jBhHemmWIdJcefdqWuu0Kw8xj49152
f7KCV3sDVZjyu8ohWRZAzuUR4hGuYAwnBzoYXvJUSGHN7hvBmMYF2i1lT9lGSKa5RRgw9A/Km+sO
zF5qKUusQs3PitUz8Da178elXrkrKGpb+nYPu9abqIqy3E3U9ba014P3umErVzJnBPhKuImZJFlT
48RkCSba6jUekpTEce/2cHqOKWuyvZaE3zYMw9a2SLKu7gkMjasWnrpbZeQSwa/pDQIytDaS98Nz
u184lpj8giXkgOabGwefH2Mua8whNQ2ATOj/xDxQ3hTS1WQ52bE/ZunWwjDrRaPTKnBnrBw8a6B9
Ftd1FuEGOmAIeCkAp6QklfAYhDtSrXB2vxST/HSkmgOI6y7y+LtEAixaEpSPjYf15pQ7ymrCcmW9
OL+yMdUlLXnbN4YhSgbJpyot9DObUDqUHY/XmBFQTtPHJTJtiWzLSJW4YHLrAz3qQIwW74/kKC20
rlhYllLqaj8Twr9hiMgGUxwJJxIm6nhH6dOxTPPL2vOsUPlxQS3FF5kJ65/M1TXKrPl/8hDLHc+T
evtPkQUPhHiV+hnOZPbtcCt1ikA3sDpuccJePj54YpbcPF3KRqTzggoYNAjNyjL3hU/ic8BnEXfs
E4XlG3xAWAAUTNhstDti/Q4PubEKRSx80VA4D78+/pDR9vivBlnHouG+hxpsTZwqaClfy3Q4Q2uF
r20bZu+PUIr2OMWzYbiAna9aO7/DQcrdpD1fGvlZXbINd8O9lMnKi1sQzf3+ztROAl0VKvSKMPvH
r1FZSwQ5mauGIgZn/h+GFKvHWe3INXvP86bPmJQcRueId5H1MFfKHnD9weFh9yiFpnAACqzI/5Ly
YMnF0DdhD+8//uGOyoKdT8IMQ3WWYNmfrhuN3T4QS61avPY3Vpn+Wgq1gTGqYbdsvfQ2Js1zx3nL
d5HioltELcUCQbyxc5wpSvinCWiycBN3xJARZnsWxuq4cU1GqMWmolXwl5a8tx7O4bldzIC2bjoD
REMWeFFlw3MeqvFWvQR97H7h0AZXae7c5dimj6wMSNhzvdlmeP5kpFMZHI/qTOx7uBF2U+mVHaVy
5hI96d7H85qcilmwnz4ZUCoMzZ0YtDJJDDDdoJFLIau7PQkAI101u3fyAxG710SCKbpaJ02u43E7
bJXnSigVWRyVQlHdatqs9PKSiLFXSs36NN77N4dtN7fvh/uOw0bPBJvA3Id1XZmrT/YOAP06IUhO
ao9cGFwDcDZAOSUgFM7SixkNSuZOvqJ2MD4Zn4Ub0kXjsO0wnKDEjmLBXue01dTmZZAi5pgQEv5L
ejeM+UQZnUL/fgjOlvpVHVYhKGrJzV4rQAInb/d2wvOZlquBrvr0TwzQUCeEhbF2uWLfEBmBjbl5
3/DPuQBp2s/S5e5P6aGXM104vHf3ccK6qXN43jiKDt6G6WLwS43uHWnU2xk5rwxmIZiatRbXnYwg
LS96o3f3yczuG8em9CeoTCoyJ/GcRd/WOy6BtKL3sd60DR22yWAY47SZDI3SIKJvZYdOeFcuHEB7
JujbcsATa5fty8jHAojrkFZFgCdiGvyfI+5rR0CDfMKvN+ALevdbNDqIbR18K9gDjY51YS3DWqlz
Pt/pMbD1ryQCbN51tUqtH2svnIQXG/gsXV115pOqvcFCJwkRkB5PQATsB+SL9gxls34RV4IUb8yD
qvlscEKnOWbi1tc94UpUFOR8zws4guCmFwRj1eYffAeXZTOHrP6wA6hxhlEI819MbYobLnQpAqaB
yQhOKw0Ayh+85VbHLczvu0ewon2ibNiNREYUzB6eLqAtxLt59YNYUlZWM/FKDKxJZs1/GNaJ9lle
qE0WAa6B7l+SZ+HbpQKryWrNyWww2X+DLObK78bHM1KjKnYL6JcEE6oq1B0cFq1V6YV9D5ZSqTDA
kchBaKzziRl3MBQgNNvecNS/DytoVLwD+HPAqPtWWygc7F7ru32PVT6pLbVrXqFytdRN8UwEZlfS
94EjTalkSdvD7TOSTK057yppJIlB0ZrwuwIDfimdZw+Oy6vaICByMsg0Pfjchy4LqkbPi+SUwaEq
lfANORHApr248N763PuhpdpduRQORxD6O81QAOuY01jWs8JyCXsBT4YU6vJ+bn2ykk/mkGmYcQ40
vHO4IOZClqXBVKnTuVnnqKh6fM6LLGrzo8rx8aFIvjlu18CdJ8V10q0YV0L4HFmKWPZ6wL4Cmd9k
PHggTQGMy1UgKfafGav0jEyKTYZWBPevtOv+0h3DzsmUJ4muvTjRt56qKuac9hQ/kiHzh00F9ZJC
M35w2UCmk4o8Ax3iob3Rcbn+teXBiheBAvYFyf7rsqz7jkhLXsfWuZkSP3LoY+EYkyZS8vNyQXFU
cFoKg8RzyYN7ci7zFTq6Wes0KQWK426hDfV6E7J5LRVnb0Ujlkm5dKgq1dfAc1YUYonoTXEpQK3p
/JlV9lbN23kM+UtxghRYoEqf//PXvcYyGPBXd8dpBBLIQjYBz7DBGGdjoyuQcYDlIl+pu8jxsMsA
BN9IMn0QLqE6KMiZCm2FGQNmg/eqC6ug/n4X68K3f46Ttgu552GyLKPec7kn4LCf6FpZqqnYhOxa
x0cees9bSSA2ZZw8Ew+oyf1Hn5qDOPdUkuZmmj1JKDwALyBvOY+QfAkqqMM1ce58QEe7uS7bJkku
1f0+cLyGZlV1Dvll60h1UTsk6V2wCR7bVt6498oXjcZeqoEoi3ytdx81z6uKDW/IKpq2kOYoA5ah
/aQclkQMFirF8rUaqVIwGvVNrPpjFBVVltLkRqxeuH5uirjA1T2RMwe+g62vwHWLpOO7sNsloKOQ
/RFggojNAn/eM1Fgx5Vrj8G22XPQrPfkt0KUsTsiBB7a7pHMAEifXI3nrCu1PonR6e2fBxtTnFRB
QaTGvnWsiYJR1UeIlQ/064/DC/2Kv/qwsZkfpwdWdE8n7xZIYnDKPgiNSGE6xBf6/3B/PscSJv+n
PXZFKv57fLclf9ogRyLeRH+tvpxmXkl8IBmoD6tZkA7hlYqGhANATDmYMVtwduquwFKClUQRiap/
31NbBQUZLbJABfKae45Qjf/fqQenrQMmujEBeoVpEghXtQ90JQrG8oM5YUdq5N6dtcYLJdBD7D8y
Ah9oYSG8djNIQ9QFD4Szk84Dh2q65GI6ik82p7K40IiSRhQz6UyjZMsr5uJsnd4EDQyFZlc7i2Eb
lrBt/6OLv4J6CI4UiiS+vrIeVfDTFOHIUngAmBGD7qm+1Sg742skBZFWC06aK67tOpaSjOrSuRm2
1T2A7iHpnTe6+ahNWcJu5NC/H5jIYq9czqMODA2euEKjWQsGIkH5hSwRUi/aiI8Dg2ynxOTKbirK
4ld2rfrcQRXQ1SB9xKckC6x7UAEoAhXktqRo1bzr9QUyyLMR4zsKsxBm9GnWB+2EcZDrJ1TV8SIV
7wes4Rg+m5WBZZnRzHIoQ6dXdU04uHsxaYMxeQfKLxENcb10iJ1k/prqYnOOA/v/S6Zffg+NkaG4
KIWSXYaAezRqPcjCGy2UluEfy5k14gDYQGHKY70kFPkWB+ZzErk7uCrWq/FZEfXTiwOT5sgiOY61
TE8t+zI0Ceq0aUu7h1JaS6uWktLySl/SS/4VPIEsde0q2K8f2SLMxfNaS/P0Xlx6jcZxzLcBLnyR
Xw/F1P8DmBwW9n1DmVaNVKChsMDmR/hX/2biU5Q5Y5qEeewEEy72DwJtvB1aGbEfT3oQJ7TU+6gQ
jLZJsRRba0pTiuIue2kHQoC5X8fdtLlhIym4D70FzXk3Wuh6sUCaCGe/4zC88AibdLeb2XctuyfI
E1BYfKQR9eG+/UdBFuRcksp7OIaGFYUFrSqcn5d88DSMw/fxDgP8f+v9on56Gn/8G6RJKW1f8hAp
RKSgWeQQlp30Fj3wXsOOj2bYAEvR8rRjmgw/6ylXpCnq2aLDt89l7hlQ0vAYgTUuD7KlJmv/HLSu
FhvjpcqrXd39zRt8291g+fPIxqinOPb8qTUShcWU4p5ict1owSW98KVKJ4SrKrkGHnSJ1+axCCzy
i1Mb+hp4KCVziixJ3aYcKif77pMbDWePvHhetVQ35p4ksSlm8Rt25/I6krh1PwVOI+JslOezN/x8
49imSsc9IqpQiAzPa3kWHvHBzRkPvs+W92aV6t8ovyiGl+lwY9/pL6rEkqHxB9pLTW3WPQ0gwYc0
Pr2S8UMRYJkbGNJyfk/It9GFj/GbjnE3K6TcHqFyNJ0zhyS0MbdEACPXrGqzCVv6VC++APcSsVPX
xz1neQhIyp1o30bTwRJfh7QPjFAJajLlm3QdDHLbKG22bT0YNpd5ug2jK2U17EM2+ybeUtllPM9e
TEwddXl5Meklx1ydCfs1xbbBMPo1PrEgHnsgV66JJN1IAQ2AddWeSWPyvCbkBiw6L2lgV3rugh0k
b5LepaeOtnV649oiFMLjNRBK+H++0F8Dt6sOmsQ6ZSoZCzfaeWtoEQrbZGq6d6dQtMEB0xNgBK2e
gl+6hhkweGOKCKiKeQvgtgG32LQhBdolFhv64EZ2bwKIunCbjIlN/8vxGTTiqCcgv2x8NFslk89f
GNRlotBGAE+Z9U1G7kzgaoyPjFvTgV+z7C0n7TOK5fvQwqXrs7oxPGSz++Z0lQPUfJ/YCc2/ZgUb
J5h/g12Kc3Yi4z7YiKt2+j6FocNLohyI6SeGnrc6UX3mOXHX1SpM2f09gjMamU6fleOyKL0ZHutQ
VMnYzCtn281AugA7ZRkhES0Na//n//XIQPlArfOcDTDmJg8Kfb1NLbydnW6vusatiJJgHFxbsSGY
CrUVdeAW5NRv+8d4tTDwUNvxe2o4OBLFv2z0w4qzw/E+5BIDicEQ1yFnjrMhy1vhyOG1F0vgvrX4
yaSn7fV6lt59VrTGIEl3ByNldv/3KdoSXJDNJtPMETyo7oOJOaNFOl2p0JD81v/rOy1LwvCHucVl
n+zMnIrP5IDOlHjNXz4s7IVvEIqW6c+kzNTZCFc9ZU/qwWLAu4e66rddKwtSmAqB4MSJ3x8Hyr0G
kOjxoBdztRCz2corj3bwwInTGmdJxrLsYj8qltoubdrng0o8lpNUUGKFCrWZkcfSokooW26yCddE
IPbf1I2IKX7WQI7aC3kbuenvKRgtbrckoteVVh/rks2AFKI5h7NaxFoy9mDrvNoqKXuU7F/VUk5N
8Coja1aGLST5KeYxootJyZMcrbDhohikzChqF0npz8qV3AmYLqGKR+AO5s6jd0eXZBnqp/alIptn
jvlmxELnenwoCwUSddLCZ3UwUlUT4Q2sSw7C3gLNUbPf2kZz4g9XqF4hWF7kn2DXB0VB9fRScT7Q
7mbub1v1K5f4TMTvb8XSLtu8YbQR6b2Q6sUfcU97/qyJci9Ttw/SI/sZ6IuEApIU1m7q5zNMgauV
+sSBYhZfrFohYDOIav6tmuodec68M6uc7kRUoAlnRMJPGa93rck+6GxeRS8LWv8DdJOiyCv54DKU
VApDFdb/1d3P7eJPoDvJ/SeGbyvlITm5fdjms0MBr8SL+GMiUXRfKpGeJZSoxiYoWMdZNMbniZUc
UlIy0mLzyC12GfX/o1rQRobrBt1Xw33vIegZJ7Pf2sriywqSkuDm71Os4avenC0MCwfmvJfwEG1S
DERW9QVoA2zBJaZ3rN0Y8Uf/+EXzb1c9wNO9/sXRWb8wyLBWrRVb2YcrUC8kgCEJ43snYOml37Dn
YgWKGc83MjNKjIZo053y7l8ynihJguFDYm4XYgksJOxwCZQDHa1qb8anvNiL7HRUXF6RzkqrE5vW
bSvFG8m3M5pXckwDsCOY/Tvlcq8B4ubF2FrUtd6bG/5MiAFbPqONfSryy0FTPpqnestmJTV3NEfo
xXOEBmANVMU6hEhGbXIzP/skEMjlpPBFb99JSmiTabsD3jwNFLKNd0LkwhFPZLjmh1uPCSK1kr8q
dl2c3ZQbiSWVx2tlcq3m2HwHENyRTx/veq/IUksG2sb3Yx9es0Xk4kATLJJkSF1eCP+rMs/Ryj7C
ZweUDofQcYvW849w6GYXIoKXbRUGNiu57gLSYwsOyD0T8cExqC9fa7m1MoPXmDVXjyg4pTrNpJA+
soMAzG922lvnVAyjjRMhZMaTqKL1F/MLzBx5WdThTniRJNHWo1eMyoolrsjA3MqTWEGODm95pjoA
3md2YKyBSH6NDUnFmzdU+yqgBIryxZp3oP2wnIt03kDgnjbkNWiUegKj2ar+Ep77lr4+qC5/osDL
TclPFFSTalRN+k0tcJkndiyy6jWwE5SZYMXMdSG0/ZojgVBhlpFO0WlRRqcDkSnDrbDxoYVTUk88
Flx0IJhC2sZHkUZjxIi89e+7zZvuymivwA8yFpyioEBjVPY6fJzQysaPWKOabwTDC137H5XsWu18
rt2R7itPp63ySK5IQjF5JRPQlfr5Jr5+Olfds/En7BcqhLRFIkvDm329K9bgTJmRfoQhHGv7StLi
O9VoolnbY+5NcrMpXxQozlhqDwAYAN6es/9Cr9eeUqT7gQQM1fVgdgeFjGKTjbh3RybOIHI5Qs/m
Yh4AxTYWftxSAVSjOMHirc0JvcJUaW8Hs+ku87Tb0uBs86s+me6KsmhH5tb8QIWHIc44lmZukEKO
TCYb1IhmsKxVGwSQ476yOApjHxVbjXmG2SC1a9XPxUhO392xqxeQdTFValLGm2N8gGMS5x2ge1/W
L3E1Tl18FHXyuUJsDrNXDKhGrMIJsUGXzvFmwxTvQATdVJdxS9Tp6ds5sozqPsGtxK6DExCtckXo
3t89Dg6HJvQqtKJ19W+atA+1W9Iemr14SE3oeaEsCu25q43vTDzUyA/ST4/Tzw6LQ/1d132mdFe8
F82npl+aoXIFUHv8BWMTEhm7PB9NFQLMKQ1C9K0TjtahfxyREDCT8WQO9Mws65Mvtd4WXNqGQVkt
PBFhXXOD7Tx2XV6BatMP/lsZSsh0wNO/Y0wLvHSijqGZX3G7J/toazNnUwOvdb/ny34IMRa0MFfC
4IcwDB0RaIDRcr067ZvoIDF+uBAzXdBFxd/q9fP9CukV8muAZ9uxlNrj4gwUeG6zlAf5ex7cDj0B
f4hrS00skfigurUbxJIgEzbtHnH/qVqCyuc8Aob9GmyS+E8qfgkO8H51HqIX4/jz3AFP4X+zn5fT
h2b9k6BX4BJyBBuftjP9OJkijJEz08hNHbZmNNDFboqcSpsvudjTN8QP0ytRL6jBMOwShiGxwrgz
YFE/8NMTo+Fo3Kt27oUUVzTp5F5A/fnj/SVecRQ4RRvmY4GU4KdleOwrj+XmF9ELutVogBz6KYmT
tayI3jOYoIAUJsDTPqc5311r11dmgKoANMlbZpdNK5KbJsbqS4HQg2NRH/UOTZvIVWZ1YUxduG4W
73aqB7Yx46+0pw9PyIt1oNkYX9KNTbUeg4ON3IeosBVlYZydzPLRuphqjXWhynTWquNnbYb/s1M8
aWYGN2VVIFc5PPFD+eQtYsRnJ2jsTZqC07UKoK8Oi9qNA83xtrQWknUd1V/FlE8naVRIaYe5s/il
7ZuWqcKVlu7+cdjrDGMj+dw8wLF0wWIcZV56KZg7JNFjjg9qQODlkfBDe5UsHBTNDj6Zu//CzD9n
zC6fGPkrnsR7U4976LvDESnbO3fDHa6NRRS+9FUtKAh0CnSPYcH5UpwFTZaCXxSTi/WPLMbETNuX
oVXCjsGpIxMMjUc+AARvR/kP5m0exANcOX3v4CeJYkB9Tib7kUgv3Gt65iDRpl2AdMeRYGoPuMcZ
q1U2jMFHAl0UTLYv/8yR1inVhmvlAIFyfxttokaoWg6J05s1fzbPGx57MCSU0M8fRLzTJ38g6zdR
OXIg6jRCY68Wco1vWrAX9KuEx9LfZbr37wtpr8jZIdlOD4DDemBg4VycsTM71ksKLYmGF8wla8qn
phR9dOyz6holmBxf8SJSvl66TMKh/m/Qn0ecjVtySjyoK5vB48J9kLSOHXqbF+i/L4AUUPsB9AiH
9F/IMZ2BiA+AVwPfe89suRA+BYNLKXF+ohSbaGm+7tfo7odnC/plMD+4ivOe13IMwns4nkrqmcGy
MLAuI3sXEFy1CZxeEZkUBRA+7dPWUaTE8eLIkjmUW0XVfS/+VVads0hvitAeborPEpr+bxBQWndw
m2mGbmXCCMlFx/bkau2gRBedydvI8nGEZEvxjI+EIVnfbqhb9hrpZsb3NO2UDaNrPUq+WMKnDy6i
Y9McC13o4Gg4nUegeg+nggpGXubkDO2V1Oy756GOqwRHfrRlNp4LUja2VqYzWNLn+aVKKJhxcNgb
+A42zrKVAXR1qklziCj+tbB67Y3yNgM4cpMfPijDt4c/yORFC/inaFenrUgtRVfVZbyIgORbYkA1
1C5g+x1ALiUbrUeF1V9vwIuD6zATPfKW3GsgP9o6On7FlbtROo+9LfuhEGZE89wUbW43lcUxIKo0
Jd0ZceX4D4VroOOMcvTTMbOSds+P2TVePWnra3E0xBxXkFTkXLbu8FZJYpEcqZO2GvSfmz3IK92V
pwdnzpA60u6+eA8qk+7GbcugwTf5+DlH3NlF6+074ANYuebIZFRGRdanPe5ijkq82kAI8/HUXasc
h2g7RTqDHqoUYTGXwQBOcGCAveoFd4z6UcGHuvCuU3hJmOKCXSm/EA4n4uoIxOJTYXseluR5bty5
w9jvIkdA187OdWsOzaJ8D2aAw99FbMpN+1XPS4yI/erGrHqHEXgR9jtqvjasXwX3Drcw012Kv0+C
KvJ8MpzdQA8n3Cx0LYDvmcvDVae2siaPgorRaup888BSgKU+/fNuM+Q45TOiE2ll3eLsle4VEJLD
NE1Bn9B+jYGiBAniS5vpqduPE2etXS0CK/yXqydeiSOX1wlF0NQLckGEFSd7eUey/JNW00CC6zGv
UrLnUOjrCgj6C9CcCFzBjd6Y7c2sCJAuE5Xlx7/RRo9WGP1LTdU77P2DghSp8ttDh+GEsQ5iPcZ6
YJf+JseGGf6vY5ExU618XbzAXf7+hlTAbCZwSTjOtfP+kMTpX5ZwujHCph11UMOx6bHTbTTZpl07
bJw/Vpr1nJ2IFktVxYdR9RH6C9aZ8oCo5DIRCAEaFmgQSyGjJxmwxlleu3sD59XVTxVkSl6PYuMM
AEyobbXkWZeVt/JyRhKwnOazKVa2TIeWX0f4ZzYrjTuvASkJYVvpd8Cz3P6BJJRpWnuihFWsHIyg
AmEB65Z4Ve+BlUJD612KuPZva3X6zKLdRdmXVU+5LPascmtjLCbGAXgbeQFKlajzjREcwFvR2QQ1
+zkl5UsJYxmA3BiZINfvMi7JHyrK9XkXUyzq6i6Dq5lDHCvEuqM7ZIw6OrKCoIm0XPiZsYiRdhdj
Z4JqjuJKJBKRmLNh4M2WMB22eY09orRdatjmROUAWtOqSADbzgq8MI2Tyrsw9kQVP+pny4gl3sYw
0UuxoNuWzfbyMuvTK9e9uwquJ7SyVUu8JdWpfIfuTE/jAcmks1D27ku8bG973je/U75sxMY3Dwuu
P/ecxDxmmwtuyBzMW7WMNjqzKuB+yag3q5gwcasuJtMUFiX0/aIPsEguHkTlNG2GabUQSrGqjE+I
yjpmmpExi1gCvJ1zhiolkbPgedFbRwD8VW153rrRohQOrvEPPLuoTB7D5iF40SX2IvhBpkkNKBrn
TQA1Vmd/1GS5r7EaiX1GX4hpR4GVlGCRuW1xbwrdHoiV9bwXd3rtBjMpk592NI3PMHNzB0OUpxhB
ZTrVNFGa61dXLjAM/4tUXesV2WyBX0PndKpFHvaSWXFjfrePAco8Efct+f9Q3egmDMwd3aXhKR0A
2nW/JLsjoBiMuUyZ/glB8QTnXaPWAwMbfNgg1n1SjRGURXX0Ew5M3Pqj6Fc/rT3mcfZHjRgSmT2p
8ziXfyAQ81OuEc+6OtMXizQZEjCpLQeaNnte8c86KYy9BKuCEIGXTIr7MocsFyudPmlbi2gzkLHj
3UecmFNnM8SR+BKLVmV5c/Zo0vWkHRBDc0sZfn+M1eZLKP8IpaX64kOLfTGpqczsql2gYYb75EHY
G3W/4JPz2qEch+1u4u7Gdy8huuyjOS5HfRLi0+3jZicnIx3RrM/+69VJbOoQv91eENta1gvJqi3W
eJuCSgH6jxG+YLyI+vyN8DhCQbaHlt81k3gedpmWwLDS5kHv3KD3mTeuTD6yuoTS4CXYNDp5MrqG
KcbPHTxrg50HtG8F6sl7gEjxgGu5t9bswrL1qwIuPLlyObG4Jc/aU9ZSvdZpICYnEtHecKPrrPmV
bw2RFC2SsR8ef2+ucLhrFb1jY9Rt7h/A7eqboOumduvJBudSGYo3A2NnQsRYJzNQ1w9RuHFONW+M
ShI0uNsNo+yGvVCEAPb/S7TTUOZhy/BC24VFokGo9+/JE0j8yxO3HI6CQyw48s2OIPhLSgDnDML1
VnFpwk+2mSAwvkH93XPu+N/9CCKKM9yZ7PgN9fm8AWtuvDKmxs2SCqxFjlL+ZOAk7ByMs/lkS0Fa
UfJvgdzV3hRV7kMryQ827MbexYOP/eGzIvb2xkZAurZXhYP9pe7dfrKMcfa807KzKCwRPEXOiw+h
1F477dTljitbY9JL8AjNAz6gaHixQ0KUPF29NTvsSI6etsKztFWV/nEHCLO4V6Nygi6zRkNfXpdr
x5CX5TGHckV71wEmlFtVtouur9SMbgJmXn8zrMlTHeEqpDewlVyw0GJox8b9erAFfXMDFOXPh/b6
nVT5r/ESBbgmT3DlvY1BqphQZb9/KuQmOE9MJD88dq9WgM9p/Gp+oASIbIUZaMQUPg951Cn2oE2l
eFLWdd9vYZt1iiws6lOqYZcsqS37LwQQUIZIQofHZ3jk8NR8I60cVk46pYeGFL+TdnkmQZSeCbNj
cKOeIXGOVB023wTVAFKAiCSUYLcw0Fz59JRymg27l3GscvzyI5IZDUMa3ViSYWYoZbxX+LpuqTw0
8WWQOUQGhFi6Tlj4wD3c3F6nGUgAPmrxZr7EhxM0cry1MCVKpZ/5zj8qTwQ4mXA/gIj1W/TuePsx
l51mXsrk9V1MQAZ0kpY8gPdlm4FaoaaI0OdrvHTs3B+e7Ld0H+yRUV56e9Pn74iSaIQq122uuw0Q
iMw0NqxTwpw26PLZl20CaXma7oecWbwNT+vRKp2XH0vpANBnm2Zi2f3rdDHGn/LOLPOKEnx2HkDL
Zlud9GtLlShTpzlQ7nauDlVK/uj7qP/GXWQKmglrmPCTlsTfFPGn0j8IJxR46ZlydOL6cbGiOoRq
xlgWVGw54dV9FZL7bAvTkOHkXdRajM+BStE1QWbrTrGgOjlg3ri8JTBktiyWUr3/+no9M5bETeVo
jK6ynw9QXdmkiAbBZGxKfLZySzX9QZi8Bw19fXXIc9hRB3dT3pFcuuaxO3qIHgbRg990EV6tkHSW
CNc1zmljOOpKbEq217MKAmRPYFtsfShRg/nEC2CuGc6VXbWtYvTAdQLQBJb1fZkGNEgDWkkyvPtH
CNx0s614gXsfPRReOfQnubbKCbuUk00wXyqd3QVMI+R1xc7GdsSLhPX7Nx0qtxMd86wliaVOPuPY
DnOP11/7CZxTc4new/GN1isv2UiRJIV/1MVrQYHs2HNOLIXG5ITygcg7V0p3+akVMEqetAbCE8j9
esHQFt/fdpOzguibF6hI3TrrB+fmCefaIlywjAYqlf7Xt4T/2WfPr+CtDeREmE1guLErWszaTVax
fyIIlOaGnsr/6frLK3E5r2TJ7onG/2HzzJLS3cR/gCuvJG1nWDRVm7eHJ07L3B5cVS83evCm06Qv
siADfymbKCmpwd/1CK8nzdbL/XydHItGamf9EBKW6S9lEfP0YSptByi50qWW+s5gNS1yg0gRLmVa
0qX3D7fF2gYcIDteW5OM8lLTGRrgds0bhOX+/4nZNwShVp4NsPGl9VL0MrAkWkG7w2wUEOdVvTJg
2icOVcqDIdN9hpM/cBolPB5Pprr2M5OnXOFzSq6pIz2O1eeOtFtdOBQNdMjGcwrtXSjgvIZK2zeN
bZK11xfyEaX7xtT0tLTYWbEFnD88KG8jvBWiVd/KhemGbQGJot7M9GvmhSh9LTVj60kdor7WAAMS
h7/OPInZNM2DLlWKEa1n8A7VGY2oAn5RhYPolJvf8+GIhDzk7sy9tgXkoJxe2g4d+VqodZXP4ETS
sI+9eMkylzgPG2NBgsW/vhrE8mO/M5/V3ly8VG6/mA4mD1avi/eNe6PULZmhx0yADtMQ8hX+ZHEd
kG/RlFNJVnmxy1AqGpMxVOUDF89Y4ABJV0TYjJP/8cP0pnY3VeWi7mGzikUw5DxEg1kL0peSgfbq
444erNPKnlJfywLxSArDSZoWpvUndQ8DEXCHbYM5wF+Au98qRVuU5+sO/OLifV7V741sc5kX0uk5
VF4FM7qjYyY9oxl595CEtP5dmyRnUWYYyP2+ebXz4rzBgDuWDR1XmcLuaZDjUxj74ZL7z/6NaCAV
1uAKOtGzsJUnWwmpTkNQZSoZ+yUmqH6pHZsG0g8hafRGJ3pUDtnPfBktBIMFwels6ToKKRNT2HBT
BISNlnY8MPmz+mvwIBiUnIopAtA62SiUhmr64N7lSauxAtZuOxGnyEdB8CcKeexOAx4+uuJvKshc
LRqn/WDjb0a6A87MEzALRg480T0V7NtEjzT/JpgbHKOs/21d+Oj+TjEBPaX71h0lzut2L1io48Rp
jjODwvHs0ZWYFjmGQwyfmo8tbDrE0RGW+OLyrqPxWSF4Wo4Q4sklRpp/XtxbavHaz6JzwaJVe0Iy
2RNXgVSrP9UqeS3WvA6YcPf2CZdB/BDSjttVwB4YcUBmnYZxAbd4chARQU77XUnrTWKLxJgbeec/
jYYZm3RPKvef0ikEX0aW2aYIf3C25yfi3Xt8mFseCDY8VA7QnJ0aD1g8162uB1k8rq29+nyyHOFe
q1XG6md5B7/cQGI39m0a32AfnnXp2/CSW/s70myjGA6Yz94jXa5vtrwVuGZlB4JZSfNAucWTWN1+
YF3R2/X977/RTQHXMEID73MaUNCzsYgMVFY32hLoAGxSk4+EFXh/NHlgweGnQSuzK6OSWacLj8a8
8trNkiipcMci7nGjjCLJNnWNJAnhALzVk588SxdE9ijQs2GvTCk4jSEOQZitYfgoP5gXzEQgh95G
46m8gLrQ0uhrfymuSPjYsZggHKJE/Itk8amSaJh01lqYUHaIW86NMbHxTwYgb5ljclGY6rkK/LMM
7+P2D7zvZYpLyd+p5ChHVKaoGq9M9d2CniCTGjyDjunETNshJCdGk6Z2iBGvPsO3+FPr8mAHwXTo
foF4LrVzAPCf1wuSkDgI8dJ7IBiYaERXwa1plC3SLvbIyyMoRiLK5AEY9Us1+Tc2Akad/+9px01g
ClSJfq0ruBDLvuyHs1RhkANOIS9BPXzMM3eOQC6eNeKGPhsdgIcybuturZKzk9f5BIAosJVEWgSO
qd2sLFjlJmI7FuJux3LzMzHH8MrDVyQpRuPG43CyC7fd6ja4d0YJPYn39tKzmPFrzmnd/zqq+9j8
plksb5uBHRoMivNUrzyoDM7mgjmQ+S8cDxUfIdzevDh3J2KtOUoaOPAYz0wEY1t8JjF38qmsS8TL
ledrto3lmIQ9p4XGV+tzXmpkfol+P26lowgGzGZIx6z/t1JDAv6YVYoxbb/VM2JGLMFO+JxTD6n4
PA3sVCxR2MDzcnFsy2GWtqScGQzesTptXuudCqLOLO+lHkFBXy9L96CWmZm162P20yNd4Q5kIvyO
CnCvfUO7H55IH80VOoK1KFaU2NvFHIfLAlC0Xl75h4E6smSnVG+I7MswYrOac1Sew6cUav/E54dm
D1pSP19m44EMhPfZT2DZZpEHpvbMx0waV1BKyHSlTRQztohZiYl34iCv6v4vNBXOiUj/XDVcJ+GV
1KFz0SZTa6zpo603sPb7WaDaeWbvddNnVB+cZ+I6Hb+z0LaoVbZyuXdudnb7mT+Ti2b5sxd+njlv
rZn01IlyBWOGBruHHWl7jmtg9SKSUK01uFRK+64dIDOpmh+lpF0D3q7/SK1CI9Mp79tTyknmsw0Z
D3o0SdEpZ5nQQ4P+W56Fjx2iZRJQ74nP5VNzXEPLYFQ88g9TpzNFF2qSxPfJoY9KFYLc2DCxOd4U
kfrFQv9Gnz3489zOBEcPEazbcjhf8XPQs7oz1iNW80ZffhnJw3Dc79180NiPxS8bONQPsIjKoc4x
Kvp5O6eIBDix1EgvF3TmjDvU22rMWsuhiQNQam4Om5w/ZMdl2/zE6KMadlv1dYuRnMXM5LykCQGS
aM30OSFGuJBC3pMV+nHoiCbG5ktmwa9mvB/Q+nu2CkEpwrkZ6Hk6GdyDHz8sw5TY91W5cpMyGC0V
fakrYm4o5l1SLsJPToVnOxU1hC0eY74GIpZwlNC9HRPYWTgS945O1H+WxgbothnuQGCPk/xMbUiS
Zrm0DRRIak5s2aOYPUchaAOPdR+V3jz75smrRoQEzRMAAp7Cl3gJYyonmFtfi7Cxy/02TkWViwyr
z+SCdK1zloEz5GRa8/YGyS39ZKaIkkBqFSeam76EjxeBEf7oC9zQgxYqUQ1nT8hYDah5DdyKU/lS
XoK6d7MrsU2rXU3jg3qB6ze2r93fE29P0+pzVd5+ffiotFdkejI7QHVkLTXjnblzed7IKJrHd2FA
svsetc0QIcWXa210ZTgXkXPEdUAFLC78DTeIquTAENFPbJ1sOwHjpheDt7QVCsAvvTIHmUif4o2T
7Qd7/2Tz/6Bei4Ay1ZaTiXTP/Qp+GNvMcbNdEAip8PAX4Tznax32yHULP7hFQ9rJc6chb846PlGJ
d3E720jHLblVtKFI5cGC0OWwj82FhUieGSNXuJAeMTEuHOk7s24wO2WfM0YAHb0F5DF148y6KFzv
7YIqHOWNg1Vzn17s9Q8FP/rz52xdQptbNNnMNinMKjQeLffzHfYLVAaKdzVbcB0qzbOkjIiiDKV4
8CzobmBBSmHZRH7dr49cWKZZ2h2DMy3IwFg72kWHMlrVm40wHVSsxWxasrKM3j4Sn6+/gYt5WokY
WV5tQrrEQL9TY3wZgClPiWuou6rUyMDEbjo6Az7qijsIRbJi/0bx/FFcQlI3b8Cg0qRneFIrLier
WNTF//paSXdIrfTSFsufi++ZygBGsqV44PivHURjhKs08fOEsH+MZhbn94LqB79a8Jium+VoODAy
HM+mzGlDB9WhDWvrhIhdN4WD1rsIciaUK+LO7nA/T0EcP690KcBD4BY/eF3iyShbRfmbabc2tuBd
wfnBBweTcY0J8tYZQiXNsoXePxU8P7+1gtcW3osb8lotPyxNma8gzWzNwUrqR/D2wIEdob2dHBw3
rLxEulnDKcBBMfJbTK6ZinT59bsP6c8WIwcBoJALbnYd6/Wefv+6TH0sGxts4wNERXSbaDVMl5Ig
fCTyamU0N0eMxZs5tfmL+tfsAa99SqlnTwiC4t4wEyiBeX/VhHTMEhK+DuqSzKpze3XbTzVlI0jP
w0HcIMV9NqjVWyiFf55jK97aSdX7kpK6bIXWfj+0TBbZF1u+ud1hLBFzq3kctlV49j8ymDRsCdjt
2GFmBmaqcJYeikt3ABU0Kjj42TzX7NQ7Lrm+THxueOQPKuQMYiKW/NfPI25XTySsjxCXb28+1YBs
Dil+0DuMRe7w3QroXUHp6+hxVFM8n3JP3L5hmZY0GRAq8x4AzGBVbPXzR0ETY8woAJ5uezCx54FK
h1gSmAke29hH4qgUlh2XVQOPjQ15qe9bSqZ0TqE74BkY/1njDNmJoEuBQNq4ywHoy2YzxEyKw3Pm
CPDJvsDiQi/suWGZs3BgI6FPNbUHdjywSveaFFviz+fsfHHNAZk6xUcHUvvcmno/iwf8DHam/wtD
x6dyVI2PCQniqyyznrawtncqnMWoNSM/JGQ5bcpEBDTDrxIw1gs8hid2WWMlvDDQy6NJFTP6KhHm
fuOjMlIZiauH+xMqSBH7WAAG3PuyFAjmqL/R9FDNKGfoYDrKtcr+ukOw4HXUMZmnwJGadBb4DRYg
H5OHHMKFMH5tPaCw5h9LafgvPtjBDNf3QoeacIM3ZANJoLbjiYBaj2eMl9VvZ2zXcjH+QA1+wpyR
7OZ/c51ws5mTgjKExm5XK93Uwz6eHTgJKtfiXf6PEupOKCudednOPeVpU/SxnGKUbN0iY5F42y/c
OA8kxRmt5E3NzaoeNE/N5R1gs13m8jpy+4HMIEibCBxKSjhwjXCEgjcjVQD8KyPacyDl47OTPN6z
QsANhqAgAcLsURRCwzSgUnOc5UfDaQ/2Dl60mfAb5qe8J5ZQ0BmWtKCHVXSc/7sFz1QYYsxKi4lC
uwQuf7XOfbOp2p0CrBcxPpXp577nLWZ0uuHy65aMftj9TDmtNGhQS/SMXCti+vn5jVEXXlhsJJrL
cmyvrYZLWnPoM2o0kuolXM0uI4E1exWUvGjhP9b7CK7VOY8MCxH8UXq/pveJ4vQt6iVPCyGkyiew
DBkE42XTTqyALM3EH3sNd4tl0LtUJaG4+mj+TbFZd2x9JQFoRYWJyuudnMYeOXCUlXHajCD7PSZv
/q9wU6Tc102YepBbcZS78xeqiLLT588K6mqV5TeEt9ROnCXqtpbrEyHYrUsIPeFCtG5rOQOy8P5Y
iz5k5DFJdhhkUZtzQ9pDbVtNT4DEMVJO5efYrDYDhrPfaczGdl6S43G7vms4nBXqR8K0ZIxunrRi
95ibZwKix7fJazxVd+sIBZO5wBB49Ey0LwI6dEcKcGjj4eWYZmVcjyJgbmGl7LIRmjodb2MLxv8m
Oa0euWXnPCUZyvjsJzXa1Av7VjRKEtrwQzdJasAdEbUyiUuYqtcFSuxbcJmWjWldtOwKKg4PW6EE
itydRgecBNgGBPkm1+19ckwsI4O0X2zL9abR14spIPRhFwKDU96LcvxfBY2XnqcF5d9UxP7Kb08B
d+ppYHgdfqVcoKbaK2b4zbhKNdOiltkYnwDYT+xjznnBh8KkxxrSkSXYf0Ur0JrFed8CGnMfy8iy
NaLNcViDST/fajI5f9/pO29JLWrv0EC6mWMSPQKKTpjLmt6Ux92vCqhU0ubvwTmeSdsCb9JtypAk
fesgpMiUEQ0gAWkEFlbBTeZdtxT22h8GXW4593KTioQi+u87bxMMVS3aWGgaQngJ9Aqnp8lijwSL
oZLyv8QSH7e87Uarxw4Z0Dx2j6rZWRVJRUm9QJzOfrx+TUzg8F8faccX7p0b080Z335ACAGkVkXJ
+X5sZPZurt/3YCZNiaQPq7oKe9a8NBc5Et1f3NZ0BEOw4fiqG31xASMjDYdEbJ/JIq9szkW83s5l
akc54ihEtBPsBYk8jA7q1f/uEaomhWo6qa3NjuRRshRHVqFqk1yp7DdPe/eY+fByvSw+XYkw5q+m
RJq64Pm5074MPKNXpznDOFafyQmqV3XgfF6vN+p+rkwfWsYLEUYq0NWAX3uJqPQqfNe+EX/VtqOY
Q4zlhUt/Zqm4aeqiVKLev0FG8hHy7zfCnPO0e+XPZ5Q/zgLJXdfVo5SsZLIOK66W7rOu1N8t3OP3
nKB7e49x80qW1xoO8Orqg3TeneFzvrWwnnIHHWaabgiEDL1oUYE6HAgzADH6j6d1jXuf4C/I3wGq
UE/tB9b4MkEvmfMCr+fwa7CUuwMskEVhLkwOJydxGqLOZ7hVByHQu5VgMSP0ltxTpLQMNJ80WZUu
jZir6MDWop3VxaOFc1rUATN/hIu4KtMfeC6sN/mdsGZJc6wDFg0JIOPNLE4ifL+VdfDCgDus4nt1
5MTLLDmO3twPgmT+JH3AU7Qt760UZEWECfAnlZ0AwjfyJ+IT0bH0tsUQ16Cd7MkwZukDo38Y5roM
qsQCfDU5nbCtnvQQRG+MmrN9Fz/+iip0HSfMrtUzQpW6wxpeRFqTC88EQ0EXcOnSX4QvUkUz7A8E
vsOJxtEHMYemWQd2We44OAehQAg3J4LWGgEW8kyL5clvZ4pQdEqUTpFDY8xMWE2NaY7Yc6DOHoJj
uk7heuJxPknp0kkFpReq8r8K2VPTERvWwUf4LxeUbdWM4eoGMALKIpLHKkFz1PfG6uapOAbEjpRd
4g5Du1ASAIWoJvnq47fiVOg7AKXK97HUX4kyiPav61vbXsl0R0OKEm/rLT7ETgZTlkBTS6F0m/kO
mWtYqdnWe07N8tzWNpi8Y5Mn9xrcuAoWiVjz2d8EN5VKdze5qPLr2JVPSTK8Zm9cyEFydRUf7Ut9
wiwXpfoK5JdZLtGIfx8zcC59NKpefMtzBwIlILCYF0Y/Jx6FAHMmdrjQfHuqvtNkv5zMekC/kaH7
t+lJFWmDN8LU6wuE38Y8xMnsxjrXPJ1MggWUqYT1+MyGxhGcY076UOt4LyCg9qeWgsRNiZe/quUH
m7zXEQla0BkULNpglUJqfbrn4ieBRrTVEopruY/twoZ7d/IxGb9Gnll3Sns56ugPrd6thc0sSOb+
8F+kK6An4pVXy9CnO05vC9vSCLyilqhWfLx/xb4fDKpIrvyMT+d+7ORjLT+Pqe+uCtZvX0qITTN8
mzOn2yCUiWwBkrmaAV+ejw1WfQGB5O9z5RCSOpx8azZZCj1ZkcSAQaxCCamK/e6fvuPbqfH5f31p
6nqPLOIsnk9+mvUoEf0A4GB/elpfBqslvHuABUQYSPVH/RFhMCxv1Jy4fYSKTFCVKp+8i3E02mZ7
kXpCUCk34ryznONZrjnZx4bFeRmVQYA9+C0FHXixNwqonncyZmVNU0C1OXL2T6mbOUOUJxDfK93Y
SIp+mXRixlAXezmLGwnmmU1K2jpzWERASdZ2tQEsDhWGBxed0Od+5dpBse4OsS7XrMVP/uHKGPjr
8LVsjBaHkHD4JTAqvv/iGbLuXBUljBN7GXWnc1lqtRmNmKplA1zElv8KPkC11sNYiHcLfs55aOLd
d4uadRD7IJoze4nMVHuHUnGXOVYRE40dYLs/vY4qNeSxzOWgPPHEJiJKXyhLCVt3gUxR9JDLAvYr
OJskNzQr5GS8AGZ/Ov1b436g722OWgJU4eeHzkan/uwAR+BDcM4rULmg2ozK8jDymGCyRS5nG2kt
EmQqO+95oV0W+2/5D2u7nmmLTOdiahhSK6dbqtSFhPMdbLqlhlXZW7o5I8kIIcLuB5e9v4N1dVnK
RnlDh9dlxJ246iDpenwDpPueanBndDwOnrj/lIptitUyg7jxsKT7ZfCfOkxD0zRlZUtwRHrYeALA
ovDq8mNOq5Y6Py0zYo60moUa4R6aUyAwcQvnuYLb15/HPeSqy8T8VTaTOwSN9SjuhnNOGLt0382D
VpmUDuAhMtMNHNz0Aomv7mUG+mFdmjGoir4qEpaPbh6yKzaryhyuXJ0mOgdDjxQwrPbPR+4YA1v2
KnQ0YPZqlKA9dC26FeGZCHWGPgDWVpV9JDZ4DazNi1hV0CWg+y61RZZDtIAKPFncb2U1yS3taFYn
JDbugo/aVhf03foWqr//L3VdgPf9tNHZMC5JE42QcmWUKCRCrE1GdMDxx3GBJGHlUVK2bRhbs3pk
qLHCv/WSCpRsExJNmZd1gOgiUUlM1fGEp8iPiGyOKHQoL6K10q9EJI+6c3CJcUYFmCHV14SXT3u/
4yfAWgTpSptdK4Ajqnx5QddoULkVkHTwWNWg/EX4jqESdBSTGmJvclyFWfyqKp6qra3hFbzmXdYK
3O3eTMor2o32WSggbXjVjWjUHCpo4n2Xs+CGYlmAdGKig4EnTpliBDcr0W7Ezw1eH1XyV0Y2/JFH
y++fUETCPOccGhg1qqZY29EsPHoSYfjBtSYgW4RnxW//fM7Uw9VpLk5GX5Oh+q4+4b9ofNgAPWLd
454WFmqZGZCv1otJ6lFrr2ZhN36lL24pZ5AohG4dnFGz0owGgal/bawwWIP/D2QwmFIscRQT42If
8ENfnxKyh4KyIzHvMWST5i3L94cgKOpgMYuuz58X3Lg+3/pni52Vai7l/rohvdJJmyD8bSHAHZf2
tu5GPTwd1t+pyd+NrpCK9oK/FJYqm8WP3tpLaAytiJUOPtbqESj1jiGyRms+XrgtmHuSSp5LpwAU
+6bQGsdMLA41Y1fCu2Qi2vPCo5HGUaPx3pmrpT43q9Hhnnqhf1SiT/cr0Ay547SAp8Diq1V2j15v
e1lXKtGAmv+XNf2UBwLkVqXHXmLgCuUvu5kbphIWGZ1PDUfTajhaFKwZn35Hkx8ozf+oSv+ctNMk
FOHmNhHEHZYzemZQLD4h72KgLV0XC17y0P8xdHSzR2F64/9V+AJym8QEfrop8TE+EGRyUG8ohX+S
GdKAyHIzmNrci7/Klta15ECA+aEDps3t1msvt0tCaYQkZXqZ7FYdTDKHHAHnIT1nVtXpAq5sUxM7
HDszuFuwRLcg+ZnWGjklCrisUVhQnvSE2/TGNjA15B4+KGEZU8MfgsEZtfu1ESCTuy2xnL4pJIRt
gOc1x8mvibZEpQP4FaZpjwp0Y/wgs1s73w/y6DC0OtU7Ykphh1/SLt+jE+6TxgwjxRS5eOi3PVau
bwHRyYU/0nMFXS4Ave3LmUMslnDpzETlioaBkcFbh8fzzIKgvaty3EPh9A8RywnvmBniq9ow2uwT
H7goALJk6q+jEwU71FhyxfmhUOqo7PVo/RhHCTR9fwRLh1UVAODrFxHw0IRYVZOL7wXvujN640Cs
LqgQ6o7e1uKPa1o8nde/vhSyNr6ZSlB+sk5qB3Ty4lJjoHAkut/SUMI+f/jZ+BtNwowiqRJntVuj
3WRUAkzxDqBT4ZIxYQetPorLb8ZI3m5KyQurgmUiLQakPzP2jzmxAcTVEkfT/wGMk8aU5cn5xjiM
zJhXLRSWSmlTxgPBvbY6eCuYBTrWZR77yiXtICkEi+RCnn8PV3te34BXyPx+3HtlluBWWo/PAvo4
anKqnkTJ2pnuuHstFULJ2u5TVUo2tS7vtT5WXyPehF37UqhijiKGP1oa3VBWvwBBoC9+AOjrAfZA
ey33pvoKzZMBl4Xd9zfqnO2ovMnxqP83q5Jzr3/zGGQKhNuYxp8qgiXJnCtvmO4Kp8b421ZCXyr5
5griCiWNNPb410795ygBt0dENEtmmhDpDRV0l8Cb3D2kpcwTv6oK0chV9jqKo6f5z65EsJjruYY7
drAxNn5NeGhK5BqmfjIBYDbCiHnnu6lEi/I4KXEed+M5fY9ukZkABP1LhPZJWD6nhJ8CwsSY36g1
OBHQNvHpLw01Xdk/xO0xP8nkY2hU3atmX+3nDVFqTFfDU66XsUClWXJy0JaUtR53cBU51SVGAF8f
kdM4yeijUdARIPNoKxcF6KgOuTv8WJpWKhfdNCBRZluCP0poc1634IR+IBQ8HdypC4Pus3UjfGK2
Ad43Dk8Z2Uy6k94+JKLoYDcVWPOKI8hQ6VuEg/nunAKHgXrS/7ZSCTacivmUvZPjo7ePBDJq6SA7
dwzQrA+1dz7YwIJ5TY+D8hEXs5yiA51z8hsb7OJ5mKcgZGqaRh9VHlCa8zYI2RxWm4YFGU+ELsp/
b9wYvS8ZV1LTGDHBG25E8sSvn21U2fAUZyA2I4GuYlWW4XA7p6lUv5V6U9irpvet2svh+2jpHFpY
GWKaCW4+dpfDC8HjecWK0Sm14Zzw5YI036c5wRBYW0z2NLTSOSEcSp0gYQOXsm1pF51bxSz9XoXm
ewP4Ad5W4F8y5sOfdRrJvnvh5dtO9RwmkJ0Vv1qA3e8WHa0a657S/ANKWyJv5Aa7/jD0a3gTixhN
dwex085Wf4UcSWNl/kQ+oieuPrJlEbXG8mtPgRqUs1LvZImkMnaouT+9M1xOBquLfZ4pOcgjxM4f
3afKVYaMVylawrV7sMhlenQ3Ebh8DlKKRiecdmBe+6rMxfFE7EvVpOsS3GkmpCmLNirmg7WBRcOf
+OLOEq6865459v+50QjqfL0dZyTSCYn+tGfIm6B0NNn4Ardql/co12rtPvVemr2ynfSHNAmAzHNg
PjqcDdrQchXMBXfZjLjTbH7OYsJEeOJ2Akw3kVLewRBXZj/B1gEiEz/uJxZ1sLMQeXpUnX7N+au8
xD7XNl8hDSS+uvTDJhZ/xgPggBSu7bk6LqG59kkQsh8NwaotLd409lB6tbX7SUtCql0nvaH8hu1x
RZhxeV/NaRekjwBAMeo7MSmB0n9+nrcBEDlzqMPgj+uTHudS+9GiavO7lQv3umQ/U1IiundVCEsh
s2F6CeeWtG4W2WZwkM2G4QTi+pf4gM/THxLaXfHfTHe7psfWBbjtnuStXl16Ffxm/kfNBHGr6v06
aOctQeDwbngcqFiPYWq1XKZ2bUkK+/K78UUAn7ZtkRLGAEdTNLWmZKD1vJxY9uKTfFDn7z7W8VKn
yshj1CzhuoVQrhf+SYNxGH9/2Tgy4iTfROPtJTasgq5um14V6m2ZK0V4iWVn27csT5eeEGhBAgaV
fSM1QsyxbhmomFb2nfX/kvjnVsMYnTmIh+0QGgTqf7RVtpSk0lKWlvYn52P7mN7Q1uqbo+LjALds
brWwt1NL6dg+9zX8c5skuXI5ckm+lBEQR1Y95/451K9YxIbNPBybuMG+X++MR07SyXAMaLf6if7k
oll0FBmuEaK+kxxePiuTZloiuV2j/FQCh8XKwH0oPUh2JMmpxta7P8aJk5kHCjtoZuWscF7ZrO3+
7d2w31oj9BzVJrNb8u08qx1MbwJa+3pga8oWWDY3GrTLnan28Edr8uIYus2FzunwWH8oN0OMvQXf
FcH/o0Kf/GysFpE/8nNHkmzOE6jlJKOrRpeX186aQmOD5J7Wixi1BXGueW/jDAng4HD/T9/5vpaR
3PoPqR6wAOLAJ8hE8kvHOcD1R+n3CBHaHuTskE57xLcYyZpSGwbmz/1jp0mtEwi/Ph9EHAa7Bemo
NKLpG96KjtAGtE+8xY8qB3EGQwQ1iKjoyD6hGy9ToU3uUfSX9k9FKS8Rguvx1HYJrRq3ZMK2qUZi
hRoLQ5iyNbq8c5rJCeXC9kSm7XM7TeuFJcin6mKTJ/OFoSb9EzpkIMP8wZMZynRHlzzzSluAEiot
ZPwrdCCcDLkDZB+1DJukl0ufIUgc4DdreVtzcjIEsxHvlB/pX/uckjsKwAHgfm8LuYLVY35s0+JK
HZprUXC8hDhC6AJEXQ++i+qrFbLe2AcgipewAFtgSBfid2N/LadG8CI2gB7ZMZKAJ6rzbkDvRlxw
QTKgJTB8LJXqADiXjYjSifmoVIt1/O9xsFnmm8zKDf82kMPMHRVn0St9KiSWDp2RO202V/ua5s4g
7Bykej83fn7tNhveD79MOcLhHWd3jSB237XFOVxmWXKMWi6ju2SgslTpVwa+B5q9JXYDa6K8OtAE
UevuXXzj23csR/FX1kiZAgzy5RZAhMe0+AyQalDUBMmN6eZJ71tcMm/IAucpvzjC37bkInbZwzTQ
j4MMrHyly9RbrBExacBKddF4XzM6IilRWDfK2TTcPmYgfnlQUG1WnYIDNyCTBoS5SnY2L8pcZzhr
T2qkWFImxrOhBGnKJ5cEMPNRt7xiz58+rHc/vxZASwTKcrhj8v1FmZ+Eu2YzL9PpZOty1s6swoo0
yLVB6viE1VPsUbBO6W8gYm6CbRHzYzF8Pf6cod9zH058+g+oCO2A8B3KeeK1S3BDdYHyXylkiskV
y9S/odZYIUGjDzu/ApC2QITcPT4VqhZ8U8MLcTjaql5lM2CjbB7kOjvzvODjKQxngkRR9yKfD1WL
HrOmmXsLvm5JFRLD2nJ+J6wwelkCmDqci6PLeMr97ATbfwIc4+IMmUC0etymNSLPvEQoRZORhyO2
EbJLNCs/HXC4qvNgfiZP0dzBsfmsHHl718MshVvi9cLrJzmyDwuCNnJ/eAgqzfqJmwVVIs/lf66x
DKwnSaUDHLXGFhFbhX69DjAA4wNLfxVMgxf60FpGEb2KvrH2JMzUszPRpxHa/rjmPDeD3u3b3qzc
yIBVOszn/TAMTIWGGxYGfLeBsvbcb5mfhRN1CtV7WlwEG4A1i6mxpGMiMNzp1W3D3dkr/mYcfEp+
9Q+mMCJ16LC7Vdk9/3AtKa7t6eGE88R9Sr1JFOi8K2oUMneQ0N7M5t9AW6GUnKVV9YfSnSdNr6rl
wBCTvX6OIpzu7GzQ/cZ1CYd1M/2L4DF+ZSNmsY0X5Wqdn/+NyPt519Qtmo9Dicz4D+baY+4KB57s
Eyo5QitdZvFXqTgxjfdeV7jhEqZT1ZvFcVaOxjx1ZUn2brYxMInVq2Lmq+3HOjX6gsLAOUYAIcdZ
tDOjY9vNIDejgERuN+wfpowgxC4Ooi0oSsGo4ux/PldcFnaIiaVsEoZX2gImRguUIRO8eYh6iM7Q
npTGJ2D3HRub7xrEm1UCCEH6suP4HAmto7RGe22EnUKm663/VnjF1Atn4VP9makj1+MI4bem0B0U
Q6ieKOLUD8rEs1zhHPea67qFbRPHZzI8XNBsosQ8Bjyy5RUp/YAAm5P71b8h3zS8wStQbdhQvetd
YrMbOYb/dtqs7Yfzw44gBjS3jvoG+S3T5GBpFRlZthLPuEBiwJXi+sXXdAtkCEHqG/40Jog6q4CD
DjJw+zAJ2X1jum/dIXdywN6ehR0iViSOlKutGNZ5uMqIvi0GY1oYdatkiF8I0sE6djLUcAIKh8yP
LyseAMMwNdeaDDQatVMm6hW75YqEhx4yNqRJuDla5UKBMd5eG64MxkixJeMc56nc0d5IK08YAO60
b3zfTB7WGLW/z2ZCF0osikY2+xHSZbNilAqGM9grII1SSe1aFkbEwyA6xma1ulW3zwbnPaeOIs39
dXSxeYKRrcHW3R+ooonPIEq84sMyv3f7VTNQBkBSRP1yLbpKdEhcTFBEt7ctmrWVfAsj6UZBXH1S
sxNz4IoOATv18n01UrR6EYq5SDiNcC+wapAgFlJf8CyJ1Kgjzl9KenD+yEPd/I2+hlhI6PXsbS+V
+zkheBNvJE/g4DXim2gwJxMyEVjlgSwq+fRwAJ1cCl3u/xyzURQiK3DbegKCXOGTIHkMULsgskm0
KjcIvrf+OIFTakjV7tZpjIrAvDlJNJUJYyjFcPir/1sFe9jHO3NIpVMM/OEIpO1RbJ5rJcMKnfuU
NgNiPovtH0pIzd2/r/KEGNEpQSkM1tIFV0d/uKjg0KrRg+4lXH+UoAggIwJEpCt38Vd0IHoaEwUJ
cqWN3FHBLY99DYSbJDE6pXE+SSMD0TNv+5g6J7mHHl/KYwA1DYdswE69IvoH2DQna3RLP+o/7aa3
fT4Ag6S6YL6uF6ZY7obNYdSrlr7QtzoaWn4KeozT+Of+dnBjMFO6NwWxKaUM1QP8LJAl3XNxhqrd
Yz8ww6W1zd1eEaCYOApMajlJiYUTTleG7UwI6vz/i1ySGNWJlP8RJVxNQugXwnWpML4zZoqqSWCJ
gA/C4iIIhiSU34HroChj59BPJsIzXc+bTISJ3n74XlllJOqyrTgy4qDO87KatHJl/aifdNjLDBQZ
lMRukxwga6TCAq6Ia/SGs9gm9JXPEMvXu3oULUlExgHgUy4C3uJdnMMGv9OVQ7tQSkpnHSKFwq7j
3Geuk+xIlbi26CeXNEktrAtmem1JOB61Y+KTRHx9dji6Fe72w4nDKkT7gQUD+iVGfd+ZgQPbaqSh
0fbtU5i/lXBwe8W4dR6JOKWnpWjBBV7N0+r2ZZpcxJrlBobMDQw/DKPU3jto1aA6oiM4YiQZrRFy
F3g7b/ScWgsPJM9jj6WJ92XXYmdT36MMYZanSJy5USrlYC7diDgGMWocLXRC5q5vIGb4PZwM668S
jIEc+ZR0LisL0/Y0pSk8Q+GBr1+JLAkzB/0JMLR/GCTRJJ2FfHl+yuReRXYveCfHrbY1xoKLuWsH
Qp72DhvXyxc29RrreKrgrfEVFikxMd6CLwxx5mICMOnMab7TJba258QPKOrKfQj1OvKnF4ce3tlF
3aNFAldriSCUGIj4u8rtmG+sXkaEPy3bnmnNvHM8iynG1D7byTiORrZoyt51UqoiErE/eGt51VK+
YZQxFZvRvDetiMelDzlh1iKImrIVGPy46oa4vcEtC1eajFB7RTUlRPmkyfNyoXNrO0+I8YqB8bvN
gs5SxxzPUWxnV8DnNecrK1f8eLLbaH1ArxMtxqDPEdCpueRY9A+wZ8YStsR34EFho9KIKeUH11Ci
inlL9O5z9ERRMODYrNHI/XPIUZgZcK+hMYKocnnYoSzppOcYrSPotmbyueYfgMrqWNEcB0pVLNd1
LANwpCyEc00tgy1NssypTaYIjCQTvLIfLSdZogKdLFWAXro4DEsFE5dDHj1C1TBrF8qPC4MDF9g8
cC0Huiv/SwbkdT22dk6NBJKrT/kJMokgVrkJEQ5xtHOe3nwiDzVI0uOc5rSxDMzs77y+85hLb7mm
VyXptw3PqzhxIAxGCoQ+PPQqqFqBxhiELFEMKF/9Gnw2fcFGDSiPIcXEhnja0dDN25iPsPo9xH+R
rGPDAyqHIZ5hH88qR4SgLYXM2EoSbQNClFwWT25HRXaQp9nlj0/YZS8zsH0AdB55O6LOtaNvdoRW
FOoQqP181Xc0bjm1ocXG+6yb8BQL5QH3dOZKwPi4ucfIf2dxeOG5GWv9oenOG8pXXx72HCVbM6Cu
1/hmaZFVkh0B/vJnay88HBpU6EfDuvm90A7iJC5ddawDe9+mjwFyPH+3BaA7OdzCG2g8RvWoDSzJ
QlIYoi89CN6Op1s+temXNI1XJL7tOrofnBAmKOk2qS3Itwag0ig13GN95E0Ig7qEpprZRNckmbgI
viQ4VJ+k9ODfc6bga3DaEa9jlhLMp8yEcbVUAGRVVvdPR14OIY4QXqMhH0KW+ZpA10xEObRYd7yY
WrU8LbEgPKfjon7wzLXw9KhElW/zM1fqWJXTe4yZ3t4y0r2eY7P+S5Nn9PsnVLUX/WxccM6VNxIq
DVWsE+CWyu4YVfOBt5xPrJNVHGRn07V4pTPz/tIgkY34WFmJC6Vx1dH2mmPTTrBFRc+p5rBid7vd
xU6jh7IJKvudAVSxyOzIKV8NmRTcLDv5FpbbtFA6iqG3lVn4e7CNfP/NExI+aIVKO9/ZNUMwJ0k4
e1JwLIbaqzdEl4DB7pgZhcVPAHA9vsKkBjNreOImpjJsOdAMQWuUDJdTPJeGvpGUUO6CD3ndARZ2
HYgRsSR6iN622LUt4qH+Jtq3B0wfph61W/tCpaXPgr2lIJbcgJ7yXQHZ9cBJi+ZsR6TVF2uvy+Mz
QQCwxG2TAm4iexwcDDVQNK6P5gsfb315ZzKAVD0O3rOSSqSGA1blMkF5nPkZTBh2oC4rZR94Ro0B
Yay9XwFO6NL2eomH7sWe/1G7R9UaCymKbHyQXtnE9z8/+EwoUacwVOVtNO9DAZq7UE/EuMMTLaID
v0WljA9DRhSrLhYYflnotD1Yhc0o6wknbciKCIAHCXhwUfh0W4fntmQSess+0+6k321mNGyafXuo
bCqmh4gAUF5YD4fHzAKV/darqywpIY2PlxlaA1GrVHnWvocSXBG3pPz9M2dKe7xido5lwyCz97WO
JkT/mXOCOHxPKG4lhm8hvS4lwumgp/WKMP53v3WtJAc/Bb2W5SLIKLkXJFeXcXURLY95FMCc21zg
VjB9oajRvzOutlobqaCHQXWPABAT/M8r/Z5QB1N1g/eBssZai4ZGhVeY8gA2MbVzb8H7vJBKWZKg
atmPnlfNDX8qzP1kHYPjsKNve3SrLlrXl82gsxGxXScYjtB7sY/puHOu8tmN3Zjagp7qV1iyOS8G
2v7LYkjLrN0LwEBu8akj53UDDk/ZzmloV+8oAmU8qSlHtnbQGnlBb1uGTlofqcYNM9pAmrDByxz8
vwN4/B6kgX5Px96+CAXkxn5GCX/toZg0iNKHyBwHypR9GKSNAWXyug6HgOspEs5573J5nPUetvhT
ic52nuIH0pKrA6+Bq7WsLEozlcOFP4wum5tw70rKO2LgnxKvzHQzIruq77G7sZAQoxds5TBuYXZm
ReJCGE4m0log4pvrliaCDX+zarbLA6CCcvf4MooX97Jz7LRvHf/e4udLiM7VQeRFX7mzVs8eyLHa
NM7HbRTe41OdUJFmIyJFbFsu89gdjMTdopYr0TFaVl+OC5sYOeCt6BbAiTWr4e8C6q3KaegTq6uw
PApwZ7DOkEuczeF2K0AbnJ+Em0cSLgtH4meuPoZkolXoI+eQF2f58PilM0B3R2W6XYonvPBuJdND
d8RExb5dVS9Ie5kFDG9BgZdJwIk1gd07w22Q5Dnz65g2OZ1fcUXkuRdCPkSc6e9Mq8spd5q1ixGE
TwWyeFOs/sqsEDUvieTNOXy2DQfw057cVIom3hH1IZ2REquIaAoTA0zJ1MJ69vmMXYJ5g8BcDCN0
iM6d+9lq0LXVv9FotjlOJ+44VrOukRO3hupdUxtxz7c33EyBNlth0ee1PxCqAxf21GKx15w04hZ8
Z+ZHJemNU4UsjX8JzJ8OClnteBcUJ0HK07sOOoccp+VCrW442wvQLjFj27EVgL8ozUlCgAsr/LeT
AhGeOE0Vuxslh6SsasGBd5R3cm2NGggwT5WQYZWd6N4IA1ZYev23554LVk30DF3AriZC8s1Km+kl
2xdtCARRK4cOsg9ByoVB9fVrIDGk5D4CviqHSGT6o3HX9oL8zKafBkzaF4EE2en2SKNs6MGQFlN5
mYnyOjWmJRyQWRjrN4i8OB5sd00lGx5z0pyJnio1kHlui9Je7MQSSbyygpUp3pSi/nproEBPXtul
TofbgRo8y4mNLDieOA+PNqczoLk5SXGtzzP5AXUyybxhIpvvEBRAnvzxgvioU/9avEq5T9ayIPuf
apF2VIj0WKXmIoQJ/mZN6l2f7Qf3Ysvb4m/CTtXs/rAJrY0edNe3w46Av1pFE7Qrjj4g14xb7VrF
D2k0vRcqqv5lFrai1gM4pUUK3SxoDYXLng/eyeQFhBXrqxTygTVquJOibnfK5KpfY9VWg5PPoVsn
VlXbmObrcKKXFHsbmTp28fOweXog76QPcMmNhYvXLOIJs0fjW2A5wp3QbjeuLvNIHJNVh8bfIO/8
7TryRJy6vVvYb4hysijl7uKvV18UzStFNX8d6+acG/nMNsNpXw4SobTt8hUnjdCQZ35PirjuhoBM
0AihBEKGZ3hBQl/u39eBsTtiUUblH0BBC/+TDY22cpW/4QSv9y+5dY/+CWjXdxePp3jJKpD+9yCj
lp2WdRnoFHhSSlVx2sOdeSPKVDxc3+IwXP53br89ZpP66hTczjuDPPUD8LKZnteaU3BtTR3rsjQk
rtgRdHaCUDqIvUHstmYydmwkopZA0Y5sc1Xos9pwUihrUfzQGoW3Ugd3v29UXkjqp0sA6Dqnkkbs
+8fOHKOGwV23/Xf6osj9A1kUzhaIR9IndipdB6xoior48a5g+qURW5fSaEHPzhZnyBOBIskP3Mqu
90Iai9DUGjD9edGnn8v0hm25mtb7CNzVWTApZ0VtlZPHLzYVP82EC7MKC3gGCWk5RAlHNELIImiK
E1gpsJ8ovuRZsS6kTINRF6Fy4VKPgr1wtESCUqyaYErzsaO4/yyHI5sSwpewC1PlN+RYKZqXMzOu
r5O00h63/szJKl0aVs7sq5Y8YuOS9OvdF0npsh4Li6GigbentOCSU3v3I8wqAXIi94EQ8fRTW32J
7IJR8N5ecXGq/Zu2arJH49wdd6GC9s7oDMOdiIDkdhlIvp+YO+hUXigNeybvymQieQydLWdfQRTs
MlcOSKwMS4rzM0AYfWVW9HuqV5U5n6qbPHLMU2U+29cwlpetc/5gvZxfYtP+T/HGY/yAqJNc0YAo
LaAOb5ceGKYVPfL++lduUjWIyPuKfc7unaTyGtCMvBUlqf0IqYHxOQ+IYxn/OBLUgvd7AVi1iP78
3oQ8DV1hKzauSpOi+a5AsLPteIA3gsBBODRyWFrab82RpD7ILhnGFd7XKrrvvASt6V+9o9ywHK6q
S+D10cWJqAWFehycgXN2cJeTdRolgc5ef+I/DTzGqrh1uPdelCvEE/BI6cHs3fMFDNorRmY89AZQ
6P9OmB111WiIWpIZNFK3oPAKBE/S/k8GDw8khUwyWA2SnFGPzQQP5rGshIULFyHaEl5HYoTnHznZ
DlIe7FpYMn2qTuPX0H7BinV+CfiPbiUbZhQn6LmmpaWFIlnn66yrEkJoWcqTjou14PSiHoF7rIGB
8DD7d9Z2pHdEIgviZmXE91PXsFcFgUBxFdTb4h+m4MKF4/hWZePqqJsssUyyTcqt7TIRxGjfescR
57SCbIRVzWxzXKh91AtkJ4SYENQbrUSHseDkjUWEQTSq0OqZaOJJWUHoa/R32LJjLzeUtkxOoO7f
QNkULyrJqqvohiCfMN4hZQrqNdiKtcaGKCPvry3onmF6ZQBV0vVpug0W+GV5/8hPu8s3CIQIt/AX
mwmvaqy9s+fU751X5+SzFlVCpxRo/ti32wWQ6Z/gg37eovK5DGYItkKnJH89NMrhVDHPRhgisVXC
dhJ2nraK4kgCnf2q+vO6TAuvmuQKN6ZZrCMOBZ0AyowcOzHqBQRHWth+7B1SUuq614ejJvUQDqMm
Ukj5tOTPIM2JL9L34ySmUUX0CGjc/NuCiZJFdPxqSfJi9ZoVn4+Ibei6F7zlRFApvkcJTtUbbW/v
I9sSRIRkAo4orNn5IRBKiDVjs/leZh0l/obwP2lomrMbCXW9p3FAZaI3SassR9S1QX5+L3gQtLu4
bEJl+nfbiG3xUNz3VWLHQNuqfm7g5ELpzRQp/bkrjYxAiPae74vEbrjS5UKu4V/7l9lyc3zUgf0z
GWdHdrworI3O5qbP5ZpRiK+b8irhfKBkNqyYwS4LWU9hsMsG26+jIoy2WVrAeQtHTGrePz3qxs4K
yr10EOFLDgKJYNneVkze3n2Nf+LIQI+kt5m4cgf7FZJyPosRX4fxgcpR2Ngx9imQJMHvcS0NC7dU
TLKbmx0G9URQRCmZcfPog20iTYrAdzZ06LVe0pDODfkqkbIP6rx7qN81Y3xc57j+M73YGoVW5gy+
99uTrrM9lBTGzaUYe1QgoOTH6uv7RDX/qWRCABLIUpxCXTV2KzVm7KaPqExsJDpVQWJ+aGAAP63L
Xja9HAX2GQZpl7XHhdMnXIU619M/H/IFEmeGqkTfO7lufuP2KuUmiBPcmoE8G5ngqKN4dqe9Rp11
kSSgfTZLofejErZkn2+SP2N7DxW6FsLZiENG7bZ6Ikb2diDQtFqS562mJQwIi5/u9eAR2bWckcAE
0RuG/XilDw7zecHritk9ILjvrLD7pLhXTJYZ+U1CbFRvPpc70eiqC4O+M/4bBYMgeCWYZ8smO/PX
uukGrUau2un982Fy4D1J7CJhxRu6ZPANLslH2mqypDA49QwU7KpPxAS1PQprU01sPflTRpJOT3nE
0EX4YqVGIOb4mcO+Vi9zdd2/knSm8/jUnILpdbAjknIi3vnw7cfytW7bBWtTJihZ8zdQVJ3E765w
rqU9EeD62ij1TMWzC0/RjI5TRt8UH9TyOmsrpOH7K6pvfb9KmHD+9L8KRgUeswp27rOi+0QD1fVg
sjj2IkXp5GLK5lJrZbxYR7PK9C1RjkTvOZR5blYtLelFTk9vi7yijPw7Z6OCVcrf86Z1tSffXEhF
yGYFuylTS16WGkSL8pa4y0XFk0lTkIhrq1zqcibxqkz++1LkRJQmP5FuiC3tECp6NyljMFAemxoi
4o2mbwEHr169pfhF3GNPbK27j23zL5608q0YlGb1QMaL/NJ6tJKXy7KHdb5AoQA9TPT0YdlHjkfY
ExQmwolmgXHTsEZO1UdRmaFRdRwihSeXU7JnasVEA3QFSOLA9J6o8mQM9Owuuce3kAVGGVfi2UaR
NMM24/w36Noz7364FZlIn66f4vG43gcsAu+bpm+cTA7eA9x7NIzigxM6ZwI8QrT07hz8YzDYiSfx
P06R+fngqPFEyrGEPiO+YKhSf7KGdoNT1i01LjKu0/FUC5H4Pd/19+DQsHvPNyfZ6szIikl26dgQ
ReoPbvC2t0n0oCyalxQ7Qd/rgEdleZNK48ySHFOrBg5OUqk5QZ2/e3hzrxT4cVAZxkpXX8FHMHFZ
WRgpHe6UepztNU2eu2EPOR7lhxINuTPAFIcF+DQqx6m9n10icHmhFKHOovt0PG0Fq0hu668f8gO4
Fby/9s33uOtCxMqbHh+WR6UGtfHn5Yx0i32b8IK8Z4Q4aLfR+2lIbdDPolU/Vim9JfsIN/JnAuS/
fzJLwH8gBE7/tBDXRwg0Ny8bJtc2zIHOPh6d4KAgQWclmMpOP/AVOmg5HtrcHrtkS1xXPgkR97Fc
BC7C/LHPnWGpPM+lR/rFE8HqSRb50nEXq5UVHf1mx6Xn2M/7W6EBA0bIJS9pUNUKrBdA+hE2SmJv
X6nhXfl9iMXpBHVz2eOAjOobMxdGuPpqjxg/3jdMUfbGr7z2uICXpBtKUXM7qA7IK/NVdFUnxDpv
UYdxwt4lYZAMosyuufTv9Rry2A4Z/gSH32FgUnz5pE7lyJXNnbiOye4dD1LA+vMA68sUxJ2YPUSw
BnN7lZUmjsfIj35hMB+pPCbAez5QpgLd8XbS9AdjKaSv+fUWo9vAGLoAdolcc+1pEFIlcuCVQZ3u
Vhw4+jqc1KTWIMaZkNqJH2hU5SmVO7YW9iA3PNmai6IryAlSYbtYvVLtFSYNOEAaCDPUIJkJlIpb
a/g7oX1vHdg/R5EjnVq0i45Ph5ayLq5Dd3zjPua2JRPT2N9gv1AIjM0evFfLavL9Hnu7hyJ8tXCP
unRFO73X/qSPSEShn9hJKvXdevmfR1zMPngx4m+8QVeHoBlSwPvhpRUUmXYNS8/gzQJMh8cyGvDZ
6hq4G8xVEYtVLMUSH/HdpgxmrixTEffLPPLNLRBZPsPic9JKVTSWQO0qTLvwKM+9NruoVPJpxRSO
VZpeirmJSNg148pdTMEW4JZnFD1LIvVF0wDP5spFx/ldmOUowUqifpTtleYrkBPUH2u1cS3wDKm6
faoHACVL+cHfswve6zSH4UMJz7uLsbCqYRxj6TOu9ZCLDA9YJ8mcWFry99LMzLNl1oc66uqLCer8
dQLR33f3tz8XtczWwnEYVUU+OOmzcVY8I59oPojFspywiqU0sFXHfXHPd+TFmdmhUwF/lrNRvNaB
YWRvWyfmKIiEcNV1sKxCaqvVSVTYXKtuYsrhrO8WcgZ0P+8HuhOUnfhMCayMxeoNWVuya7m5BXi8
FLDKqfTv9e35ztdHtkQorkOOezYZvoDzwJ5RobK/jbI945hZZzLg5GXvrnp4nQXyo6HC7dyh+Xso
zQLjOAFuD7Ax/W/4iIOJ4NX27llVZKDaFzzWwut055HJ8hMjJsuHG8tBZJGOPKZX3mKcm/NnubWR
mv7MGwJZ3wJsPVodMLdwOU54oKcGh1fDpWcgDsqkdCguhDXv579AJu8KYlMbIoqvIXFrmHQLTvh0
y1gk/I8PG2wT3+Ei5dyiqKRrJTO89UZl5grco8KNDN+GnVubGlSPvfzv/cauCc06d63x5XRxuj8I
8UzMfTkT+ZzevHy17HWsu32wYelQ2cZqonwlUV2rCMn1Kr3yAD0wZQUtKQ7r2HY4wYVXsUnZ7j80
BbQSynGOJnDahPRhN87iMPx6T1GomNiyGkq8bdydFlJt5OpfgAJcZbt3SybyzFllsKnqjXp9f+uA
ruJP6tPXP6ngb0Ug7TPfUMvVh+Dux/UKFOX0RA3nnfly8feBtyIJ21TIgegTcF9ioiOlKxsEGKV4
+PklogKosr9TJ9SV5QfifCMuEWa2wM6X/5oUBsfqGqMqNmtEmW1XHxuSMQyeNXsR0V+tUfcPpwtb
MnheNijCoRW3AtHjpuLpvcqkwb+8YglFCw6fp+keOm4vr71g3B2rAKhIrBBbtY9Up/AeJPk8S/wS
OxSSB3Qi8BlZ7Z/q5UbiaSNTv3b1yLpsN4XBpMFW8vyBPrx47q1j0fNutKVpdj6doxnhzHMfni56
mtiJx46IunqgO9hy3nFpi+R6azUCGY4JivFBuvtX2N2ezUNxVT5h+IPM203LOdLC9OHmV7cCChHH
dT6XEOMs7Ba72UcWG7+PD8Q/m3BjtPqV7Tl+ksbnmO3yah765MyTcbifVJi799PZ4k3tholnBSwH
7pPsZ86ZvHk5QA6AUIWLx8gahaDah93X9IgW66pCzIp++84RNv6R5ofRxMkwGbBDTqshwxg0o0kB
m1Zi8QETD/PzBLDU/KAkm0bQgz1zTQXgC7niX8IoIra7+1JmMpAHDjwfgboce6cuIwIfi7om5SlQ
pDrWJh3a5JA6/I8SrBHk4BuUK3xlbrhRvBDyum22RNKEwKGsAKY+++8OqwAp96LsAVkid3DAdQ6y
98C8jwsBpAEwXAqMcpBD6wreWRbhZjW+lq9uSruLGuvShsXUVf2iSHA87aqcTT0MTSgdsjpi0eWu
sWZoCuZYfRvEf+eh2Mrl8PVy+KJcoIcyM62LvrNZWQbzb6vhK5IXR/ak8BDreqLBgn8vcfKomX3h
jvPnc3VXyszxpORENUp9wbW1MuIHKTkHO8os9KLGGHwL4ETl2ekDDaMKoalsPRZcngBA5mfWr47u
zNrZAe2yrRU5VdzHHrdGyEBvhuQKRIIQBZFrVDg51vW77CKluuXpjr4xn+iXDYcGrSowUVg+m6+4
7jszWu8qQ6Nnnf5+ZGqWVZLDcnBchKOGfXxcdfPzmf+Jx5TGkFRwB2u0KwkfISgJyGlCitCaqRkl
JvO+wWVZP4KLbO2G916aJRBUpcxtfsl/lxocgiakRXbOdUOljgHeYIjd88EJjY+LroOzbL/FDAIL
Wrf0ia6A8haqofmq3yEfTpVjBMVDUAUg/WO+PgDJcSuzz/f/VMEo5UFs4wGb1/pc3zFItz17dtTX
QLIX1jy75BX3T/m3M3cuHb5WSfXf+ANLkCzg7Y48ZE5ncNKmvoX0c5IF4hTMg4p6MU4mRJqRENZF
CWNk2QfpRrLsWMWlmt20kqDNVM4tNuMvbr7l/baxHMalkYkiNwx9/I9xMqpetwyWThS91owgPqUF
npnz7sESrwb+bLUGbjntiiHb7KD0M2u91vO8LcBrNXwrMk9vNBONezk3N7nyDQxn1pIEJQyjAOmP
gZyaWmpEykMO5yuRHxRzeOkNrtGMBsKmq0qZ9Rt2451qrwWfXJ3DNaQ2D7JZq8j0Q8WGla6Qt5dF
SUQKhalEARPv9aEBlR1X3OKewoFMI0Si2S2D2PFBlzn8CQAnRhPidWP8SjonLMHmIYdUGjc4d3p0
buCgo2PzDgQA5fBMY5hHXYo0MNCGQOzpPZP1eIviMumhP4LVqRcVaxfc73o5PRe34KR5tQmaOjB0
SaOqnhjgdIuxBogtJyVNcgxPdylKIEHV9JpRKqPuZMOsYYoFqAGEn+zkaa5ydoh1hjTpUcvRKOJe
8qprMBA2EjHNmk4ND5Bx0bWcMCZP2CYToNuKYIhDZtTOrmQDaRgsPDm7s1C8rF92Ulnq3L73lcmB
Mv8CccvR9K2f9WkMgHmD1GoaXFfbLYsn6B36HvPMJbjkO53LCMB0PlClXIf2w049nL5PkFEn6mLI
k+pY88gg5IlueYhGij14bfQ4B6Bd49QGc/THXxHVls1o9QnDBcU3yExVZWKcXeyX05pzAgTYjU4r
jQSmpUH7IxXFHfImfdRbQQ5aG96kOa9/eT0xBDqkHhevLMz4gf385tFUc2+rQAoHH53SdyMheu5S
3hvKKUUAXWENC56ruYmDSxysFzQ8S29ve7kQycbalYF7O5ThAQl85dk6X7l+x5UB6ehcL2hYQsrc
f+HQLA8TuDHP3N3jY7TclV6jfeI49bhkEp5AOk78T2xr5MV8F4rnjMzMMG0YiIx6or3oUvpRm5o+
HbsIrvSXimEF5wp14SkWWD0hjhVmepIyDbyL/2G0mns4r7UFD8d/F+tvyBaD8IjdSFLxzuljKv6N
p93WPV7EzTMo2vGm5B8zQP3Mh4KjAdmpXKodqnKC4A4Hz/NFL26dDlNfh6DxGhzsE/v1v2vD1vMN
WFfwbmYNsFKbwvEvjj3+vn0+DpjC8BrTec76qx+G4tk/nIxqwGA6qZeif+fJq4gd+UnfBGgRTdv2
ybMnXu74N8E3jzXp2VaHJNePl5QKWuvHc27nJOHpjWLWY77d+iT07eVSSUegsF+ZVCrCFJ5ogYzp
Is6ihVTjZiyxvhYWjVKydmx0Veoz+pDvU33zdar40mEivGJpqrkMPfADV3zywHqKf7DAJ563gPxa
SL1yDsGKfQlCPx7TK7MI4txVn2DF3hck7XH7isF3hfN3Ado5qLH88aO+Z91QadNLNsIgvctC2gK3
5GBM084wk0VTxiEWQViaQ5Sqq9oUkWoBZgPAbjBWapsTO3jwDnWQ+hbp7HoTC81j8FnwQ5iN7qTy
T8X9Mu3tjjq2c+2KlPH3h+E2RDIeNdSCQWORjJhtdDdwHza2PX1Ppx+SmeYEpmlV+wCEMfNlEcRL
dBxRxaqGCjABInB1udI9+pJZHb4QXVB73fn/8eMigjcNpWtbKoU4zHyOJQNv0KOivGSZZ4juf1dn
ipne8Acu728zekkeXzk+U46DMXl4m4imtg68rJACtdnaK5haJfAMyMhA3D6Gf+GEFR1g7PxqyFOB
2WPI5OhzQmibMTvX0hIe9JWRNiBXYqG9Bggwo+5Wa3ff8kiQh2ROOfWb+IZvqXUbAym0yFqN3IOT
SLSROG0ocB/XEkIxiDaqBcsSGeshwVeYPYb66ASv9/jVC516/VOGk9ACx4oKWfQjDqQkFDYMj0bx
jnl7Ju4DhQ6f5NVTaVcED9Lx9VF5w9BQiOyNA3ZS4y88IkdlXwWc3vhAXwPfIWaNgydf6M4uHa+i
wXxvX++vUGinoWqU+OgevhFa9RyqA3YSlOMph/CtiOUhGILnt6MoO92Db8OL0hcfoD+JSTqGpLb+
asuCOUnlpwfi39PAmLRpYrlLSSKkqYr3Fd8EVvWnjp9AmJsMPkxnSB4wuVKkWjBHSvL00tADgOB0
RyTbRiZhooy+qLQnEuabtRbLnfXxfzUw6etm/tIKZA5550pPfhA6HlVs6eQ32+j2tP/64w9DCwCd
U5aypU0/rUxV0P45hcxbEMmGknaFKaQa+gg/dsGP1S+CHj2vz5imZwj4sQnSAy2hTDechTw1jO0y
P8JFrdg2uJxuIGYzg0MBXGA5UPUg4W6NEO2hQOAwOBA6BU+49a5443uw1wfqhUQiTMplS/1rBW4i
TT2glJfdIHhbv9K003I1EhJfljTxjWCLY1/62CQB5B6MULaG+Sguj6CHnzaASGqyZ64qHtaGBNSj
E6k2Yh5jJXg2lddOQ9J9ai+mTkJfoywG5pox3wl5O9zOuHr22MG4pyzcdEoMlrE07LaAo/U7CaKj
sWogB6U35vSVfcQ8/uCFGkifvM57MMOXgrJOr6mM5rgk/QTACo4Emm1Vu056aygiujKlqwHo4cTx
LHab4k+Cv9r+2wLad9FxtnUhi+5qnCc2rj8zjmPVhjAgJnmh/gotVq5Ce662ai6q/OJAwT9OcFTj
leYIdIFqSMoLx7SssZAjUUirYVZt9KqqPA792Sn6LXfkJDyqgsc5bSeoqBDzQ+MHkYwK+L8EhaYj
WBwBwOy4lYrdA4bBuSRKmfSb5fqAArR/E7zAuWTtKSjRhyDdQIDswP/QnJeFCE/xXxlX2uJjrEc1
5KP4Hn0lHK4Fj5XUw7U9ODlCUe007o1ZOFom/nQpabb8trMz3O/7T4qv6VWJdCUKifXP82tuKed5
2Ig1kHJQ4tyvhE6i3wiQtmhi3vFg1xxoOqy92nEjXcGSvpDuRAYfs728y3N30hyG4+hiwX25AXO6
iv95sCnv0LyDkBYwp28VHxU1iNEzcwNsceCKIqLWiZnIkNyhrzbFo3LWahA7AEtdelWXrZ/K3KhG
Z7BzAYMcbTOZkapSYog5nkTvCSFQvdKDrUzbpeqX7q6b3tgRGGSjWrbNrv4kMETYO2S64gfgo8hY
SMFfjQVM5yPeckZldRIh1Xni1ciIDc+o82JqLqZdEHMeiNBdMeqM4QyPl3cxwzTSuxCSqV219aVk
ANgeTgW9bEJJ2k1qgfbGUm4pNrPJzR4vLY98xuzLEDwVgcs2JLmXUKb85jVHNP/yRulng0a4mZc6
lvOlyXDtFNW7QIL0VvW4KQSdHULwe3dMC8DCFMSjBDdNSvtqIaxJAQ3oBLciS1DiKke97v7yfThp
mK8RThGwm0rDF/DbbvpIyVcBt9f3pZ8WLBKmmkii5zdBiFhHuZajWMRYIiXR9W7yOZs21whIws1n
3uBgmiO/Z0jSgjOhcMNMDT8GA4lgNLt5lCquHLVlJC6GPGyJS7J09EkQFeTVqlENPgDWLH1FJn6W
k08WfMvp0zzDszZo6ydVCmjxRbhjOPCfA1VHwr87CvCQiFnLI9V78blUhwKp7dcidRPHEPYvY8TC
983yPSAdaE8fJmNXpHArF/KTyRSCE6ynuM6IU3r4CwRuMbT1wFbpsnTakt2hr/7dbm1t2IN8L1tR
1o2Fsv5Tvombl6QPckvhXuzs9R9VyHESeaR9ewmlc91BIstOJJtZLQ1bMRgTuTdmHfrNlNlMs4m3
yofVdixdZ6J+yGQvz3O6uZq/HJWrW3EUSpl5uXODyLdRydVByWJEOVdFHvZPFZ9We2taKPSiMmsl
Ic9TGIgterst57ge9qE2IU2upax21HZmq//ZDQ6mZ7Fol+sfJ3SPS3tyy9bB5lKq9kN15NI26HBj
lx/vBjG4JodLzjcnFC0w8v/sWwdBHvDDjQ5gZMFeUoJU4p5y9HFQeE9lY7s/BT3g6U3H2VTH2Ggt
1JIldptXxrm09S5EQOKuXLRHRqzlwmfHhLilLTjSSdy8QZjg7OmkbKBHGXfHK6i9/xp/+uKWupoa
rkEEEywzXN/LWFyaFAwt591UMKOjB3X1alwQLAfDbcM5YeA8BxO8784jUosHkCf7V30mqctao3sR
kQm9Cn9rCJgYNnfj8+rLUtoFm1SWYjB4nbXb239jRGDEi5yynaOBzov7ag+vimYAb/W6akzK98YQ
x+RICSV5SvUiJyX3p+yeuqd3f6qy6IPuuF4U/UV+cwqjQZqu+eRfw58vZDFGu0cMXquGXbXJymss
HVzHZTYd13sTL7VkhIAgUA+a290vcgxq5NDPBB4zhgwyUSYCtORnHnx0SZ2bTE1lMomQ/SNjsTC3
olSJu2m7ImpZMb5ZrDUyeHuuaUjscPRxUzE/kXmGXnf07LCpOzZTZCZmri1yoXZPSe+g6js5XLoe
BUz/mAPRXvhfaEHyN9+AAMjCZJC9h+qKtr1qygCMdXgPZRIn1hr/as+OpEnS229fANlfWx2Fb/SY
Zu9lEwsT6dsggI6SKg6a27WpS/T5LjYsXpxn7ryMYcloIYtJM3d15eAePSjmFSTry8RNPCDYQrrV
e3UxVq2ct7Kwdw7w0gI7En5+2tLUDaIZwBwNwXlYv9j2lLpPjPvEV9XRg5Pa+q+q8rOeAq4zWcix
cQfCIzrrggkXblYgP4FIUZxvP8YgzTqucO/vUS/dtTCErE5QVaw9FznyLY639S5KAj0diAevIQlc
qrWhLsYwXl1IyaXQ6piFtos59AJ+8l89QQ7gL9V4SYoUPDTAPWNGnoc4/cfWPYDoX8g8Fuk8BEp8
BiwHTFNMdMSb3b1m5X6KjmFTRMsnaq7UH+dCnmpb3TgzgwBuNHAYFOTLqPfB6CsEX4SybibeKVsY
JSOo5vAKxwGmtnK6X4IBOcC3kwj1vnn5x75wH9bsg6YAgRvO1GXcPf42lt5nmJ0/S4C10D5gdnD0
4wCEqY45KFbiS7G/tkHyFFemxkUjHo7BcPGOCfw/CSl0EjkD840KR7aPU0gbsRNetULL8lkgGeJc
DoaYb3lt+e9n0uYi1MKurtq5ccOhWtPE1+Nq4t2yi+kG8ERQfwta4cr2L9ghEMmIrMgxrsg+1i3T
PzFJQPCdL0hilQssPLOUfaxqPBl6e4DAvd3QRDVDm1ZCGkRWQF/6B6mdh/ZCFkHQGm6R0bWzfccx
YnC8MCIWvPTdDdEIR+IQ5SzxC4zezSNRVBamYYZilhzZirqStdwpyX9NAxI+L7kQw06KCWcyneAK
do85jRU+TIHBrQ2DrJ76b5SXnye4CeGXh46lTEqI2D/cWEruyH+LzlJ6VxOce2Iz+bwUbX9EQQj0
ST7wwvB12k7I4JxdU7VK/BVTnjkGTLaJYSJV8TA0Twjv26iizn0TTdhYB7psYtPOm2uG/5WEn+RB
9bHb2dVP/v5V01jNTRISFzSi8zKjTQcWSxvV1fTIGoC5ldTrtgLy2S5VVC2n8rjrOGIU08hbvU9C
For7W0hLi5rZqNBTHR1TV2hIXCt8Al3VIJfQIvvCF3Huag2uXEmewNac1MgfxZ/9QHeSa3vW8PO7
l9BzzJ19B9Z3Yu7ijJvh38TSGCvYUJRbZbSi3PrYjlArnLfPfn+HJ8Dlnfog0R9/1yjyxeOuTA+R
3Oxj5Eq5lCdK13vFtUUUiCu0LUctyhNM+OTvSPkwQJsw2OLipSWrVPpagezjF2K3NjoW14efNgYr
Ev23htfqBpP2b1bh/KTabNwf/GD54Kbxz513tse1LVmMDYYp8ZlVy9YCnidIPZlI1T5LrukThiAi
jFKbjUy8Vhl5CGvnYbJmWqQ2YnxilxO63zMWQORoVZTZ3ScD8ZcKREoLUpvlgujK3RCxSLW5g0sW
1Na1uxjiotqCqu+EIgpvij/DxrZuYx/lJ2gDJBRN1RpugonilHCkw1uNmvDHumiL3GEN9g47TYt+
BcfTZUnKAHhmumQmrjSqSjlalH7hW1D3QhNCHVQwhFPzIG1L0RSSdQ8NxhR1mSVFsEV7GhYDQ/Q5
lw70T45AHR+9k37DLpW4u+S8pbPI/LTvnmKt4mqmghP18Vm1VEMaaDEqaeHM0QOXVwjLR6n0uJZK
hUEK7KZPu8XAnciAWOzjTn1ZLl6mhq1W36OU7FO90kkV7kj/dkKiwJsyGTkcU/wqACxAWxKqfhBI
7t1BjBCLCb+UwHDygUt49L9D1qoUuKZQyt4Q6/LKjxuZnzn5LB1NU2u8faeCUDPOwanXq8p96ncT
89M6ZOiKsmsRS4vQkTSgXm3PIw+7w4hZMCxEU1a1IrK1Lt0zTOlPB8K/tcKU1zYzypQvtZLiSNEM
cSaAAmX46wiP9Njj8H5vCp/FP+FeBpZdgUC9eqEj8nfzmCHCwEtKNTk3dDS6NOY4yMWSWeuLIH3f
6RQF7IGspev151uIJDavI7bkxANq2ZKQtamLuK9WiHQ8Z6OjPkCRb8Ov75wKMEFZN3zzjMT9j/Vq
zPvLFLVJzDZlA4Kt0ICCjfR7wsvsNlcPhxOqh6pGUaBhQYECsHNz/eAytWGtD9pwcaAfNa4ah7u2
DbCyqIC22045YemxdZIi29Tku9drknAlIAToUVEcoqsRF85JBs3wHVCF7JwIvFjM1j+6Uj2i5QWx
CnxR5BpKuGKMGAo2T6uwR472e1ekyqXe6jC1i/0vgg6elU1pmEh/icrCYWRNVYNWuM+XpwF3wVS0
eXDFiKu1iOEHluLvM5QDFiTqsHAVrr0jlJ9wOnYEtqgQZYI9+SVOJitTwHFZCLz4ca2PwcSUgjBV
QvqFg+KXqyOBNFYBGmNcwelEDSeQEbuO/xBFZJKTcQuvU3fu+Tgy1VCMeqMoOQbeJhOKktuOeHU9
hXbKTM3+qbBl7jU1RdsFfnHuvjTGjarkA30f/aeigz4jK9RfNk9ZikPrtkIwHQ3r1z1uWgp0B4zX
/F2lqksK6QoVl6dSp2Q/YoUkkRjfHrLQ6j27jhYXnosKD4Uh0O75ZSXjFah59NkRsU/z5D6eQGYe
eDfmAlRpSo+8Lnqgav5z6IiwdTUjz/b458dX8lU1pMv0OZITX4QjG7karZKGJTy83Ak43HeH0xDP
eQqfPdWKzRy0KxjWqSFeMhzQ7hUpc0XJbMDU3l81qPovQnbdRI6R32E/VNKLCSyu8ojr/Bi0cFw6
w9aB8uId/SxjFsTLpn/yrU9Iu7BeHosMimU97mV6xOXUppslirC/qhogSRsy5vgPqgmQcMK3yZ5q
iOu/puLv0Ytd6u4gznKNP8yk2OCRh+hd0/pJOf/fW8qkRXWKkWK9fMYj08yAvgrH9xKU6yHfKm9z
6pyqtMhobk9l3leDDPLJ3PFj5T796YGYnBZviauFgBfoCz9l9zsViUoiPTv5OSr8xe2KP48q4hpz
Dlz0QjkzYh8pBPsJ6Tx7tWJKrNjGD2DnBel6vrfc0bpUAojLczkwLkWRJYUXNXGE1JzmpHzx/Hes
Uec++pby/im0opwz/L0ti+pagZ3V/nurZq6izpLAYYLuk4SGJQr6LwVdkoA5pJuSqhTDx5P5laAu
GrtLG7VgEpIMDGaWq7nvvOYz7ICyZsgAKt97jL+sAhMQTjm63V7oViDEdoBX9SMrGB21Xx7kge+L
Lx1CeM6syfiRSHhmJDPFF3qpCZf2pkhbyorgcLKZPjOB4ET7a3QGWmryjh288FjMJZ98i8d1DU9B
3fHioylTekuMjy5f1qnWQFlDGqejmQE8T/aC6G7H9ymoR5AOw9xmP4VceZSoUMd8B5tNP52cMbDa
FLcWVSc26DgLl2VdOhBt+AJO6DuTb4oXMgDzgDgIqDnv/aa0hK1WTl8MSr3RtxuvYz9p/+75Apkk
5cUbvDKr/zS1uMCSc4qMcsguP2nMkMZ8+YJGRuGZunG9h+LeuUVPk7YoJNVsTiw6i+UFQwBJ1s3p
TxCP5WwEvQ2VPHWemPTsbarEXEZF/Hg64lsGR5cyyYUbjHviyYLGT90hwwshxb5ONBbAFk44JNBU
Sb2HppsBCeFouy4xonezrIzaj1EQmU+YYVB+pEbNNDyFoCgmlD3mYaF271PXuYuVnNeTyzrmnRPy
6tSoHJqAHZT/bAKnDHMUoETeKgmJZZawWOBoOh4FJ2/xnMMwNuiS5/p1TZnLAuEJPPLLrfMCGKeX
liFUxUGAQGDAfOeS9uvz/8qi/txZ5r9rZldprnYACz40tCJesRRVD+YSlDpbNWwMWz8qjJ+SKmWz
nEin53IvrHeJ1vkVs3SzQb+TWgFTNaGeQBUMiJB+I1t3u4piDd1tSwQTjuEbwWHSUky+cZLHKQoW
SIkZVEhmciOm0lPDiXJFn4Rdp4+ez04sPiQWsaJ/Ix/XAfnZMtHgz5/uZQVQ/9vwAWU5Y4fGqvis
x1QSMZJJSoSF4LkySU+aS0FP0N/w8qE85q2uflpg4xHwcE/818ZYLPacp2dQtenNweviffXfbsOx
3qG2DEWGiMNHnTDO/IOfc08IzM+5gOETuKshnCilnI7Nliqq5/iHBkaCeDr+bThswUU3eZr6XCkP
AQE+0nglsNJ27i2a1ZgpCiFptnIyBLwAFlcLHz/YxtN9jwbOFbU+qZkzAYtzAcJ9xQGfok0LbS0K
CgDLe5tILj6qTPhcTouMdjIYpmKnxZYh7OltWqI2N9Gyb/jt97PSN5iv75LBL5LFPda3yjKX20B7
xQmvjP5VuuMNShw8hoQyTbIuapKb5ZdOX4nW2XW9W6OdEYEPKR9Iu6XTH8RMbfcSYC6DDj/Glc7V
CTQqNXR/1hgkwXuh6ZfA163zPv8da02gNjNR+09L0wTaO58TB3/izs/hXcaH+nanbAbZXyLbV1y5
yOZwvVvQf24P+1OGfD+NKCVWGbGxodJD6GaqUGA/jzWaaNUTu6DTyxy8BYL5COaP/ZPykI+LxKEl
yHuR6N4BJfIOnRpM+9fR0bvizdBz1hJD6OyLA0C5rNNJDVz6OTO/Z+uYNDGCjUOJmOw6OhDSJEIh
2pjQmRmYG1nTHvQ8h4S7isaREi7dqQDJ8uD/LvmHt8pATNwH8bfVMA8JnuPclZtYIfubHY24JzbZ
GBdXSZiiCdtdDFdFt5ffYxytir1TFI4LKnhuCauppcFD3DW4PawOO8wz8D3RTTiZ/3yhOCU3jS+7
2+J9CR6H1FJHXs41hUXOXz0gD3no5EVBUPDpSlTxgtDGdPnKJ2Fflqp8+jFtdPuFHJlsMZHbuv/5
j0qt33NszTaYdDCxAUZ2fK/wKv9NzYTWoedDFcGkKEGobadhmHYXfpYJU9Vz14BmLhXlX+hZ6dq2
2OAEtxlpb3IN9M8u3VoXJTXyl/xI1o34Z6Va1cY35njz0+kJL2qAajPirSyhjUJEUyTcJRcf1+P6
SceiZK+b5iKaQHQhkSubmu+SSy+oylYl53SlFlh6yOEjZ49y+roRC26QjGpyaX7pXRGT5rBN+85H
x3j3IvKRtHOu24lYw6M5AYZU59EsXxSNFh45GDUXUcnne/oyPRcGbsMH5t+nXGARmBCCYZ9YKNRw
6VjnYxNBXjrZEDEltFYxAIt8X75Jo94MZ3YZj96jnHYHqnLU9T6hDHmHGooiF0qaew5YkZfSw560
TKTGLQR9WIts8A5HYedYdlLtEOBqet/ZaNoGPehu4+whFsiU9W3jlk6PcbEhlQiR06WvSJtNw4nb
+E31tPqs6dX3nOA8oZIusqZBFtBH4u685J8Ul4eXUqDSqTISstnBfqrbgK14vPEMnTbZp2Adpgnt
cSqesCvIZPFrNyavQPoDVbhBIAgHg4PwF5xspJmA6qhQIdXNptlxuqttKBNxBAQaoltQdzAV/Uyj
PP4Zd3aviJajTIQ6anxxCMnlm+xD+fHWuEeZ96240U6T6CjxoRTbUiZdEHalPUKpj04ROqqsIaAA
+wkWArOb4CHNOU6AGdoUAGkQZcE+B2ZWtM0X3ffWdokTqpO3FGUUloe44seh2JesBCXXw3ySHkDj
VByi3nsT7b6LnGPBKQGzrvSTi/YomD5Rd681bOuOCyaqeuk03xzcLEKnOwaLtwbqX1tQ2oWqac02
07zFIm679EwPCmZKU5DgkKQhCcMwUWnhnoSNCGUIdElmhg15lINwwNaPT+589Gyn9yygDL4YPW4N
fxsr98f/1WvMH34bB7rDHlI4hu3TT9KfEAEtHQWZmhx1XWQktcM8fsxXP+G8xz+mVCvenIE83YTX
XXD2boSLYr6sYKnP0UPU5lYnt7XLMX72zVXltIU2DVnHS9/RGJlpIyz0L1OKjhm5hWCjajwuooSK
Fqj5PAgUL3SrqZ6vBPAQQafGk5OorhUh3mB4+WeyF8558iTtpn0lVjubLUsIBJVlkPIEdvvsX63a
uv7Sv87yj076nRz/b4R+mcX4XmAYkvyONuBqnjO/ST+pfPoF6lDbRwZBrV9+nN666t2K+431CqJk
+nGTQw02PYEWRM+vg+dwuJduALkNlebHPJupZnZnTF8pzdMMkFDS3jlINkVoRk5BXXpsEVS2P9Aa
AmqqiehZml2snlbbNpiiV8oH7k/3VSnjlrjeIFFsYA2NvgY41QJMTJ8kLqrvnsywPvTDhAhdhR0Q
ReXtNpWGcG0BOBlfXK90Ydti1/Tc/Gdh5tnzGrM4BDBL4RCbOxZGp1X2fNKIXY2vG9wxzJ2ENJSS
lMHMybJ8wH3y1sLUmnTvxsoXJ5oy99TT5hhxUxYrvPWMhTH/7vEQ3OZXi3/Fap7/hAzFsMU1Zb1e
mk/jP7gThmYdk4muyRDfLElBflf4RqZO0s49QvNZ4CRU1n/2xBkRl54k5NFS6eB6nnJV0R0roh9Z
mEnpkBjE6BGapFNhUfRhDIHavaMpUawNASRNGJ6oWQx6Lruu8UShgZ3fcfedLpYiPFZ5Eaij2yuC
8nLgEmXWxDrm0k34KxocJvGZCLVu4eBbDPDl4i124v5KkqxJVVLY0E/To//iT+zq7ENKtKhCSdjU
xAxGXe1wCGP0eIx7dL4Brj3GT7ei9PfNNDCUfwozHqChb/LuR/8nR83M5VVUHBIVfQUQFwIOvTAT
2WHJgg2xMpfRo5Nli9LmSFIpgwX13U2VnxUHbwqrb0/0+zQAosFqvPvaxChULDb6as0WHnj2Q9Ie
VeGnfWNZLhLvQQtJYqjHPs08nCPxnJxsRH+yQVtc6sdn/A1MmvdSDRf2RiuTrfau3rejlzdD8JVE
qO6GHOs5ys7UjJgpEN5BhX6Bb6G1f+/Cu4JDDBlqQnlN9skn5F2G1Tu2ySHtlo6oK0hlSTsWue9K
rTbwTafPuirlSsVUtY6On3Q4Xc+8x4+g300b0TiIohE0ymTHVsfGN1+E/kZsxJ2W2q1/QYJSwr+N
ivjZTpV1sSL5Q4yfs4aSHmTJgSOYBgQ7UGc3ynXNCsivECtRuNZehzPJi71VQmETV3G+vKGsU2eY
v8+B3lOiUEHTi8mFX+e48wuSstmfElK0Mhbz00SJIl9OP7R44KMUsyuqOMDyj4gwo9HAP6bLWTNA
DTKmYZv2isLsuWMpETsb5NKG5E49t6fSum+ovpIA4BaIbIBOpZ9589wgl6bcYzUBKIqJhHmTrNJB
b6ku3shJVWpq+wVxFt5NT05J6uJlsxbRALlSGYz3OjBwzMZG92qCyNIPxPs0Ohqhg9nm9/AHB27B
Er7zTDRo6Sp/c3KnF8ricEBW/OvI9l1jyMtu7kOQbN+QQRl+jACrIx9coS+0kRufWxMDaTqrCjtO
0TVeQZzrdPzUlJYDZPLXLF7xsq9iDug/2yVbKGWPqR2YNYrmNE2pTSsbD7SfjV4bcKeY+1lDTObL
cTak765vtHJpwHojG4kloUkQanEkIRr60FWhODZYKKF/cr2GmHHW8nJ0DzJDaaZPQY4wTJRBU464
CfEUIjCnjwG8FrfoFF13FWHf5Jd+5QU2PHmhr0WH2e6s7jSfjpnhy3/nwLr5PzJ6NLnpDMoWjMTf
KXqo6p2bp2GbHMSJXQKQmPAUsIakAknuLWrElcdN2EwRopdRR73ZALwmjTxLL2AyI+NkI4wWKONS
5VvecXOvnloIkUByrDZXl4F+sG3FF6oKUYzjqPKzLGDA0B8IyOVxpUvX1JQtdDI+ZLUURZS8UoRv
9mqEdCF8h0mLhFN0oG5fFSOsGQ+GR8aVLdaisA9EBtON2fI0q2bg1CuZyfP4Avh02/GPKbQ7AY6f
n6W2KR+P3ZnSkErLyKMaAzNCW1sesw7vq7Si+HPBnlM0F5/V1uFXmAlo21WNfK8vDLC7aF0Jbpun
0yM9rT4zzc+qx+EXHJdHmk1unjomc+LT+ZktB7BjteWflYncODQ28nd6yj5pbPqBYkW1iYI1RhfM
3MVo9fXg4B2Z6Av+uqeD2t0Hn8MxUG0Vpg1DryJ0PdU7dENk7jy+S2dAUBIo81l4YOxwl6jNMnJu
HTZm+rzLLtF/y37B1qWNKIb1Q0Ow+3eWULzYybpHzxdr06X3hB++uh6tk45DenppecXezmVQRCaO
iCRfbL+Plwbp6mQOeR0uF/GoAGBmVj7DrFhllo/9ZK3iczIxOtYMgRpRQ64MwtQSF76tt+c9TkSO
UrM0Zq9u+L+Q4wyKMBL9xBpVilas/FdzV7cBPGKrxtGZtqrxBSbK/xlybDtPzU2JDqtdMAqw6hO/
jVvs4JpXYwhX5B4qjOESAnvhi7OjpvhNGG94F4Qc249RkheyJlCEp0jPkxSC+cixcXKJFmcWKEJI
YgsBsR1iwLS2/hiv2D75o64fhA8EmErzmoWWKLhCD+ZmO9sbujJRuoiHDHBjjIlzbWPXfXyj1qX7
vkzxgka3+U/R4b1sFJ9WFD2zgD//6G9To3Ccm2TanwKUZRIrMswJsGkZcoOnodN6NAhMCb+GAZgs
JH9gF9qaDyVQfEE8pGjMkcF32/wmOiWqRibsPXjw+olP9N8f4ecGV3IdlGGdipG1h8oa9bvcMp8E
3wkhd+NiyunC09NEXO8ZdK3zu9nfTCWY9iPgQFybavZY5LopLLdrOKXa6IEX8fVEFmRgx7WQfjK6
CqWE07qXq1Io8ZGfpf+Av2X28vqZ2xh5TFkw/wDWu07vfQQEdCR2uXjicsVtOTrU3d+UZctzwzyQ
2KAYSpB1mTSe1YYaOuTKdWGSgAKNdzS5S0Cvdd7g50bxQc1OItNgHpNWDun/i0FFvnDNPfITGwpA
WQv1yO4oykY6OrszAmLsb7WApe/krEqp4TkmHIcBIDHb5mBJ6IJyaMdDPVscem9LY216W9tq2F6v
AixPGxL3uF81m8lV9T9KbGINJw6bmwgJNOWEKsBydlWwuVQeqZ24M9xRfquS/+MJY68Ft5F5TZZa
kSIO/DguQH96ssUNvUxN9+c39DDw8ZQK13T/fuzRZyVHLCcJO9reJSmHXg8s7cYksiNxEwtBSfGF
I5FxTOcAlBpsYDDid49FF0mhJ9xVffd4pe+9E8ua8N/V6JpabI/aYoep8hXqp99O4KxWOTG6KJdK
/cHsykOftiIQuBFGbsF4I+2mwwRToROzfI2Qe1qBN7USyAnmki1z5G9gQf//bK1LLsAAIKbCAnHM
Ac1rDvhoc1LRgJ+wpK0mRRtJykG/ZDg/BJOf7FGV8KnmqQTytf8j0G3y5NomBKbxcokrAeJ67d0r
0EJsJVtExVchgiinQARpvWoa0ePcRBi3cckaRf/W9ZZrI2/nGL3Aj/jVSuIlg0ffP1HUoNfOywnC
yD1/4N0NDzrbYm5Ao0j6SwJ+VDJDH2vROkiHHMD6AsXD83j47a6RpreeJzPqbb4KqjsKthInXnDS
K0nYZ1paRWHNUgBNeobb1t10hZVQBKu0TOd4ybbj5ooWW7f/kbQUUm1HHr899cD0MiiXMme7yDqm
3pfTu2mePJhgqk4RTWPFxbesSThTc1CHO/vX0wmdyjqLkpUBK6hWirwtiL4jPuAWVNFyCyBc6rjR
jhvfvhL8NxIt9aRdNr45kn6uKFa+Uc0Tig2XFfQCjuaDerv5pWo6u42lhbzE+InVVepSJuY3IZSO
/XbS+Bro8HsIZs+8lCEwFGnQdRM1Myv+h+A1Duc5BOautL1x7acOpTrPUAeg3U1wfaMnBiwC7DAg
bcD5qRsboA/o+HusNXI2hc+QuSQ6OHwf8TZoYaAdYtm4eHIULBjX0HeF3PPQ53ncA+JA4sNfRKu+
xnPtzxegrVvy+GDnqmhAg2rydkGarH8RPMJIdHxaPGCHqsYnapKQMsYVhFgXglxizquBeNHog2wx
1N5EsNsCKwd5Tf+NSOhHPAI972sLwDz7mkMC/oLQ54D8afCHfNiC1V/2uanpWejG49yeuh0S71Q3
Y2qX4poiWmVaduN6AWx7xoh6pHM+5rPqpMGf45l6jW+MHzeLaxMNoVt9PoWOHCOZtHEvV27viOVR
bJGShXfUVlgSS7qin8I9mCIqLGWZWA/pfLaBdVvULElixXrQq0QUbUAtWMJfymP7ZZ3RNT6FAdvw
+SkEMdOxqyDbHR9K1ewMuSMjSMx2S2vT4PXm1ECThktD3JCK3GG47SjhrumrFWQEEljiydzwBRv/
8SotPZoftavBBVwy6PsefyWlQg74oef9kJJK9OlOsQLOmh+andobuqHLKQ3skFrt5z5Oc/kyuDHh
d6nj4On+HWUkD34LechNKsTK2iVn+iDIl5oGR/1vgdpXEzCBEdB1bwJzrXaOKEI3osEHFgm0dzNL
veYb++r2kLT6LdYol02f0UtjakEhhOHv7Slh9tm7FYSkPLKPqXgAchMVjUGQrZKgRKwzHmyLNrBJ
qIOUYltkpf0/9hSH+MqBQe8lCmKJL/lV/LtxAmtMCfXdpqiFgAXss0v+In8apGHpl9t2UliSGCHv
EYlw+g//vl9vjsHthO+4IIKNjaKo8XlqzH8EHDRfIcKUM9MoeCSXYUvPiFwvIFxTUJgFckgIgYjd
nE724y+RB/NzbC4oFq7p+HI9EhmYXWgfMpyFpghvfaqUsL0+UA1HK0KQG7Pqgy6urAITFGCS1tcD
OJuwlTJs9sqvlp8p3Gyo8Y7t5tFhPW7lslRs33oHt75k1d8ZCJcvf+YKjypnKhiznG/H3a6Xit46
+OwtTerVIAqzUpvKUrZAhlfCyCi222Mwl0cGegK9NDXb7CjIjg6bxX+dhAosTfuMmPwTr+qlL6Up
xBpWl/g1x4CMCgQ7hmFUr6Lc9x/6vrz9yl74mvCTEUy/QFQ5Pl4LTWh5rtZ65THZVFb1RDJ3B1H3
3WluUQElNR8ZJJm/2rYZJxZJEXslo4i4sFboYeVIjTxDrXiozOKZroOa/4jgHIlJ+uI5ssJFGWyU
XKbqQMYHBuqhfAtVXEgK++oI8zTiCpOZfsY8R0c0zFsAm15ZlwMfaH4jk9QoL3qDaY36gQ62hTGx
6AMzPqAJJy8ZUoLkgBzqHBcsRp77LGTElUzxClbC9xZ6TUBgRFCY6b5CC+Id0KbJZLMbH28ZJShc
/XWe5l+Y/2aqeDJL9oqbqe/WiobakkeyEYCuxpetNl1jJsWgz504En65ZfrcnhA9mYDs64TESpaM
UTuLb0CP8U6+F9mu2H2Etx3lLlCfdZ/0SGv/Gi5PDXg7fB+k8FfeqnPRuLS0MVxQtSOi2KCSjrSs
aXJhW9jYY4fgl6nEYUjWUxFQvGCSN2IBENHYgz8q4DkeixjULMD/0591tyPs1mHVKmh2iyPh25b1
fCWaEy3zxGN7BWQ5iDZOHhwyM0qS1ZWQi7O2VbUqhV6NxmI1gcvT6U05OtTVPJ6vXA63M6CIw6r+
vwFNc0Dy00B/0ND/PYiUv3p3BeG6hyh7qoGbWzIt05gccWsy4OP96uBSpiDiSxoHBHGmrDFbdJzh
s+gnyvKkIXRLr1wNa8B7XpAOCf2w2poDcb7ZvFuK39NEyF65ouskBSRhKcoArV1XiL+Kp7iAVDOk
a0UmIKJSiJvGExOByarojZIcs5LpI/wZE9VfBVcdd2kVYFFLaRJ6mnkkRlN/c53HnOvGMBTLxPWM
wv2y+2lmfpA9TaSsAOKNFhcD5FPvB6ZRNYO/b1pbxE7mD4Wf9sQYS0UMjk3aiH9Vya1tWqb4e5TX
3beJ61PsptDtCax8QD+TU8hmwMecp3C/2Dme6k13Kw/GSZ72YLr0GXmyRIj5415oEp6Nh6k+xHaD
hdilax+Vd+1PRag64ejpDC+l6FL5KbS0OLUS+fJK7YZkAGlgQhbhvtA4ixKiLSztYn1qZ67TGRLj
S0HvoJtzv9vcVUXRgFo5v98aCRz674BmL8lVBMk/9Zl5xVaqQW2rmZJhlhS4Ni1ZAIP9LTLwRCoa
dhwZLV9vkC/GQdeRw/AXEV1+wc+l95s1AQ24Ia8QiP8IsMdDz+SON51PM98EAnGzk26tVEJ7F+FN
vhHwUZPytfmP9A1XSX5fei2XbUCJoBrHz5ByXdz8Z44DnVgdHOboqog2ZSq1WQrih2Dp0u5KqYk4
PDBokiLboaIWgBeBygRaW/be2acHWBN8BI68MkGIQ+3V1IT9WOo/w7as4Erf305P2GuvVw4n6xpH
S0hRJOfdOpAgN1m6XZqbG0AyaiFhsEGBIJKVzRBsLvw9pgOwL01fwJIaIVJfUYPM6lSCiu1NL3wS
/khdupZVOO4wV7kSrb0spVSzSxwsJLBWOOxt9yAGf8mDhoe0VABF+b3DdRZI43GneK0QEdGrUcTu
3yp0zvpO02zZpPEnIbpnDNWhKRKELk9KCBxNXLhsKYB3TuvrpfnctzoopEKenS2KWqeJTMjs/yx8
a9eJhXRv7nDxma7l9JcYlFr3dHz3a2q4nJlJ0gaa1OaZlLL1VgppKHsBiwFEGM3uv635BZZyVq0J
OaV8JRwej3+tky0LuKPFFkHb6umbU0UmLlEDbsLvVZI14ifSxq/gUUsmYSrjAGbFGI8hEXSpSBUd
J0Hx3r/G1kQq7GqvfCntIMfiB2eDjrTFEZVMIvYEfTbLgiFlUb+9HVmKGVlE10l8LGmt29b0DFHQ
nevEDNubDwo9g6knYe2D80bO4Z8aO5cVdBpUvzblFGvo4qxzLDeUXkGg+FGab+ZhKd8kej1GhhvR
xRO/czrn3BTcXnSfN7HZstcU2IVZVpoCeDbvizQuJxaTo8WsmFJgAh4Ac6KCMSLXWXay5PSqmK72
58Na6mi1J3JXUYgamypNUty61reejQ8zfky3SkvvoDP8LzklWg1Yf3yuKeVZxPl4vEiSW1MhA27Z
VDaZEpH+vaHpkj1Vfw/n7tCR59jUUEnx9VB/cI8LmpbsARqVe6i7m8nfnIM4Dg7p814h9b9ORK89
ekiMwOKkPIFENA7Me+hNJnSTL5eFSCmibsj/c81n0ogFHRihdqoFM+enZyM6hGnlUC6sO4VUX1Gx
WGllBIpOT6Vj6qJnJ/qB/Qao3e9wvii2vxrY27FowhgAv34Bd20QUJihyHBQfIpdVzNClTKQ6Can
IQEiWoN66h8g7cUaChnji9FNiS3IzEuFVmOz5h2M4jOconyiz+KNeH083i8rRx9PR4LNgB42jR2G
vaM9XIHa3a/suoz092o60IW6BomLrPMBOvh3lM/cxGk+0aGW4uDGMIe5tRCrK+OBuyttBM5lpG1k
dd89i2XoanwoC76/92+bzUfZkVKLKOt4Kd70zaGhmYzIEcXdqA+BvqmxtIV2EE8CP3+DUT4NPfy0
JaQ/oT4eD7ERZ4iGK21ZcyoXy6BENMlFqWvPJYVCotjwIhnjPzKnAHaOcIb6SGnNAcpkhajtCVEK
PS4NTw64f2A5WVUTKCb6BHvMsV02C1upVm75mh45AxgcLfrNW42pytvWpCDEwWsAhoKEO1XBAjR2
/dXFFRlh8gRSt7QiMp96pXoMtdgHLEEU1TAOPJQYtj9K4NoDMTYs69nf9nQj8qvG4knTWCieSjVE
qhtYjvkZHLQcyMOBlXK4mR/yQwSQA4Pd6Mlk/Zwv5wgauRag4uh9rD4RbGWEJJwyBf3Jq6puTyeC
0r+0oYOvZHqqLWJYIiI+/WfrRkxtT0xF+mEgMIOt/0lh5oabPH7idd7Q4AiltsagjMSorcGTvvJt
sMAz/oo4LpDFeHn02sV7ukaRTq1cdOO90DidZ0hxFfizUDZzpBStT28y0RA/lPeD6wzUxAF78LPr
1kRv5dFV3Wz9sUaXf1JOP5cGCbxULbiNxsSn/6ubbtT6xHXsS0rzvw+4FGpf64jzrpy56kmmu96M
vtTIuPM7VsPCmzSJoV0MPLzvtZc91tz9FmUCVVehXcU1vzsIxnnS8Tbm/pO1Umoy3kblR/hqtIKM
LyawZ0Wihgl+ZF8S/hFhsY8mxXE0ya3buetWtrfKkjFQ6cbzK8CAPd7n2NYtl429vwONsyWeF12d
k4Ax/J7GQV8mycVppwBQxiYPeGkR81/H+yxm6gf4yqpU4Jh+pSLYkA7Z59QxYfSXY86IK9SoBnRN
ORtUXjIGnQKiTXLfPP7v0xFG4//u9zZVfH0kz9yw0kOVQBsmhNa06lSXY6kkzQ9taBeDKx/U/moU
MPmJgoNL8G6FECySH8ZVVZwV3x49O9tA77ok8t0q/bYgzsimKkpa/kXIbN5AGZFoEMQhRttVQKu0
QFYXPkxnyzmG79BscugCP3nxM1VtkLvpmh/uGyPDmlew/b4NfMOQkIsQRVTu0JYo0PhXoZoRJ8gM
xyR40axWzZDi0Gs7/J0YNdCrJUbbcrjaRR18+9YHNrH7YSr+l8udJdBVt/TtoKDZCGWRWmfe5/xM
gLspfcY4Uc2+PR+7iYQVCvjTowoTLKQAuzBpx/1zm5yT2XIp6f2TJMFefwR9jLo0zRfRNxP7XdAJ
efsxHNaxSTtXlF7g5esjnbzaqdZ4R5Vto7ganvRRTV7nA/Y2iOFvR5+XRkfnwdr6uwqGQAGsU9rQ
XjoJ6y9kfuJL6IC9LOd3YRKDrtYepOlNDKpQFaW5W+5mxMQ7Sqmw+X2HEugEQRjGvwffKdDVaeW0
NY7fyOxF6dPw38VNVeGL6+MrEzgY0N8z9KJhQwx+h7CUa+QoDC1ZgYt+bBLURFGNt60aoE6cwnoV
lZugl2q2LVKT+8ozt83Vb2Zxc2WZNb2krsiAterU/5Y4Qwb7Nwbg6USJeDERdAjSiXN2u5jfWyVW
7Ar+eQYkElhVD+fV9srcRIcly7QCs+0RlPZ1rLITzESo9TXav00AySbtYwTDEaD2lDiYqWmX7N0A
yRZVNwADGDoFxfIQivIvSIbrE2CQVEmXrw7ylWlQqXZELhrAbTV8MiamDrLNUK4r7QacYcHTokV7
Qf2pzDsqz4pHCNBP7xQl337rhYC5ahFfH4/M9hQg7ey9DMWV4RWRvdGUpWftHZQPZxkY4k6pM6eY
S+0QWzNd87ccpHC4Q2hv6enTuijK4G8NfOSo+TK2UTjGE9G+cucGj4O25RJgQYJY27flVV5uTXGZ
K46PJYxcUnYGRqIrwSN1QQ1ObMPh8vFwNpRlIYsFIvZsBltXQD5VMSlVFzKlTSMcVGbIxYdOENfx
9cB3L26k/CtwbxAd3xdFNF7zwBbdfwWUzrZxsO3FYrG2FX7VNKcai4TKjbWtZz8LslkIGjyVd2BH
v0L1z3CEiDr1yezV+jWsBjOPZgj0CEKgzKcbNZU3cWULgQfGCdpJSF+q0V/mSJ6nPG+geDKwv4RH
mbnc6MgsrXph6qhO6RQ/EZXe8F6OqpKXglWopDuoxrZtcUPaf2RhtUGpT/2Q+smcIliXzKQMVaC7
sel5+DXVVbHXvLGxYgEG2ot25wVPojItI97XZdavqW2kfeITgsSmbNDeggLcdbeW7834QBPqSzrF
wdx4x2xNGLkwqfz75fFBPuJoj9rZ6gK0sSvdVYYDQqwxe/XRwflC40prZqm6SRWG5F0SkUEAoSeM
kxjsewpxCmkAXdCreaoIM91Wm4qRnBtXB2bqBvqqUFh+CNrwdFRgS/m6EvmYd+xlHSwL3uepWtpQ
DxcNzFp5Abxyx7K6Ut9zSsRV+Du1VoA++g/46EPVB3JRgV5MCqctDHuh8w/+kDrJjyzLMFa7E/mc
l1pic3qctH1Ix6eIXYr3yrcOes2V9qDEqZg4sRKPWJfoznBMtKElwJW988djufMMXe3WL38Xsgg0
Qfnnb/txnwo50gPtfg/WYIbjz4yTdFMUwsLjAItOUiSrfUO68Zrd1VmZ30g8G/ZGEb3qMoo6LRWu
jHeaElXxB9XNnnsKVSFnvVw463HH9hEqssJpfDB+sxbdhddj7wjhylpZUgSLBPsjJraXFeK3KRNb
jiSE73ditM++s/LR/kSP609US8nzLtJbS3XjSd4G00sGwkyrqsb+v/ToF+yrgacl/38my1AvfpmW
GALym1nUnLPHIx+TH8MTg4zQzVrJKC/Mtm6nv79y6T2YREh0GvomW/u+udl9Wj0wWL0eBbqqWRM0
Yvq8MHDEvCiSOa1tHRs0kdoJQAgdJvHEyRs11rtw5FdVazq4YOsjsNikbZaUvVQkwh+MGfDeFmXL
IlgAdpy9I9x6ill6CF2dgA3L3jZdhNt/gON14YtScdvcsiFKxmdKQzF9eg5eFM8z3Xm02foqkgng
mKDpoKrobWsxFpTrpCiq3wxSqSEYbi+x4TehW1Je3DX9Yk3IqCl8r4FMIZ5HO32t6BB6X8dSeXYF
/jFuc0qtYoyIhbxIl2hPJGasmMHBHfrYB0Mmi5b++eKdPd3X1QgWhHd2lqBTU96D3WrDKsQajf0n
jAQuMk/IqgDLusU1J4+G5hig6+4gpN28OUK+aX//dXqIzoKOyaI4ooLihm0QecJOI1FgRk3Hj8vw
rKY7ugluOWeOmda8ZJd7hNn3RbGsrFUlWrp2ynDOQM3dOtIbwqKG1kSwriIJGVPXo7lge/4wZTFk
SgnYXAQu0MJAiHGuLr9MkV4mgO38yxA1ObH/WUcd/Mi6ihnSlD84eZHj5p7QcLt91R3kgH8COmfK
3KxZmTKiqEB/Cb9gU3N8LPA2sa4tx0RIHHOZvsfUBbPWSwk1G0hi9JG3UFZv2c2Pjug5KbpVUwiE
G14bSWpkSTAxw9vmhTknP1x1yLMqdm1OP6VkRafVaCu8BI+MyPBcE1pWjSPVCDuHOp3fVw+xv6st
x2tkx/Q9nwg6XkxkYZC68XBiritrnk6tq9KEG44g6kqMdtgwNYkPRMupYgUGhSHzonPJMYKcZuxy
NVgMvlAN/ta0WHG7HvgPPkn8CFdVRrnt+Jy3hKUADV354JrB2CXyDlbjMKSncKqK3dErooSD8I8n
HUZejSMan/U97Q/pA9x0tNz85JAaLPnGVpt7nnRTaoSwCcm+xiieHCy8UuXwAbC0pYYBk4Vuc27n
TspCGQuP/QyuLJkxCG118omOskfQ/SpqAJ/ZwXMKCw6sHNjHE+duzDMzob3jl9zQM16Nc8Qc2OEF
PLsAjCejLtERqcmv2t5d7ff58zpDDfrJcXMEv8NamV0REDqJsti4KvJnM29GowURTp4Fi3XbPTQa
KriSqDfKvTilvMOHv6udzqon5SnOgLKXP6GSRfIv54GRfCrvhX79lhw7q+B55/jpYfsikLL576ay
aD2GTUYuGwBaFtIio56OlZB6mn5mEijO9sEsos6+Vlsumu24hINrOm8ZgwM4s/pkIvZXlh8hsxbR
ExwKiMG1iISTlrrtCKzRZXHkeQyGj1IW7ap43W6lhejBsFm0H3itcIbI8gSYcCsYRSd8uebYrdeR
/V6qNrnuqOJ+6tlOWRmtGfsYSNUQZTh1MXOq941s7KGmFg1LGVeC9SgBAYj2BblzODUr38zTGOf9
DS24bQOYeG5PSe7vTIGFjjJLNMicCKc1fcO/Zq/xF+bknqu1I/vCfkIQnD6nMGzSnVmvUToiyPMF
gkBYjwlC3zuHMEOBhJfc+W+oLElxPiwJwOME55BaIWuxlbt9Iqsm6gjveNpA2WZCNkZU++K/iLUM
YwZM02YKN8k7ODBQ2ik5+5kaxvB0A9B3CywS06CLYkXqB/G6R/wrJOj4LbR8TSbMALnXR20tB5y0
u/3XfFCGdVQyTfjZaTUIREf8Fq1GMy5DeXJz+L95Y/52pWMd/SWt83IHHdoVQmJDtHPvWdillewf
3waK90EQZjPQtukeC319QL0TtjqLV5ywmcmtVyDoPhXHizRe9VOi7l8ApK1PgqOXqjhHbsj9fvgT
fgwkiSHSJ2zCRLTGkuvUWiaSOQrFmTZ1fhE4ghJNY3B6qs2PpjdhCjEUz15qT1KwApVcdVoumBjX
ThonCjp/q2RMiBgRs4K6OSXyc96d3EMABuaujlIy5mRDpmdfrYPFrsQiUeRIlbm68OW0DS4bq8KW
0zi1e/+zLJ8qbMBS883wAn39JeDPFzgrcgqRYK6esv/8pW29p22zdNAJMEVujtknXjxtAIAI2R5E
KbBwPZGBa/eWUXMQjhivILehiLQ8U7xtvXUVFaRJVsSM8TyBJ61eVOv8NuZfjvfakqiZvSEoAuNl
QfXhSVsfdIu1p5hg3HljdKqgEm4/djynAGYYo1IHsFBAH1I9y0dAkFmiXyi/P0SbWFhN8EOVbtbs
NDyoZZ/Fp+Cd0962GjzYLHVH6e3hMmcaVY9W161kNBKZK0E7Kbx1nz/YKyi/Z95ZQ6p4Yb+MK3lf
1ZewAWeP1H1cBNJj+ecDU3IOi3v7rbFW170XwapmKlUHDvKq2yCLfTFq1qqFdHIIkE/oBcOvj5Bw
kVlTEO8ghCqVEM51H6b1qkkhsmaj2ewf4WTPl5bQnmEZw//6CdzeAuUqRKe+WUjWyTzRFf3bGjK2
hPeWhlVvtvQ5RhEuDGaUk9WqQ5KaKbN6ngk/62fizdsUqFN51jxQnGyt1VkIGH+LkVBK3DiEzfNt
qHGvkIZPqpfHNa33JdfqVMqkgwEdhTBA1DG47AglCsFS4fuXGXmBZy6q8knRWJl8Q/Rz0w3p3Vpa
XtTHsf1DCMO2Iu18oqIVp9ev1tx2kUvsjTo5ePo85gdxfaBjnGqY7h6pzcX4Da47sVRJm6tF2Qj/
sDzVzCKmtnsiKBN7eBNdst8K0vDfMHTccfTSkWbzbamZ6YIZvaShXd/FVMqYMN4gLFeLsbx0Ob6F
R3XTB56yK0jbq2d1PvmxQmRuP0GYT4NJBdEL6lOsjATfEMEin7b8Dv6pnHYsMncQW8YPtqjL3ARX
oyqlVCG0zrtl2KBu23B08b08R+9NHILZfV+WbqrAd3K7rHGDxEN7ddwEi39Q+dt3xBVMcedSPGjm
GkgFtkMIMv/OtHangA2xEU5pkW5veIHZG1PadtzdcATtwE33nnkvc7s1MJhfUKDaGYLPJwZStmYW
RnQJCl9RfylwojPgA0UwYyAMLZq6ovuPL3ncQmFSsvaSZ8bLeEAOCE6tvxMF1y7dN+sj2lAzDvm5
ZTCxNL6ZB7J30bVKctHEjteXJMwN9cJYzZU7LypRnGwESFHrxv2LjiXG7YV261wffYTJJH73IhnO
rCSb1plH9bvfoePAkh7z9exrQSfRqzkJ6kEHZRkyguhy7aqaKYSCwGYJ151s0YZSUIwpaasJ3aUB
nFPDvVfipH8JNF/PNRS7HpobSN2rmYKrbAhgZOv7Gky/03UKRtM1P10Yori7QGJQjK6Ir5FR/lYc
0a94SrnrB5iO5MoA5mXOvEPupVK+kTwhlsB5nbkur686emRs23vJOaM0dRoRxPH9Vf/W2Wkk1Uo1
/BV2vKxXtjWAncsNVDVzeWdls7CvnKLqTxBcCdrK5vew+ytQCrFZpxVsL3tp6r6bz+SNlbFGpPpw
pc3EdjzLvM82lAwZhRGb/cvgdxPPWOf7SrdpufKeAllWw10txQTUoxNO2N2ky9nw68w1FjGVxD69
k8JcRvA5QTG7teBEZw4miyeqqJNHNc5UNUDnUExIhoAq2aiEFXe06TrgVI1QRD55QoHGZwGNDX/Y
m7D2uUS1y1EmOjtC/zYY86n5geGrviOBPzindS5eZaM0uS+DYfKT7FYv7Fp3gPZWb1aZUZUkfk6/
wOYybvAn1G7NxtiwbDM0TQ5qBVxmB/CJsFwjetamE9t/ZMp7BFSNFLckJUm/1QmSuy0Dcv/lZ7Cm
ifGi5Whm9l/kF55U3U0pmMU+lieU88xEWqPpHzlbafS+xIjWtnT0DsR8dM5A8MSVazxa5ceiBwnE
TkMv1++uBQTHTVlDkivn2o5ev/9QKzyoP1jy3lATEWGps79isGDPDyK29gypuE6NvQ5c4Rn9gSw+
mdO/b0wnA9GPX/dRMbCgmcD0OABgUuRIhmev4g4Qz5PnoEy6MUd3qhJkfT26CTxoX/q+Rc0wwNXn
iW8lANFAZrMTqCij3iVaHKxh3Fs8Fbl2Z3GfLEd+Nh7PIsEkuu32RFsLROHANT9604iD5+qEmp+7
K15R48nU3ngCsAdX5rSDcW3Nnd8kYSr9pNzToQ42v8wnLIkhG7VXhwsItTqkksvIFq8ero7obJJa
aRa5Y/DCFXFofsHt1FBCMDfzPdWFoAW+VaOQ8L3QGRrKm2MNyNqQcxPE4EMYnI4JEozimjU1kwL6
M/032DLPMQfSlHqDPdxSCJRYt/paS33uOUpjycTTNcgMPTPHZfLPk+rHvuApO6I/y+ohh3ujWHZX
ujKW7142rmBm6tGYu0dfZzGClB4P2yy1zn1SQH13Cl3zmLQjbyN80Z/8tkA28u404zbOOoCoN3kh
5LFEJfw7DrM5EAaf+85V/3TANMtVk3+NVnya9feI55/FbdUBpZL1t6ysMKRqkGPbL0aK1GAv5ctp
TtI7oedIJVWlwYvmVMYqriCI4kFo+DoTU8FjCyllwe2iVM1wvm3rXaPdpFx9uqJ2Dhe+mGrlsI/9
dkvnVlHAvmkPK8jW5gGmbgM5QDBjaUno41POgm1pv6DCBe2rm2OWvWQyDCRtjgiLuVgeWCI/1Ve4
B0MKmuBysBE512wyRg0bKUUxeuPFzVSchvG39Z1HnazY2PhritgFWcPUpybwZvyf67ZqcWo4atsW
V9VadauLxzC0pt8++PapJKYcku0Zuds9HmoFjldthX8afhtbicjp53bgNXBvdSj9sq0sk9HXc4LQ
reyRoKP/azQrizfpIUtKE0OgkaoxGBclriLTqdqDBi6KJ1rAP7Bej/YGlBh9bSGEjIRzqJxvXqtE
cOr48YymM6PS1G6QwRr+d1kSUPX3HAgRi4cHsga0G6IPyNeczRG3xMKuS7LRtScS1FaI1nc7cFMz
WuMDd39Up54B/gpJ3rbU7DArTIBE92/EpIj17SSt2Heof+63I69aue4ETO+HLrdterSP8n2xmuWy
8UoTsSYMq1MkIQOheNOZIwY3A5mbMCi9N8N6WycbswgFDy7VhjR3YlgqWKd4AQuiGhvCzTiQvTbG
MXteFaBM38l6AekHIU7HSTZzFLO5/DF3uTY/04OKOEvTJRxHNYEJlNkRuBIBbfMm2mbvjtJ7dgyJ
R+aHDGnGZFaitUAo6wmmQg6St9WeushKOI+qVU2eupMwprip/QZoDFjoYsRsy8J/eGyl2oK9vLUv
R7hTwaga3inei8T29/hgebVzdxErK2IlT8y+hjkvKTdxws3VK9SQ+o/qSszdPlUGP/Nalm/I46Yn
PPdVdTPWeyKsgJaJNnY560majGkfUUH5TLSp2L3dyy6d7VQUzZxKLDVKFOA4AHUdYqUPOKmVdx4d
2DK/XNxWfNNpYuguFgzgOB5wseUvC2PYOxvBpbYHEpNvdIPDrqqar7JADzTKxt2sOQempqdc+SJF
XpaCBP+BscOcyrYxJ6bjZw0ZAIlPxVGlRj8MYFdDJ8qpKe7Sz1/ZPpTYa11SbXS6TKkXepBNJgXm
a13mgquPWxv3HHtt8SDxofl7mP5mrAQIpTIznXBMfjOK22ka6qA+15hBr4bBho5LYYYz2Gyckm3s
t1dKAO6cTeMBNzOxnEgRPCbc5FcIYbhbL59Ptf4rFRSfTlmJJihV/RXdsT4zKUBDobbvNIiKs/1e
xaxjZBLwoeeqoOVYAnuVTP+q2eAPDbaWu5srZmd0gN19CIXy10D24AdzJYMXwIPI4rnxg31Pca0J
zIMVA8LBHiWuJSoBgReTYBIDKXNTQnqPjuJymDjQt48l3pP1llf9Ca6gJ7mK6Q0SaehKPYuzBLvH
5jJ6JyyInNmXW5naq9iQ05coZhWu8e/ZlnRly4qxiOU1QWkHoSn2MhmlmSWb3h9+RF10VS5wUPW9
+0M20vCeSnCzc85gz/KSSTo6vqLpUsYAdo8X1apUxdfBUtfmygBIFIdv1NsJMR0UOztlkK1GNYNA
tdY4DCwLL5zwK4nFsbqIBc3Pv90h4A/LN9C8DbHhiFTuPhPhYpotd+DNHWR2FRKV6tyJXqYWrkYr
01POLeLNwTLNogH6QxdHZWig0l+pSwXXN7g5tGTgz142bS2G4bdTa2qFmuFPTyiXHPDpvBln43pO
tQAoCOiC1d5CX//nQWItLodHM5YfiAMi0QhHcOMBBwPoylrAdxUKi9WFfXLg9uyBOA7MYXJK+KEy
KpOI041dBnI+Zd8n2BAB0VW3O4dN8spAZsH3eRc1DGXtpuUt12cQ/pTyLIJp1X0pODX10rI1wFIm
ZjCf7mf/ZXJ4Hve3yVm9AGmayK4aUJUE8ftqkdg9mALRn0xHsePPUjMM3mfn8yABzo97mLOyiTT8
mjO9yL2dZbnMB2/GvkcfTZueOlt3RJYgVBhCRxTIaHAuBxELVADu6aGoIHiq5gu2kSh3CkZH9H0q
nWM80wWquBcOu2kOMq5ExJTSoXj21DJZ3teWiubgmlfUMbE7JbnWwgAZqEOdfe82GPfRxarWJfhl
MOkIa9J+bcPm/qxuio4XwKmHu+u3oFvJPVqv7LNrY92nb3JJQxCd70CnuJoncgdl9tOcgGn1Q5SO
RR+yHNvgmyilcm16PKgU7lwm8XitMSeSyKSEtDWK7xCuuPKvO3D6EGy2wq35It6nT5KO3vSeaojA
jO6DQOpfG//iIi7A9lU1ZTwyNoPwT/APkq7ELA1I//qNKv3FdVKg7Y9i3Qk0trucyHdNQjzL71Xx
T57P1ZLrF3lEcnbMr0FZqTMUX8vTNSgqJPgzD03GHA6F9cIWEt0JdAJC2ywGScMcdOLxu7AvY5vp
BvJoaEy0owvNyB1N/EwK6ElJGCietiPUfjQZ8buWlvtse69LmYgFKK7i/8azsck3Q8CEjMosQZpk
FRTiKKPylaPvLJy3HjV+t/S1goKQ4Bx7mwfz33LDthPZB24WP2ap7LrmKNlg5WFLQ6Wr0gXpnpbi
pg+goRehz2C5tPKZPJ4zEut6zIORZI+IGMEgIybj0H1qRdiLos2yk4LTBo7JIsdW+Gw7YmUmqacV
+pBdHfyIyIvBRy3DwRYXIdo4BopyzcAJEyKbw5AXmfosn14gQdxexPTa46yXNgw2JCROjYenlYdB
yOFq/Pq5mlJQxv8J/v93cA+EhtVjgRLmLYi2naMEQJNdsK+2M+3nrzTZO5XJFq49KAR/nhn96ttY
9uTBR1xP7p6k6ai0a5pj2o3gElWnV17D6rB4rUxtcewbpcrxGxl0ZvMsV/AwqeXVChvz1EFa4xfN
inM1WpjqmvOdtfRgd8Q+orY0umoLUMyDQdg/SItunFrxOKvp3WW7pbfJaZOVjM9kaZ5vMmYh6ynZ
6NHqLn2FsvJb+uVxDhIBj24RBIow5tStO52muqQPxhYhbXQDGer6/4ZfVj+hfFzwk8gPY72EQyOX
zVbSwrdzPTjHS65h3xtsz6TLRrfR9RVAzraH5MbgUs16Wee4zJ8CnwTj3dZlWxjrhHkk5aFOzNjD
lCFfA0SnwUiWjTN98QM2aDxKMuP104uM1UjKgpTB11JbPpNktrll7VAaSANX+UVhE+qeGToqP48h
V3s/enxZC2vlPuBOWXffZNDhbxSnhuE/jDRlx6/me0/t+Lj9SQWAt3LYZE1c8ewijZifeXSSM7P1
e8E9ig8r4pSFDtKdyWzFUzOKlmrADzZCKi1LQIbeU8p4tHgI9MmITtl5dWAUtqnND7O90DUxajuf
XGBMGARasbRjlnl79RzJFaq/Yf+gAyGucqzaV28RCFtNCa3Ys4OLRsPv8F+W2NUXQQRdl0Er0IhO
zT6a/CyeewpirdykTFVdunnrm3U0U7Et/h8XMLhUg2sdLFm+K/ItXinq6e+r2buOFq+9qyIBpFlQ
MzfulIh9Ng8ofjZNIZQQ5zMAoZmQ5CyZSW709TqutaXfWC28uLABehnSSbwdMtc79cIlCphu6bcd
C6klUo+1WTYlJ7F+gPe+BozRJ9iJuRQUnDUMaaKFj+EeAfidoQctDObNIKMG8x1/iFUJKOoe4alO
8XQiYrLtDz6+ZLG/kcGHRFicEmEOM/QG14zWfudW4sDnujMyiPrcMotkJDodxK9fbJjdnZRfiHLR
7nSJbyDh6CiNk8yCT77K3xwpjIy6YOK6vZhWrpyh7Ft0q5O7VfuUqJHCtwFXUw40yGeyOATTXcky
ZPHwO5iUfVB3465BM9hFzt9KkrUqh6aCRDZJ68Ffd9b4Qcx2KbCdxDJQUps/5k/6gMOPzS8pvsx+
rrxCiIF3KaZPk4KYFHOXmNh2QZ75k7cUqdh4nkvN4o6XqipcETT6jIc6IovckOHZGzj4IdyqwwdC
2pk7qvmeH2tgiZtr2JQrCjdXlAGrGYkbbsLJ3k5naEzeUCS09GklbcLbdZ7B0mcUlQibzfeysbws
chuk3WSzeNV/eF7FV5ZQ1/TE9k3kurEs0WZhKNV3aJDZy8RQCJge2d4WjMgbfKkhenfN2RqTWuxN
JvtDsZz4owSrzI/IsCRBhK+CnNOMzAoDg/JpicujtF+gx7k43Ii+U5E+mI/ft3Y2GKLjBhCRLdmX
zK9Emnee8O5rEsbf2jzBr0yL9A0wQ25YVOMgraAVxRqqaspN9p3zEOf9vRZ4YZ+R6+BzGcO4ZMbx
haj4ceubgMGSXThObCib9CPhEi+tgxFVJXzXHE/xwWlpUypACnCi+tyWWnMc81m+0L23V4Yy2sqD
Ck83Zn2y/cjsrRo2OD07GHP/4pmfHmRB43qTK0cHIgb4DiDI0GU3RVOZuW63GiFNZC1f/n6fGBsi
UWYWRXb17J3AKIvLjUx1ScA7g+P2dSJG+0vDqc5ebelW031+A14XTQZbU8Pg8vJHn15s9u+KUsca
5Sax4vk6crDVZwj9PeicS5zpD7dcDFok9I0eAJnRx7N46WT8bKaN7eEIGQV9U21J0vc+NZ22+vcb
bP4zIxeJayhmnRqw35Thixi7thXVPK4Q3pSeaFYy0JhrqsUYWiKu7xZtVdOrTGVAxcPpinHJB+t7
lZtu1PlzlDO1qSsq5JvuV5Yl5Ecllr4LfJcg5zEpeOqksJuTedJHm9SrfkIgqJWhbIcslW0f9aoO
cWmAE+VuTGDZMSaTYW4TuTRQLWv8hM3wupLCWnW9XnIc1quEEzD/K1yR66r8nWxk1dzNtG4uzyTS
6s4xgkDUg9+K0s3VK01gj+5+Re0L2L56+QJAxIMqxVRGU8J3ienp/ls63+r4GS0+XXp8dJ6qpDJE
siPhkF4XOO9HgB/+8q1je399HI8+0ZnBt98ZK5mRLg6ofK73J8jCI2Y0IQWT9cdsMTS7js9JnRP8
z7bRHh+cyTC+NOYnJ5TuvkZCh87SWKf7JnM/xivHUEotcz7Rrd2gbJyco7f8JBTmWqbHSP6rs2h6
KksrL8hFIsZfJ4OJps9n4TmxRit/jvhQAcmBpfKsz3nyTgoirjh25C9Lk01xiWRramiT58FjvbGE
pU3TQ7xohrcyIgMZ8JMCoEcTD/yr+8Xp9fZ77ES/81TpMiXlhRggVmzsutWqJNzX9PAGLUzmySGI
iBIQk+dAlMDmQ6ZB3mIUL9CxvjmFAogJ29JbQl+lP/+DAilbqfsdwO1NXAUzWMcx6eQH6aFFZ2sU
bXhrCUfAGqdcFEDFZ8XSYLdX0rB9hi9971Q3SybxmjX76VjGsPX2pJsIEwxCT4mar0cFgKYbmKMV
z5rPBF71GgX6A4VMb9p8A6ZRNGcRELr8/fgMJPUYYS5BONXSWE6L+KutLCRFcVNLygUN4DVDiv9Q
JLK5S5Uiu2ExwnZUP4MQptH4U9L0593vuC3j9Bk/Nh7pT/46ZyP55OJWPl2rvOSYHw76tokHnHXD
vHxxAw7jYCqH3QikTFrjs16WA8y1/7SZkEjZU32zzndBvepxboz6g6dGUXbXDC1JYvlTNvdxCnP1
xNy9QeKA/szXSXjno6EScK+xM6JYzJlgUEkhxgR1HKoKi0Rjq0GPLs+Umns8FJRW9W+80wHomy+e
WzfhfW9wfA43JSAHCDXLqmNWz3RJvrzTxO5v4PNYhS6bksef6eu7lMSb00jBzC5ym/9Bz6Ky2Slx
Jka/1ISobIRIi+t1rt42vUVVZqbLK/zeHvQJonIbdYq2E9miSnr6uSlajFs6LOND37li14u7yLiE
8/XNJOO5JnTwSXnw5Px9j6wSIoI/0mQndW6EVOx+kaqhS8uhD4pnCfrN9F75nicJwczU02RHds2a
bGD+IdmUOfrBAIkNNVX4a+dE+YW0GiJdfQbIH63nKYXuaRW70/g1ovbIaAIadwDZic//I/1F9YHK
y5/TVP9clBn+aC/Kj3nCv999yI1yQxXm1/D2ugJ1dsnJaEeBr9UhP+HzV3wnmbJ8s5/mq3WJsoA4
vASK/z717GkXvvLh+GRAXaaytVzCcW/+/YkA7yF7zcR69UoFTdpPDzk4x58B9qjIXRAvMLLHcqzk
7eWIQGBXw3ZXqO9tFL4AtVURSXOOpa1JKVdPgDeKI6PyOVQm5hf7mbe+YKT57WoDJk3IKktNDWd1
/XNJbeZ+HNSTFTvyiV04h45pK+WgQ5VVDUBaZQVhtSXTnlwhgVYpFjior7OLAFL/JB422nW/Yjvk
S1cz9SLVwl4bf/VXiZeH/5VqRQNjrlvDi0N2rO7K9cQQZAszBdqo9Jo149jafbtlmBvSQOgWsr8e
s8vknynC1srli9V56f3TijJyf9VcaSRRQwhsmfxGW+h//ONo7PrqOdTk6F9jD3Cwa3k6SXxxPxfA
qI5beog5MlVG7Vc+J1BA+8j1qNLXQpdtY/UdjvLUrOxi3tGiHz9rBpFJJJpif/GAmDx88vorFgjv
18/i06xrlqI+f89nDK1yg1+AXA2g2F9mOiPIHczlSjohmcP4oQ7oT/sSOzoEDtoKgyLS2NgfTjkd
NrAoVU7ZtmpP9J0wp4umH6nFQg70G3RVQuJws/9/y42u+BIPL8VA9NxXF7H8ZdTLu2CZoMy7FeE3
So6Bpr27Ui+aDO7efnaAOSxTi5d+m/EHBeVcX6V/ytk7tg11d4CSzNrmK1dqWWjEUIg0dTGQRe54
rZLrvUbmctMD++llCCzRDijs1P8+clbHfveId9Q/qwS8P3aj1r6K03p7NeI2PmJ6XFt2Dqp4ZI7q
D3OXNOiV2ofwZb4rg7ltzRdc4gMhIYW8LU/QFaTcMXgbqVxvGMMZQPwnRgfRx2m/Vn0QzRt7g5Yf
8wxShvFNO/f41YHNurHGBDKnf197og75yt4L76IwRYQnJBgv9Jg9yMJ3WWYgBvlhqKjYsXWnjldv
mCJt66u77klVQH6ql40m9Q7rgOkx+6pLAwgoD+qe85MLO+2wijknM5dADnCLPvc0R+nZjyB9Pf/c
399F9qcjlgV7zZk+oLS/XAz3X+YpDjvJfY/zfe+Ab/XAX2ixL7ppkGGvkIHD5PD5zhYySuFe9AW0
zrx6ldq9ml7LGNrNS3fJbnlfSe+AL/xgaAEPHgfuKmRy8CXkmkHuPojAqdP/TPH3CvO8XGH5AjrB
gcCjVZXCCVmDQTs5vDuWt+oH0RnsYDIXmSXzKcbUakKqkJWjhE8wSHjFTzncU5pxdZ7sMwyeVfvF
c9Caijv5/kvR7pP147tc0A32VkAlTw13aKQB+GBRcvIOrC0Hv3aOfpCHzSnhQJ5uZxpJoPipmmoE
4xHPu1jSqi1vEgCfcVbAknv4GSM/yvED2/wIWaDTylpVqzSxW2I2oPLVrLN133Yru7frBqRfP7gB
hr2ztVPwkdbqyxPSRTAj4H03RiaCNnGGvy71crzHL9YMuC0g+4OSnO+cg9zHX3737KGq0ymW3N+R
zlr9bbgu5VbtpTPbNNrs2o/FpEkw2fB/+ey3O6PRel4so//RPbgL82hLsKkbox0mK7c99/XMIlm0
9CTWAPa87X6h58nNy3IL+m8qkaauawPYzKjDu7mjgCTudQspemvDv4Ip35vYU0DnrudHCwsAOG7x
S6x8ADZbiTSx6s/j6Xr8EvfDF+4wAOMryBpum+P49CC5RqmzqOweDVqRV7mT0atSWOieR4VsiXx+
13e9nNFTZHFBweOLENuOoYUslvHH4xO4DRsnyGm+9tu23HiktCX6LStjXUlg5eiboo+tIKe+Yiue
ldlDhahPcPUZ6SYj7Z+dhvQKRKSZFGNNQXrC/7i3VmzMpKcx3DgQVB2cq5fxE2ar9zGaLV2P7aui
zJ5XNqQ3aRQg/jBNRLHpwWgCyj5Q1MFBamnT2Uj+zqO7IS3ERPJRxTYn0oZwjWrIrGGEo3hrjTk/
9oNf6IQw41bq2qbxhy025js3Zpfo13SrhhJI9oTTONkg/kj+uxnNJfWOqN6JfXew2Obdguuf9/aC
rYiZReH1NV7PvQgxkkKw6yafI3sgS4PW6hLPGrGrldMKuQSvcr7jj/CbqnAyF3SPwFqfiHNy61o1
o/j1+G5GOuGPugMUaKzLvP6e9nHOAdSFj9NTHoWowGi209ivVjbMW+KUfvKwvB/A3+inQlyeERa8
ZqklnUAjKsZhaH47O7GgnaWA+SXEGzBOojDwYVdXubYP495obnsVc8Cz4UVw+fIYRVIwLDQNBV7E
oONyUNHTLadNArPaEKCOIfbKWa2fBz2wtAq2BNQ1RXMHJ7LwZy0u/SkjhOLoEVP43vYBBJNesJOw
HEd35kjCjTxgV6ZiVzhh5QT34M5YBRUFtCkW6WiZelqms0BOrjLX9FuHwVL3NPjV2Xyp3/0A6yLk
AlxiEDaJb4OhUVHCTw2M4j5wjZXp1IxamRZDXVLfS0K//KwgiwTzc9VSGoiBKsWiGmqJJlSGsNYT
HA6/HSjKDNTCKI/8WDi9YI1hHU27Om9b8PI6HOiKEkWkRIyP6p0g1wMKnXvSQ5F5RaR8jgv9NQgU
MEbrFu/KQ+eraiQXiJDVwnUvLaXAVUHdKWUNLwRdYqVfuIP2a5aBLVYWed3ndI3XXtP6+1yLajRC
yhqOrdZs6FKsM3uMxXa/TP7AzFwp/8JbVJzrT+SOdwE9CfgNWJ2bFr6CIhX1zw9Z9dwJgOJC10/q
2VjTBRo9Uolb7rhNlI3QPcok9YzvRmxPae5LH/wZFtgggh4JF8CoNyx7RMK1LYdeCY0Zc3s5CWW3
0GdQ8NFBsmrc8KZZQ+r7JidYlDYhceqBG+onz03N0esinBEdygPIzXM+kDrRRb70SBQJEXeNbWSv
LBJsYWzhEjeCg5wjr+052RcZvWrWiXbLV1IFj4JcnEal2lb1YUCmdZEaKw78k1hMq79Npj4MQazY
i7zSPXdAJlKPY1MBOSGuJCG5HzkHDe6gFbv2KWKTGXVixKR1ip6kAIO5r/1p0LmLIRHsmyNSka0l
VBKGlYtEC6Opu1a5Oeribgg+iDtEyf6be9XeY0r1x314+LSHNZ9igLenPiAaZ0Oz5sRm046/Coix
MY8BDi4SD5omYWGARkFDEPmTui3lyx8Wyg2HXMSTomD78ACUZHIhTlH7WHPICZ8W9jzO2eNiEWwI
7gy0Koh/k9ExEeGRtYLbtakTSlpx7y6inayotp+ZivqTDinQCzcyBZUT99uJWRpCpppelrRehGZB
D3XUQcGXQDANTgK30Bfs5/bQv4q7c2Lumf6AM/uIdyZ5+ZNcFRqID4Rfb/EskW3iJhVwj1At2z19
9ZrbanJ+ejB7d1mTR5gdbpo4pU738PlsnXxHSh9DUXRMvOt7WSFI63Xy4A+XKgemCww/e6sZp8f0
jRVFyLLOZfWDc9T4CE4V4mJMy+UyEXzlcWrS1n7gSaOKQTAZbZutKje69Uvc+cXpaR6qWf9kcqcD
u1uXO50VBQnyaeumVAWSStqW534YQrsBLXv7spe5gLFMOvKDtbAsklOyHl46ACFquWXtxf0qMDLc
R7feboZBFzkzxG8KCBk0r612vzIE+E6Uo+Qo1ht2W+WRbZOq1RgTV7LmjKhRxJOMkqpxa371G/OD
ATfxwrnZwNsF7eiBptRRUZMPESbAqHTWuKaGWtS1AK05/AXHa6yq4anh4SpTRyXxVFLluaQnw4oW
/sQnD9TgJU9g5uPRT/w2CgsGjbEpxnp0+8pwGcgpLvnbSVKk9q4Pdz5Y1alxPntSJmHCMC3i4myg
fcg2PVjzDcEnjkA0OlS3510TVtCC/md8POP7W8bAPQPmQa37CHaPPPodqGxHYie2DCj2b1Nm5ZY7
tJnupUjuKK+3pRrReVhxROduWS30PVcP1sXWj9BqfVLtuocRObxoP8ieNyRHDNaHN/je7Okqeiir
gMmqzJ0NAaRYC152IVBCkN/2tb06Hwa7xwKjjs1vpTUEna525GzlV04/lZ0W0iWoBsndnD9CH/kn
3KlN2vXsb+KB0BZ4Y+ear0oWY/Vggh4zzgzgSF10z/Yk6f7JKE52zaVxj6IiSPYm+RsXOrjD06m3
nXdOmKbOF6R0qHvxXuwwpGUoSzGMFVFVYCJUob+q7v4SneLYdZAKjfZd42gq9yzGGvX7hHDZbePu
cz92AD7135a/Hc70pHoxdvUH0McNILjLSX738ohNoA9JvsEZoRTPDuGt/aMS1x1b83JZuN635Nmr
Gp50djqMxG2An6LXAk8ryb/IIo/I9WMmc2Wdp3q5i6jotMQ06THAfGgfyI2dQ/2ESvTZQGW3pJzT
WBiQmUgw8enISwlkudJj7HIUQHt1rSYrmivBiFO5+XdVa86GY8FBb4GhNnX/6BMB7IpIbJBaZqQn
C0EB/k0aNuwXfTkNZA+K+kOoP/ukHXXSUo8kZns550rrztfcsubJtj9NknDFSgMLG8OOxp5AElFq
v9j0YNjd3Jb7vl9Mp/xhw2rnLkIaMxCDWt56DcWx6usDHmSSvIxfENdmN+yNd+mWIwI4csxGk+Rs
c28PC95xhOSGy08n3bNPq+1PVU3TAymsdnuH6Sm1aqGwlaf/fOU/gxzivebrBezv2UhOYfx1Rmuh
rppC/CCKCJC5fybzxh2sieggmbaGA8DGGxAXOj5loPH7H8pZ98Ksk6RZiHVHmp3vJPSEUQbc2h4/
DU9enCGby5vTgYa1mHPltKgWP5deHYEhALaoZSop2lz3CET34MBXo2RtyAIXsmUnGdwjto1mY4mj
iYetjAzNJYVPE39Tl+3kpB060NVmT4Tk7aBeW5PODOkjp7VkTZ67oiDY4/9tnAx6TKL1sXbHrAOP
K8QvA6i3wdmnMaHBDIj/ZzdXMUR20gtrpBToNxCTO6755t3v//xAt+LCxyOA9vAhVEXtWNg1mOrE
uHEHaXmJtiqeRJnRf6JOEZsDX5Zhzk13Gm4nmPFKVWGDcc/58/M5BgCgudALg5peRd5yyo9Q0PfZ
Gm3TCohdFR8Bdyy0L3oUpFiuXirGyJ1m51UOr1X1gAZrNMT/IX8scKrY2a+2aeNDZb5+3P+OSBOz
Wzwk3FL1rcz2WAU/LByBRq0kIWHZtfxnkaaUcuN1lqMQGMYMZnt7NQ1t9wWG4cluOS5xgz/RrUn6
pvIWT6gUSEfzfnmOq22adIN6W6oUZSJm4ka7Rc9Dh2Mv5OkciRFRb9Hs0omN5vEbyuF5cEiplSEJ
8mKeQC2CJggXNzTR3HTNT/htZ+Cyduqv683bGnd3JiQrexSDdp0xocJsoEHS3kxQ7QbuDJxW1K9N
nlr6hy3df7Z30H2sK0YZuDBFM4bj1OIq2c8xR/WdXiCvAau1qGqhfWKWbgPxB4/ObnF5nlNb2Y5O
4oz6m28UDopFOSiRA4nSkyUbz9fiX2NnXfYLfdtZzEWot0HrzXSRTeOvFWetchDvx+nENjb5nLVA
WRXfK6J/r6ygB57k4Ly2cW9/ESzsQixLt01lqh+loy9C0QMOdnfBYdkXt7MseKGqFKfHeI4p8xHc
lNCPFB0nFjjCf62wodybbtMKrPktHCg1ncIwsWrWR5p126Uyo2gud+I8ZEVFiuMAKYvk4waX4ot9
kRVgBIVTb2r5DtejP0lxofBh3ToDbxK9LD7Q8IgRmLTnhbeCqitLlHWCTdj4U9U2yj1k8XNWF7bL
Jxr5sVcLpoDNn6y62cTLxg0bybphijZ09Jck8seqF7Ci/63H7KmFAUqU6ZY7BBeYtFbPcxYTlt78
+HA+/1gN6gHgf9sqYjTBv/9TbUNfImndZrahRcI3TWBF5Tu2S0bAEzPSHOMX/u4Gcjh/4iCLge+E
UlmZQZc0TYLzwkXAgAs5DgYihWxOPHK9rq8PyeWlFRsPCzQD8N3yudJhv4OeyRpIHT+R2kafIIkx
cwNk/zRPbo1Nl5//Y4fYWBVyB1WiFkulqOzymzZ4uDEjCP35/2+077fias55s9aE2HYfZ7y1bwll
bs+cxJ93TF7vnNoGig3qVrK6oQS3t6ld/E/fPHoJPS4mE14sO+7ngxKxeekIF+FImbnKHIeD/CXw
SN+cBNoXgIb5cQb+UhT0QqARuxMXlOena+9Fy6C1bNtHokSfYeB8k5t+NzKg7DLLv6YyoEE3v0wZ
zqPnhtBNs5wrLLKX6DJDUUqsmH/kemso3dVT025/b05PXbTxGiOrTLOzaLoGGIdwtGU2zk3WUtbq
7tlgHtatNKSk0X6c84DrFk7GXwEoBnIiIVXTNP6vJe1t6jQl5Gb+4d+1CE1Cnoiau/FhyI4kkLks
4maeRwPk9SrIPFUStsbpNnLDfps8j9WJY0jdUDGkaEb3hWbR9lvMkz7S17H4zvzmBPfHLvPYEGjx
anL0JGvehCfM3FWbZWszITB6VzRxdCCQgv2YiWyvOWLH5aYRYqjapnyEy5io49RM/GOB7bbJzGDS
HySXhJouYmtCPwEG7q9zPCAPzfTLICA1tqdO4wGmTY3UR0H+kaOrgNEYoujZU5h27mor1QWptS4w
h4fvBtNTM+VTjUeQtZFaiJbln40y05qhr5xPlV+nHYyhyjkw5gcMxslUc3CkD87A3ZTwbAlH31TD
pZaMf8RI95P6LkkbUb4qRs/cBSGDZ7+GpGjEVFKF4OkjqL00BYG2+q79m/JPXiM0qGHY9YfunxS9
0BXraFXkxn07VS5GzCjnxZz9SQqgTOLSck3/wwhmrkLYQs47OpmO4kyS6/Wp+bSkAM8aBK0kDLhA
x3d7nSJ2iadt0e+XooVFKXipXItulElKOWKFDexxcdB47SZlCGG39PKjY5U0KsSYix1+DOGBsmQQ
ELPS1ZvXx654aSYPWEOdSz955EF2Fr9pEYW2L1dNqUM8FfZBNAWlRLQR0XyLSRyKCK3yZy/H5PhD
PT1PW0cNOjT7cv5+uI8od+2kqgev1d5U+szBpTqB4xbo0snzHtyI5gTF/na3YvRtbhaJzg9ePQOw
ol19CtyLn+nyumXbQqynRdaO8Cvaub44qz1MgBBjiJvl2v6tUEkMSm1xFa97hrIuS2jRQ2c2dnT2
V4KstRiNlkw5tigaY++rnG8/UWhRvWcKcGpT46Obq3v0Ke1tu/SdOJ2wgI4UpTebuGhBn91ZgZVE
PZxbaImKM4U6cNf9+P8LmGL+WULVQSODS1kHuzNAhCulcx+TdZ+sQ9xQ/PaM3a/SbKXWlRG20h2L
gihCEe91+kX05o9lqwNJi1tYICV3inCY4xadEoCcqPwiITmmpoeNzu8DiomJxOYukIZJfRLH23fn
V5RX3kVXYSsOlhDJzfFF4P1wOeLBGMmjghcznMs+0nu1MQe+//4V1S3q4cJDmHfMLSnLsCpqxxpr
9SBsIUV/wha25pos8bxNdX7crsTEgFj+YjHWIMY5/ij8h13tGkf9LxcfaLt1Xl2UaMu1iaGAOtE4
tNbMHHbTxQfgxL+ACza3haYXj0Lu8UFmEaZhEVR71SpsEq+TcGENl5/JmiF7cyQNT0rPtOPaVXrK
AxwOgxVQ/XfCYEofzSc5gG1bS462ZJo2S9gyWFZD8aZ8jzjHF3FseX+TK8QZiIlGkw1T3XrqJ8VP
rf4c5Rkr51zJOEW+dOMwwPkDH3Ws3Oe75w5MfnF6sPdlNJDx8oL5V11eTnEDX4az6nFnSMXjzwJF
OzolydokezBKNYrvucP/U8Y6j5Xv6KLu981NLa8sw9lKk5WrszvGgsdeQWio2zw2AlHGoODRAx0v
UZx8ugMMKJWotEx7N71lzx+ryKyKP+bAp+jFvom0w8dQvxatl+2nVeBABuFXMCPUz670e6afj4hP
VPb5M1qMUlsyH1urmy4eySZ6j9frjOlyBQPAsGcdC7dM0DTT2513FIlk0Geo2fFxCi3II1qi6vyJ
efjImhJIPlu+AkXCoiCGqhEp6nNKMeI1b92dvpMl5TnV372p8lNjWSPWFs2RZLqggN4kzZFAfCpk
61Foy17m4d4hWGSAIK1jKncZe87ylSaDTm56R4gcUXQaHFrIXRORdh4n+jhEfFgOY19dSra1di4o
5lcn0yGPvnfw9i1FRur7PZJMQ56qfBGbP3JXsU3XOPFv+rsUP/H4J5liqHymVzpXv3D9MPYGb4ge
A7Qii/w/M7eTYI/aXj8u364HWGOf2YWDRP48KHHAPx3rqo6KibDYsBjagG77fvhkbv6+u27B3PD8
0CxToLAiH+W+0KFuTcA19XsCLFD1Id0jW7JuyQUwRck1BRq5MIR50xMKo1eRvQc1NHyvkAp/AUNJ
KkrwKgZtb2/zRG5gV0/RWtROhOLxczOGKHqB7pEL7Q+IvI+Gm61DO2wBk5Egg4363bG5E6xs/vLr
xPtcCzAplbfT90o4R4ZriHq6z4BSUbcpTX8vrkm9u/nGS/ZnKFmzkB17loLJnqu73TmgeDlwpvqz
uzIEngwwrO9+7juMFQExEDXKbLcP3ZiHdaxku9AUb6+Z3o095gYfjWi31RcU7c6X5yFIHc0CKfqd
ZvE0KXqSs/i5Se90T9oVFJ97vdVAG5Eho95UbFCje7ww82IhwE8TkyfEvwUU5yB30+ezCjALoF2G
CetU6Gly0+ryJPDEhVY48cVgg4/7swhhq/T4XfTm3EoBit7ruJrSmnRAH3142SyEGlsV6ZVwo7/p
dcuAWQx7TfjvFsF/N2E2m9RBmmMNWLonHNV23voo4dKGTjR65Fk3sI7DsWvVJGkhs79pHh8fMUgZ
QDSPUbwC0jySKKKpTJQIN+PyPGrTUO57FZt/WjdkBDjPanfZJb/Se7DLXTtxMG0u2Kd4zXuF7/VV
ZBRpyaZ6HCIkoJN7hc7sss3WdHKggemng9Hu1U7mp3/jF1AnMARts15lvr2bEs2/XmijxqfpQn9l
wC09e/y+LxwNaOeoJXLypq/1BtfqDjYqE/d1WzKeKN/4Hsp4pnYs8oD8Unjrpw3JJA5jhs+GEWUV
aI6lrOQim3qWoje+ZvzT6Hv3qDGMckNBWOcR3AHZgKPOistopxc99aLWjREB65JOcsl39ciXBD+V
I+LNT3sxdObsGkRJ9hdjCq1NCUJ8jiyp/Cd++qHJeaWQJFxDkmUntqTJUUIqX3w12ECejKkk+Dpi
XPYJ6L/4RPAF+ELz6FYJzq1aMACUsnN8OxHCp8YZDSKhZEkkY11W7hS+BeuBesoKoF4nBwn0X+M6
AUG5jqYXXnIZr5X+u0rs45uKVetk7lRieROhBXEG+dEhs7XkwF3iZmmtp4003D9aqR5aYuQM2DGJ
BlXHREZD2wsuwAMyHrWwPIg0KfD61FORISXerqniQZjJlyog0kFG4B9bIfcWgNTrnIeoqpChQbZ+
f+g/vdN9/4cgsV8QdGYG0EIH1q7hDU+TizyggwsLGjLc2mOFZZyyzdKf7q/Lx6thoSwYFS+2rXWl
/jRMzGSRR7XthrGYEXzsxZFaq/9uCefl5YXoD6U/oKHNS6RLKIBMC2OdqO4Y6oF7qWArdem1JgCo
vFBkTlG6+J4yOsCzUov7O64yc7xAxTIMBpF6wsJ9+JHya3rRj0MnL0mT93m0jy8dnvo/k4CJvS0R
/WKuJKdPkG7EKQvm6fogROaOrGiGv50khZJRviGBcBe4dD6tr28BLPsj6pUgkkAixZy1m8iYS8dl
MWmHF7DEskq5YQH0dRusf3NfTX1FoDdHBOrpUciv2vR5biPmhiF74dxH/VC24IB9Q9O4x4pk6WUF
vAsCBs6T4QFsUPm/9vSHqleleCGf2kohLf7NDvTArmfye8ttWjCn2mlNju2yklDnKXZpzd8vOW+Q
AeTsBg/SY8t24WkT2/CiKpbmYasDO0hrnF4iZfujBRdpQMnJbPlcLlFvcedMMNAx4I/uca4ZdZy4
OxLAeRyM3LwSxUQkDN75/kmElTlYm0n8fQ3LL/s08ppCIeckqavVT5ludP1AB+yhIJaFDlANBqw9
ayxDkuY4gO6WTrxiHg+A8jkb9YJztCPWSBtwSVY0TdhOlXEczLjZyvoXEXrso/Y2k2pTWPVhEPEj
WG2Cuu0UlbKOVi81bONHv0WIwcJWp/6nBFYdYMHoLMZdnBCv13AdXfuZFija4x2eTOChSpAOqf51
/mTnVB6Hs90Abs9T/3j8sJ+LyBlKbdHI6HiGCAENBghR3KgeBeTNmis2Cnd2OVuNbezfwD4PeLFQ
0IBJWOUazsaG6U6+pVLhU0HRnKL9XU3H6uEjrnIWnrstJrViedEIx6V8XgW7mWHeawvs9l32D9Br
Qpi6Wr3A5Hc17L9S4YWBzfvwiBjGaiTlw0dV5Ru4BvfJKgOQISn27C8SfN/aoTR0bq8qnlX27/8/
M9Bsmu3EuWVN+N/gLLnYjKsZSnFBETeHFSdd3Y8+mSdGgpb8m9paBZfmx1rAUfb7tz0Xwrzm3NeA
2zTnWkjWnHciUUVs2e2Wd6RAjv8m0ejJMVa2Klj0BShTgAMYguU3q+wXWsyg6/wuc8bAjI5TyPqd
lXfna/BR/pPfyZLK/z3Caz0h7Q7UK6ay+FK3TXvq7rnh8n/15cHwHOOhz6aP8gVuSTCUiZGaRw5w
Zx+iUUOPvsoirEUUQFDeta02wJt6PIdz9iSEjiFjofoKtM+8I6XL1G3NpmogqiDngLX9q59lgj7u
Dy+pjPcQCOJpo7SyRTjNMq5nErgRWUPyo63WV2cKtMPf+0Zgy3Irub6sHXF+FreC1qKGI5l+B0vE
qnJwyNk3N0CWJh/BzmQMr3yDXSQAjUJFn7uCHLqJEljmKppeJBXTGqKHkDBQK4LyLRWVw+GTQeFS
qyE9HmG8hpWnrCRe8lWocJhz/8IL1upSmy4ivSLuJaxMBx02UFfoeajsvzYi4p9LiuBti7YHRcac
8GDVuMucTlugf4yFUoLUvLbWO87EyB+JkVZ2eIHyOtYgzDsOLdp22YmBmTYSxwuslUVI52DhBLh5
HrGlqpVg9NMq8vVrDWGxVMKXpDGZt7e+lyYjVXhmMkGClYaDH55Mc523QE+91k8RLisoMFTM5oK5
3z9drF5ofTe6FAuRHns1n4c7RqMqwKYOxPlzl+lUkmgvHarj18i1oUiDcur+M8btD4MuEK5BaIrT
rJdUPTh/QKWdXVM2XjR8+asdF6pUl+HZjKXKME+FOrUchjSDTPhTHobLhb0ZgH1sn+O8fw4qUy27
sP2ycai7VLmvQiUFjwAP2qvhzy62gqYyVNNJzlr+u/bOrIZEHmbxGg+nFt94aHa58lz/uOQ9PvTW
UADRV3tsVqdIu8rXIafWY3dkEOpTDOzKMU4jVdpiIE27kyVWaMJS3Hd31D0XRMovlkPQz/npU420
vgy7otVEU1o0C6WqeOx9YplzVSWcrLYSOxm+PHb+PTXXK/ZkyL4FVZ1RU1iswyi6Fp1QXKTLj859
UkK8orL5Z+6qxJf4pdvOeDm6ku/x9ja91tF+dq6/WU5no5Py2xF2wL9mBiJqRTo4MDAhbrlHJNHb
aOEjZcwRbe+kGoxlOzlwgEf31GHkKNXsKCdlFaaQgjC+9YUQ7MYMXxwghafAOJggtX+FhpiI/rSh
Y42A9udwJbidzD2BudDbRKrelaNwHY2on4Oxdu8J7bqVquUt94sd2WAf251pwbp4hQI1XoOjDMaI
8YRlKJT1tnwybMh/SWO17txuuO6fRaqqbHi6O3fmJV/4oIR1n4jIrCZ7Hv2xeqkHAw/MaNILMnl2
6ybVZFqNESDdbQU54sqq6DjAnj/2HWeX4vAENShr2TMGp5GZ+XSR7bkq3Dyy2l8P12EIzQ+kFYmV
LeHV50Z4vQOvvZeypow13rA/6I79hsj8MKLDAJx+vBXaWfLNLjZDvaj48Bk+LUvo3KgvTOYvMod0
MMNOc0vGqTfN/DcjE3BX+wBNfMAkDZyFNkyooLuH3A1HXVVOKz5ucHR+UT8R6i3ooxMYiuP4xMRW
T8sQtYlh5V8XRz20Jxum1AIIoMO1kW5K92JAmK66g27J/u1G3uKX0M7Ae1ZbgAUOsV9rnU5AEZR/
7VGwfPPq2s9E/LGJHorx3cxCyf6m3uVgO8ENo5AF08YVKcsSNv9tbvRcDC57ZnAYYlj8b0FiyqwK
imMSuVIFHCUTKYHB72cFs0x78d5PpVHlsaTet8uYhPRq6U0ch6WrD1bRYR7XiR/LP7bLcVRthry8
iD/ggxbnfSOdz+7fPLZw9Xi3C95dHPYszUFFe6lwIPW/SniefImsXhH2+C5+buIdhIJglBPD4wyO
Y8ycxDrF2PF9iceMPMBTk1NM2G0iwAUPYMGc8ioFQqJ3PRk0bJcEBwPiNmc/yXlplIuZE+DwUMB5
vGvbOd08JZ5+q/bIFFsOA5TxBSniT7pp/zZIFMeB4Y/yQZZ5Cbu0QCtVvKywAPRQVHlBpeeLRzr+
C4Es8GYBrJ86KI/gIw29Tx8ydtNDs8c6oAL8q2S7aOxULEcDEgSwgDzjtJTqRbX6UxgEbSg3pVUF
yyNbrdQTpva+t+MUmfN2NKHSmjYM1zvKpSxvphm5VQErUlpvONQsqCKTsVJwwn+MkkSB9LH1wGsd
siHN7VEEFCz7pzbE36ir8ISKnTQ9fIKfESAeqBUgW6ioqvooQIZcTLjpf4/P+TWhGMnAXv9gnKsk
Iih3qjg0+/pMqGQcXcV+lN0+59lxlhbAhRaJ+gnvu/1fyMjVoqRPUfPg2OZ/mLZx3Aba+svp7wIR
ly9t1XHXu4lCvVmWVAnBpPW012Nvt5uJb7mIvJ2thHenegpyxbU5gwnl/sR2fhRw/NVinRqjqWpS
UNMFH/viPbmiW1WI4z4Zak4zNtzL4cZ5+E/1Vl7GOMv/1suftSGeIGAf6rAJCOxdbzmpMdKXZxKV
tM8Y2QOX7aOgFMBiFFvVqIVzt7topci3D5h0rNf0BfQ6/N5q6FwTn3VAddKAKFS+EBAMpPUlTFGK
Vyg+j2X/eRKQ9uNhRlQWQplxCMKj/C3UQkRBKPsRkRuZ7G/pfW6JgINwlyaPjHhTVQgc8VKaEwyC
Ssiz6/oIhspdfLGsFXYhv/GZOGvfJk/NjFTtXM+V2Xg5sg4/zXrnjcZxtnk+0M0P5r780EZGhki3
c6IQLlRbg1xxDYqnNttjz/B2lFZkZZ3g4OJvnGZTTvL4SQ7gnAjMlkhNRgar2vAq6W1+20TaRIhq
Ugh0lNDWMM16Di96ecmjtbLCRX996uVmchK1Dg/Tf4dV3bSHzmVqPqDc5S9htLpvd+FjBf4wGdT5
n/atAF/D/3XFLWXtJTbXGwouGA/X+tpsRYS6Tcmj4HUO75PkFR2E/wK4Yk/Nqcyvz2C/8FHnogE1
9GER9EAz2n8vIVzj9zsZ1S9x4dg3kU/lP8OdaTxkA252kCdk+QJw14qQAqRSxqFuXe90EByc4wxf
W8nHY1Zt+cYlOP+yefPxpRn2XW3Lh6rfsZsbL01kM472xCtHCf0bOyzyKIdbU6O9uuHdGNDEgf0Y
zm3PsAGbQrTIdKN8a3L+JbeK2HBHl91MTyf88j+RlMFwZrYm9e7weYJr300WUXq5DE6+lPUQ69kW
Q3wRcifEfxaYaJCjxA24jCln93nGOOLLfizieYfdCpdJd8l5U4rcAXoEh7Y4b8jeb0+w/ivKnNgQ
4c9KXLtTWOV8V+VoNZkZ0QTQg9Be2S0gep1uv6xD5nA/k3fcfcoqhzCoMSJiqAgeTYXkmTy/eJyh
Utpl9WTvy9SYlfUmbDgPK/KR8NstKWdinLOSiEagEg2KqaxMQijQWjv9+dHbeDsFNEJISNEUebeK
7o1H6yzEyVboqWCXdMyIe3IM4aoZKCm5XikF8QdTIKiKLknDFrzbcDb0M9Pr7CVixGd7j3pxaeGH
V0x0TZ4bA1LBxF5UHkq8JUv3ZhU0AFPNMbTRGzd8WfJgOmis5CtxaLYJ02SOaTUrE+vWzXmjU0Nx
cV/SmWz8JylgZhM/1et/50PwdBzBFBSKmdNvqso0PBEsP96ikxJUM2DXx0ViazzUW9JKTsg8zjkF
JkmeJZETNVd7xFZ82D+xOwZ/Kg7Z4ZFJR9afxu61l32VAGkqVBUVEu+6UKlAIMh5JBZ9w/HxdeXF
ypvtGIf/ws/Snop+V7NnRm5z4cT3KGJbuytLndzh69kv86ofkAM6uXxEj1gd64SmyYRHII67B7e7
QwaTsWeTSj0q5sYaKiVigZW+r02+vNQml5TEMC2ysKr7RMfTiQxoDvQA3t/jaxmIXNpf7C30U40K
oRa5koBpUug/MS6bubCEHDY7+edkxDXimiimrTQWzVfgxs64YMjYBabZndk06vZaAZDYsdZkn/b+
jC7aTIALfCDKfK/NZZ4099BY+lHyokU9UANs0rFeSyfJa51QuiGoDFfse2RpxRMnDjFfdtCiryzq
FzSPuChzsDO6LbrIV/YMRG0g4SYOTZ9022wXzCPzg9ysjzrBeHETE+J1yTX/MsuU0XHXjz3suyHK
jrNf3y9dA4wTswtMx0aYcQ+TjhWX4Nnps3AuBOq+1v+ggpUfPDBzd8ml4DPQSX2xv3qbpW+Bo/Fj
QGxChHIynWHiZfh19RWTYMSnD0ADdWypzzLDK2UnaGgTb0sfMzcnFYUu9BxYWGU4aNy7sz4rAKiH
EfUotmF8S45CRsY/80o66zyi55i8YszxOugWGMpLLdTRS/BTq7OlapqjRDhXZ+ykL4pXma2wfYjl
3qZpXsCdpyxZZwZC+sHzVG8Zh2FROEJlvOiFWhWaY8fFQAsl9pFOUEwnC1xw9r9jSeK9opUWEVMv
gnArPXVHzaZRYQkuIk+6A5iYRa3t6cxXUeUqB610Gx7LLZ80JUZx5LDR/fOsusYG9UdV4CUyDTGo
9TLRsvx0duRt5+le6m5jrpwcoIAe5hGdUHh86I3Ce3NX4psGNOcB8fE5lEb3ebHTAlOYcFCWvXzD
PIaohSmD/43cFNijP/pMZchWO6WqSeaGl/eNE1YFj4VIP3zMYvVYJAmaxj2C85SaGyjHiL6gdlR8
UxYu12JW3H4qojTy+6cOSF5iysWpy68Q5EXNKzN8hCcskm6yreCcR3IF9hOczEJGSB/KXR1PXeEs
dCCYfJwNxz12bcjf80afJ938Bb5kQJsF1WDNovBAkA6xk0JEfzLy5QW2c9dDzEply5+h0AqbH6OO
XcCfTSVyDEeI+OFqHcTaCOJUpUDo+FT5BEOgpVyv5pKIbV5NOjzKRltxS+AWiCeXSNC0pslciUae
DVsbfFuwJJUY82K2q57W5x7PhKGND2N/P5E3DrRMiPjULc2OKw/Hg/7jVWlOu7cyDc9cLQBsIb/f
jPpA0+iVxxbPOP4CxiFYXZeTScTMG1kyPQyxybMwwX7zDNPeeGeKuY0MqxwH5Lrylze8IApsQRa0
T/ACkek1vPFgJPeRfZbWycgwSGXFlJ50AXCZvuMDdPcgmIHFPIy2URAKqmbjCGdKlLGLuYO5iwjl
s/lEyQeZcsiuj7D04uQqqoYuZ/T7mSJo8q0+cKRyJD0CILO4LhTw3wHfXapOstjS0H28Kw0ubU3w
/efrCwKHSJpO1WyopwhyCvn4jvgxXnjJgRjLwFVMX49gaTnZDyBLMrEx9aSot+p8oIQ4RucQ/GBH
Z9J7+hw6iBae+NS+nDcRTp788Pw1ANmQxhvv0alJtsASYLh7BRUd3GvRzFheoVCrzO5MakNa6DVV
OkOkui9OL2uaK1RBQ4xdIDAjEfb/9dr7x+vLsKkaSaIP9K6cub94xqS3sxRWmv9h5uK8I5ZC/Fno
eZECJfhv+Q/pk7B14/z6Zba5qBUc+E3yiotS58XmDsRmwFUTU5ENeO3WBFTbNRHHaEIwwg48O5oy
6vb0E1Ba7G3YuJp2hsdmD7N7TRSwA6RZq3F0Di8yAYA5nnnIMFrhkHXd9m28QoXtoaIa1CZ9a98D
86QDkDK4fwbgUrSVWILAR2lKhQ+S6dAmz0pnIvUSDHJFDObQCwD16iBIoRa9mz3oAPlBybcmG+xS
26usJ7eMTGH4bAde5NTjpZWAzjCcWpmNQ3/CzhBR1Oj5LocV1l7gdZjzqXXg2Fo0Owb/fj0Bb8gp
UHc8vmIcBBGlJVht7Z80JFTMmvLumNKykQ0mHLcwcroAKR3P2py3tbPj9phcj66K6yZbl7vkecSX
qSTh6Ue954qtk0Y/+yX5al0VlxLDelsqUEY3sK+q9DTuWlxOariGRNeKq/ZTN2CJjps+dOoCa2V4
CaJY67uFMwvtGx+gL19km4BedJTCY9OEDUe/3n3WXvdKP0teKPcwaDuVn/oONq4CP9hA3FUSbDfr
zULE3/MeMY2e1OjSn5+FlKP8eXTD+A/4zocYPGRgCccb0P9Xy2IwtmN3SZdy2MqCqcVyccmUcXsF
J7CqFanQT0WWc8c8PSZaSFe1L7hE877mi8wVm/Hgf2UtTKK2ubRadTsFPDLiOTZORnLScRwL4Pwb
kcWi2F9tilStcwK/wl8J3DAQjPctFSVjtbzLtOVxGwsaXkgtgK0RayqH2GgVABApPoLa6SI1fjE8
CvdB0NE3KWpLCIQExhAASvf1a0+aG6AAfqMlLKg4y4pFRVE4PyfW47QcUn+cE8ktfYr1zrQQ6uCW
24sIzK3L+Ra0KDCDCuCx5ogzZypYn8blVJTf0d5LMXkSe2xraYOJcTDMcBr+gg53XyLAH5//Dcvy
Y16kifyKM+5Vu7lmw2AABlVPAzmONkc2CeF0BhbRN18W/dAoGaqFEYf+XyoIT3SoKCeZkmJ/5oxg
tMEeh8HTCqeZgZ9oFIzb+uYEv8enbvWLXV2fcbTawKt59/2L1oPa+xZqLAZDJHQEUKrn+mWFezsL
5bETvbjCwDAgXagwnWAMXJUWVfGT+0IynzqhgFYHdAHjQlH2OqTp8WbUnbw2yf78GFYlBvN/VrO0
opk1lvakujN58L76veFZLK3Uy+61d99jwa/o9FIi2logS6HiTYFGpGOyIGkIgzMY6d69gWiTP0WP
ZL9bVW+1I9CGIXuBNzOIBMTQVTkH0pKFbdF2HT+pBXnQet8bfMQoH9K2527xAEfp4FTceXy9RLeF
LeR5QIDBuB1PPUpubnEgCxZLZPVPlyO+78wMbvWBeYFyuvg25CpqQ9SRVKWjptEbGXwQV2Zeq+zW
5GVkJu0X9Iur1hF/75o2LjSOufIt/d/V9+6vOWMK3ZDe65DRB9mWxdjzelAUxztp02SB+oukP7bj
+1aLbCtlyyKnaJOx9olgnKel3DN9rrN/RWjI8XuOOdgZMJqu041gOaLiwyL9aYIjPMJ+w4hrimyu
qcGK2AgBOFItjGCrEjF+mVABCB+VWDG/IPc84GTS+i15C5cTV5zaOEhR6pFKeQf+qqdsEVcKJALm
ZwGGmFURxXvx47tQAdAwxzdsur+XsBz0zGMlfo0MQJ0rC3cNloVlfuuma7zhcmlGAgQP3H+Sw4Tz
va4d5E9oSArca//VvnlCjyup9QD3Q7AtDS8bo3U63Kzi+z5cwoA99zj4PhyNvKZEzztrm/rhnE/I
bbj5zQZI8ybnawYTusHG8w7A3XlgUi3fv6CWBHwobodsGpX9P7YI2SgBHG3jQhG7VIkqtTn9KTNV
79i3iivBesW6dMMJ/ihughE2oiu2pX5hahc1dI4mRFO3qY1MJCWW+oDkeagV+x5gNN8Ip0waL63t
HdplXLEtI+yCgaJ+nfzBdkyWR4YBT80u48lPxewj5Yx9KPU0rwtYU2rcVUE/Hkqtki9go3JRquU/
5GNEGI7E6BVLz/ghuHucIxgup3+HvmzRkdvxnDqG3GgFCOdhrz6eYVGE5COxV/HpDMbKeN5Auvj1
UpkUDAxQm2mbNvXWB7vnQA3pfhZzEMpidSUMw+VyxpZjOSkA+r6yZnEXj1QnZukxhIL3LiDueJeU
pitXqQK2LS1s1p0AJbcVrfvjPgmNXe0qzw1Tl/FozJjXuPW3VTGme2DhjDStgvL4UKQI+RkpZd03
II0nSaum4neh3PcLzH3rWH6feS0b9QpV7LWE9w7pOxp5J3U5GTiCUhKGNwCWdH8dIq5tDZBWBsx2
OeOE5rK2rsbGWTLp8iw3Gq31sH5ZjbbnARzYxC1VBcqBDBMFmaQA3z6tNGozTvuPoQG3Nw9z+y2f
zuZMhWhZJXguIWvKSOa5ag/vv6YABUdrrPXuAsBg5OdNzh4JhDoDJecLvatyFXqTYFiygvUuVi8A
CGfb41hsnxBaHKF3sv3Al8KKFD0ZGaAjwUWM9YvxLk2xJVkf1bfpscUX3uy7q71zNto77PGobbIw
pphWHm+VwJZFVxg2YwNyB64aclSWD9n4Hgs03S5lgdmYfM8UyciYT9iY3n3i9OgZ1nER/FYDR0aa
HsUO9hnYpSbZ196pHWyCEcIdzdZSt7JpHGjI1jN7vYOkcyNh6SU1QcsKhDHR+4qx720H9fYphyKR
0G1JZjHc5KRAuLYx/5mXjwj7Vj7Bb80Qz8ogMKITohgK4wMnF2jUd47o6LYNYaLPQeDWJ414DHoy
hYzyx/9NenYLe3QwFtZNs3TflzIL2eaxhQgDvrPdLGCa9pK2ydw4tKB/62dvUoy+A6RZo3TUCnPb
MP7lZJky53JmAWdmXnclBhmd/Iq+LXRxPmhgh4uHOnzUX+YC4eLZ0i0fHW8G4NhQby9A7KzBFKIC
JRiyRMHCty3Jx7uADUKIkDw8XjGC/PzO+x6G0bVeE1ujUVO+pMJ9g0mHFwjIjBJ2jqCYQgSka330
2aclPEzvUg2q0s+j0AUq/splGFPymR72uH5of7XndoAV3YEytWOLzbSh5bSBaP23pJqRQhmsYPaz
y5mq6BtaQb1X+HiYe6njZU8wg4C2D9V1/eO3YhyRJHGu4uOOJLA59e7t06UNb6R5ShDuWW7K5M8/
NacJ587KGDpaFkNST7b63cX4ZIPOGDM2ZA8z3cpu2fn9Gzp/SzuYZtsn+91eXkpPgDOZHzRPBrlx
xbsa7DOtJPUS2WFw/wUf09sta781rPu/cwn1t8q18PFBtdkbxcQqn/hRW7m+4ZwM7H9PCp4Nrgud
Cr2T1WTHLdbdHnRDjnAX7oNWPVGm577blTHW5VCcor5N0lYW3Z5R9qmTDw4pnSCXcJKXhSUVKdST
6g8ZbkG6jWADXF1pPjpq80+AALsKeQkOtL3eEkAoosTSiGQv9Gs+kgJid2o29nb6F/uFrsRxs931
sZ3uQL5P++b7IoumFP8OJEBsAgWuHKTvndDQx6NV8NmeDImx5ZELL4XO5req5jfiP+k0qqMgG1dt
lRIPsTJgSIBMG/O6FqzoiEvKuDSv3NJOnjrnWlgOOTD65H6h1JhjnAh3rRlOczaKLkzuU3QwTU5f
XMyk1JBiZ4MdfBN1AO9ngcXTkL4auKSU1eBxwBdvcGf4kWd6rgd6PKK0EZee68dOJOhrH/f1puda
ymT+4VXzzacyrgDCWUn1ejhWoKutVNRynqfx+kApycd72qZGddqzIaDQXIuZmQzP7S7zaxqbDtaD
ENlyx4S1xhWPjZ3B8Us59tXxMMehTisPUUWkiy+pP90NlZsXAtA7Qrix22Vmcnbg9QLMXqL6MUds
TeFpsdMQ7V4V1ozoNRD+GCXVH5yOPN5F/Y7NxO/3fbPcwb7Oqgccq5c33kkZ9R7+ELzKU16nzGBj
2AB4w6x6j4fKhjfErWjXgnOkC3HQ7iwO7iepdcJZIlX56xObmq2mkFvPMuq8cCIOUZwuS1g6YGvA
7cq9iZcG7M5+SKX4oKN0LMAaJSmq1QEJWyDQZ8Ryn7Pq9HTjKnilvRjSUu5D5tP45dKIprJniVW0
0P4e7XNPvNvVAjFVstAJpCUkNdzrvk/8JRBWDVRoMAQdf68ZGKoFbWo9DThCy9DeaZosBwhs0oMF
bYGD1XlutYfeyxJPW5AG8Am9CuYr0JDOxtCI4/8+w32S4HE1CjzTzndwed61lLglR3D1V2Y/c8iO
6IOyy5dZ+Zvj0H4mb9/vq4ZxTeMqHQ/nVQJBI8EPvWeKKyjJkAeTU1tVUym6LuqXFtIiQ/7f9QjN
/azffr71/o1I7YLUHNLa6njrLDNtR2ONjfR47OrdI5NqI0R5kSZC2auUV6trG2YSgEmzYWyGPaBf
PPjs0weACHK4X3MN2eT+35L2yeCAtTkmYeeSiubMKpUZORvltFbnRToYJkpBL87UWu0qpA8KuQ6/
yOdHxsAQTZzevtkB3H/Ay2b94mh5gNY9fiEJOze931S4hHH791r9F3NuXliG49h0naeoWU7NCHYv
rv7Y5X9K2SLysEAaAZ4XuN0sB/t/y3b1Zugrpou4P9z7NzRJoRM4iwfA/hrJ5dcpT3zdygBUlduv
3XR7uMyj+i4hOU/z22jhYpmesadrUig18khKpvsch+u8urmsibjHFnvGL6DARUzPbWkq+YjLK5kf
GG1oCIDAICf2TTDvHUaPBpM33BhctYXpiuEDFtXYtSIixaonzbV9tw6tXrmS1MJEjHlbTWa9aTSQ
F8y6AjhgJC+uW9OjxhfhjC4rBr4IAuiHFGN/kCy30uIjGKTecPOt0GbwDyUuEeQvXM759ONxsRwo
cs10qiqlGS77edaeFGomsNETzzC7Hjg6l4yCVFWx3fde6EYMfzhnQGuZytjQ51v3pgvTzNcLjd9/
3+0wuMhF/T2zIOMsRtrMLEnW0H6b8d4Eh8C+SiEM6f2dH1deRsPSqfwlJbXQLyNIIXMjTPP+j/pY
bKzRINzPQ9nIOn6AKO/gsSQE7QtoKFAatQD9ziyRsS/RRXu5DvFjoUvCJuVDSu2tTESxBql3WVji
x34/eyGYwR009KDyXjea2UeMWEmju43CP7trwLmqYrOc6Aoi4yb1xO8S1HrlBNqzAdVHYClWj3I0
Zny9h/523QcW2gwRzUKnw5qdY14hWlYqtwnrvwj63dASEm/JkcW7FkxtYe+yjsEa/lKveIxubeGo
2Tj83hxJTTQSy/uUtb8KRQ2jaPeza41Zb3F6osgXPV7blaBJPvVa+0FgQ69IoN7T4rOCuAOVBD9I
sKM9cm+fC7OsKi+U1Rhza6MWmlN8/GInKAbxYRKXn3CLl8jhZHEzktWtPuNQmxwTGfTWNqKtyHQo
sWAeI96hMIXR9LVr3WGSKzzbFfo2AbblLYxAymaTlqvxQhJlKqI+UJ7WxeXxjRn8XFmgcjLGmZfy
IdByXWHOYqxb3ffiBil8weAHzyX58NpQWRToRn5eJjqgxDJ38qeoI3q3kOSF7JchO6UvvEBfe7r9
y84SJk3JCKIPZiAb0ZHbKa8dryfp8SRM+G+XyxgB+JvQqVpDMcQoVot0HzuiCiq8eQ/qLW3x3ZcK
hyTwl3Kw3UYqeOTFgSD1/Jicfh4yaBAY0GFwg3e50ZUHF6Y/3vX1QegRXU8X+h7acKk5uaEJ3yOB
8WWteeAQu7wnC7Lvd/LPRZx4JIm2QFUcgcBVvjLlcfjLETjztkMpZB+gPu3ZbVh2BZirerQmfrAP
M+HSv0zOrbakkjdsh9S5Dj3hSEaEloTuFXu5k6Mz5+f5C70Biyna2N+cEh7570DV7J5OtvhHpO9K
j35qhhw93Das4g3oPN0bUWRRexX1mwIK8gnESzqglNgZIpNXZb/wKx7YSi49ZsKZVKFFkMzxHNu2
5EC4nMJ4sfe1RHLVdI1YTmQzRHWKVpMdLBKFYG3CmfV5bm4VNwSxeS5Jw657B69VZwBN01+CZdch
INEvhBErTUzolMX6odso/8M7RJUZIlR/WMKel2ERN1w2jXQFegFS6jv4KY1PzZfuBHIqfIdHyjsn
h8B+S1n79MtwKyfSwSv7R2RZDKZn4C2cyC/ChonBCDs9vuv2kw6F0PhkTe7TCwHNdoEqGHISri8I
XBCyxsBl1FO0sH5FUf2Jzrmr8znFbgt1dnpd4NScjyidBuoAV8hGvLwZnDxxfB/HpSNACJ8wRZoe
yybq3SQ3r0o2z3yu3kqb03UEOm++PcB9A7JCq3sDUvSIpb5LGWPWQB7Ql2nv9wlWlqBrKGuu0qHe
3F+oCcy81PbilwcgjK00oxo/iAbjEc0H+HdUH/iVe5DzUWffNq1okLV8N7QPI9HTCajyiMX5JLE9
C4i+Q1VGKUvYZSNQHn6F17QhnC5kEWmkDSP7jX22TimlR5bLjzJROjYVWO8wc+iWVYXuuda1GGHd
xDp4XZzIVFXrB0rFhDSnGA7hStkAgYguJMct60ho02sKSRIzdrrFBEA/pqJd6GinSrs8c9xnzF4G
KXmH10QEXAgwHmpbb7HVfWIpfs93Ndz0oE8I+Lg+3Qwbw/2ilikdaYBTFvqHzTXl5CiFMKoj2M/E
+oStqR3VSON81Vau8RG1Zp+qzzB/1UnNbvvYTlZym/5c09/8hhKfgAONuFN2opsnJ8OhzvU0GrjO
ln3/d1oWH+kQDxnr8I/XJRI/gvwfa0Ggdk77g8m/RytWdmZlL7zSJ0Cv1vP42yXCfWSHW9/2C7fp
2X0J2mlBw7YBWPKYGvkDyNKVJFLtDMU+YFU01nsZzKVbUuRkRHwPTuaXHci4rEln0Aa6UVDC06S5
n3p/F28ayxWRaphacJaipBJwhN/YHB/U8NtBs4iSeNzpj5Ummvzz8uQVvGcH8EQvwJvNuKDCu5c6
ujlhsqih8QtfXYUp6D7yWwTa/vnY4E9B75+l4KUXm/2+4Buv9Bd1RmzSSlEhQmdGBMcCGQs6PJdv
PrTKylbT08mzVIPE+Aeb2/EMHRrHDgPgsvQRmLAZq8X95hsi33VqqiLIhSUaYBalpx+CE3Lxuez8
0rECqNH86APABY86wfYeQSgIBXghyGsqfb11DPaJLLVgQYf71u8NthnR0ph0xhxvM1hUK/HTQIjU
2PxA/Wrcfyu3vQUbypDnjpa4LQUwaUYgfEOE8i+PekqSn9NPgoG4rLajiwEt9RNm+V+y73YXTIlP
MBA9IwSFte81SIfJQcLJsozJmX64x5Y7Q6//OQf+lqioOVM5eVIYFuP+9Z3UpYCKSB1A3kmFBqtZ
Gy4aySZzbh/YheuW/049J5+sAicZ1tYREUFExnobUA2vpokBUb7Jd+1cSBBCVKF8yqPwPfA03HYe
FotojwCZB1BDH0Nizxd6ldoLyX9157MLFv3L+Wwt8ZTYLRu5D/mCsPp44895XNmjFKqP4WFApT9p
60pSUlajddHASeOQETpl3MZqC2y680fEtWeVYd1xqW3NGXsMD7ICFVUFXWBlHNSGQPJ8FnEgMS6Z
w17b1MzKivn6MXniAy3kAXnGTPcCD6C5/dKsAqx742i90SQPBy6UUFQW8ZE0w+2VkHEUbpze56U2
SYBGK4gYOdg9+QXrqOcg3Bi07KDa7wT3wKZJKj7V4sqln/AwlP4v72/YzGdlsiZ+IyQMKaf4Gybz
9QLpjhcGBHG1hGwqe8jr+xyJMKZnZh3DsD0oO8Mtj9Xq7Vy2EZlpSvBpcUkdpK+RjiJu4q57mlEm
CHMcCb9sxSUeD+s6WUqPN7OoEmrUjyvlMDbWkMd3Q4vsrLiug60w3ty3YZTyYSKRkykBKRxxmxtw
S188WhqtfQfRmzTtH0jwQ3ctp2JgwLeVQFnSKr2XG/SCLovu5C6WZxqkyClsqCGV8NVQZ1p240U3
ip4Lk93OFBoZlBFvlFBheRkK8lYWxibdGzRj4uvFIk6Yc5ctE/5Jaxp5ZCoRhdr/1Q5UYErLs9xF
NrhQYTAm2ZryTcmjV+JJf7OFKeU9WlfR5bXcIqzok2GIt0hgi8T+9Zrtpg74Jhy6LzJlIc+EoiGg
1Ob5N2ZD9BrO0ULfwy9VFKQPN7kSEHb6OZZk6VmgucrCt0MqxvmRhhzTIWEucJgOAd4BYAwDBsNS
rRChlMuwHMG/gYebyawha9gpwoJtbtbQC181AOjDLN1IBvITM++jn1KoxxGOUGSytktEfbTFgmzf
kbl04zYkUt5VWSlCkmrbxBjFz4eO4B4YtZyaq0P2eqUDG6f7rvL/Meoc5YH6cCh8rnZKFaszqvnK
c+V4YYH0FDVE8TC9ZwbD7V7uHOQ4939PrnH4ldZrQa28xnGHUECaV53Zuv9U2G9+ePmAm7GHdpzk
psYZjZ30y+qYNxzrtUGTfC/ua3r8yRDYZhFpC8E9y2FEFMxw4H6yiaxiIxRm4xwpOUkVUE9kRRwN
xlPyeuMrgVojWO5gN3mPEw8ZkHTdtC/219T+plgh0Zgicr6POkp2/8Hiop6SLBJdWXd+czHLImr3
lnX3avSkAqUsFc1AFXEkFw5hakJHHCDrdxiwg9HqmP3j1PFezqk5FESwOihymHQKYaDP6pgjiOhV
Xg3quhIPZlvkS6R2vUpuz2eu7lNxBAuRL2pg9wR7a8mvtTgfUJ/ISCYW9TwF35mpzcbXn8MKInq6
Lrqumzg7xEI8a/CgoGEeEEcc8x4iIla1yUlDJtMgxob5KTcg8RXZF5aFiV6/ahYOdilwL3yGesJ3
TIfeGk9x9rNNcpsrzkGUgazewNZ6uKRawS8PtkwL146oxZwHI9iS42NhBWT539tflhhmJUey8sH6
IHo6niqx4PGNPMUO27nUtFp0bC4DzwCB/865FkWgUmpP20Rgvp5occLVScSArzW8lq1RWMkcSYyj
AdRYlcdkWgLpWg4XSAYsTSfd+cvWFmrochyBOel0jFduNfPNuogWzz6VG9wla8WL9+mX6gSthVzM
Z2n3HQMZOpOxWjsI3qqf9mfnEH5u4704fi5fRdPxTSTmHnzZepvwSzNKqd6QmnksdTcK0aivvoJu
CH+/jNJckGOU3CTujEcocstv1KDCWHv68GxW67qZLqTQ/txD69Nv434EJjhoUNV06AbjC2go77gs
ndIfGNuUxKlDeXddRQZIQfgf00F7Ff7j4UtIJ8vvJV3H0RLv9Blx6gP6LIH3OtNJQ19F5CCXnorZ
Pahxgs98SZWCBHVL3mbdLxHMvaLtVROmXgEDBhUcCP1Yi5JBgDNLm3XQSsB/bBEveAi6T6a2BQDQ
JO5Qh6GYLx0uKMUA+fpWmi9DrQQ59yN8ZFNTB4DUsr+pFmzFkYuz9i3TmHRSMJTQ6SLX0D/n5q4e
ksFBJDXEyLrae4KR6/8ih1vNdN5WySKKRZbQuorFF288i0kFlJ6O8ChbtB5Mpv7cD4wTzkMBaa4R
L1N7cFPkux7d2gJtnpvoznjmVnaAen81rsPiidha7f70zrL0AxXGurB8g7Ma7z32Z01c7RVAbfVu
BPBkj68vVCCp02vvfmSScLT8WO32NUL2vZZUo98RdilES/Ym6Duqp1czP1SIKT2qHJjZR9Cq9fmW
zcKovX0H4cubCzAhAeZr1/BvEUMJR1kND9zft85XE984xPQv6dp4w7cp9Wbxkgypl0MfFqMqW3Z7
gPmgFfe83HUtIMOEXx4rOXuR1jMEqYPc8i2PhMOwnyqkHwCNa8NzZQW1BpjisWeKXa0rYha8XE08
xIslr/V67Y6A0NtzKS1B3eePbL89Cp+dPYoffgzm8FeDwdBsYNjWFu9I01ki7rtZFqq8ceGtrR9k
sBpU8w3ncuwnH0v0U7ceKruB735ZvQeETl1El3x7fBEjaPqSQS/b6jcwneJwrbpSRRD5+OkG34jJ
KL3eIQlNK/L78S1vgDTvXb7aQfCMp4cvsWAXGx8cINL4k6Om32JZSAROgUmb3WMEZF1W6tFzCLeW
qrIt8k9PJT7KGj/7NYS//e1AlOiFOSbfRNCSNUodvt0hxJjEff2v9MPcaeIbqJ74rXbWEIOSWF25
InAI+mQsSZqfJhahdfIOjsvsZx4g8BNMF2oB8GVKdESbTVTn4/CM13SemIS+ze+mOycV4fCf/pUG
DKjcbNV+Q7wMJ7sSsVaAdd62T+a6oEGXzq4Ty8jKThrakIutqpCa27HxTp1KZKWitbkjrkf2U2L7
1ms8+qrcakwaHfwhWiHuqFi/HmUQ+8PQw0+c6dEI5hnhN0RDTnVZtRVCbbfoc/GahNutAlj2Z7M3
CTooiVEC+GTnItXOetkRThISOf5N4LSEOlpfGRQXD2WgQSWKhyNJV0PTZgVsk357BCiNRXU+KrEi
U3RVF1ZS9AJzK5uJEHTzJeKovWQiaDdNQygD5E6xFW24ZASRU4k7i0oijy2P0+mVjJAN30B/WVBh
8pVfpnRz09dblQQDYAhKwftzeRbJK9GVVKT2gRelMBswATD5cHYHMyX5QacRw6gQ8Zj+NaHtz1MB
HIHyIvBHjSyHaA8MEgGgvYw0mt9FPk2aR+kjiwppTJNLvmqXKNhXm91q3y0tcwGLHzccypYwE4PW
O03FhSVA6zADMQorO6GnAOQA+Vq//a9zV0WqhjUEwpmRCdTb9U0l/eOG6wjMkyZmw1yGynEVkHOC
LaGPPvmBdmzWCphGtSUTp9OqmBMUI+sLE4z45Qm2uyvpfA1vLpFhha6S8U6ouO3ehkhzv/mxpvMR
GHQ0G/lI3k0o8isrFFz7ONZYg/ZDxNvW0RQy8jy4CuVo7oFKMzTAFB8rpcDU3StN9T5bixUq9zkv
7P+4ydrnuLpBQp0uPsfjrtewgkCejUsQ+z0egN4W8R+i9eqDE7dOpC98KaiutEQU7tFQig/TETYo
fgYxQR+z9GmFiY3KN+tbi3uBTiXem8lTYEWIBJwGHSZAY4tVjQUWcjdnbdLg354PSdxIBTkUwKh+
4fI9uLTjyjfg9ZD6xGFXNYR7WG0igdjZqNUpcayL0AgBsHnBA3bj56MMlSPLAEX7hCSiAi4QG7J/
oAW6Uv29IV7E8rB5j4UXBMNkW2fdAJ0wL/3cWC5HGYWMjCGveARAkVftXm+BXuaj6Cf93ORAu7Qw
TBqcEZVTro+3wqw/coM/R76rzUHN/TMl5bQnoqAxdchrz1gieKZ5t/yIAwtUI3akMXnMfGJfau2G
ANxqEafjaOiNzN7pfPt35jN4l1GEJjCFE9yBnRa17gSanTfNGxzG1nNw+BUO4cqEL7JpcbhYYZ2D
7IiQt6Ikx//b2+nnHGhdTg2tvuxNjN0eiaPQsbiTU2DajK8AH13z0UGnD0WITfvodU62KYcctCge
EdepTP/VMjKZBR6+D5q3QDjAoe6KnJ0pr699wdFoNYEnqVSB85qw3mIcg1baTCqo3L3exX0ZmiPm
lm81URyRqIolpCnUkU2T79reKFWZFIknerXxnUhw4ugL+yvmvDn7A69WQkjgc3bG3j89dS3xUpVi
wUdmLiOPUn9hetFiOcbyIq/ewF/AbLwmw89Wh2sfYfb8dVMDJjE0H6uQ/Ouwn3cy6fMuwUpnn2tB
p5Qyfyr/OdQI2tJfXVrlNPx6aL3QkajbVsAqcjdMDmoysZMl1qAJ3YtSaL3za2eqt/7aqjlJ84Xb
nEJYf0bdaCk5U2d74g42nwBeIV5C+tbaC64qA1QTkTzyAwwiAzM/X+pQlWS1yGbZp6eb8rcbXBIS
Bxk86r7fx5D4TWVZmAZaSuB1ulQN/lkO4WNmHilZru67aleXKbKVyVZ4MNZ9GdAHe+WHZU2Jl4Ov
IxciAooV61yLabBEATt13CitAyd3fpZ1FDsO1qlkhBIT9fbydFVVfBLV3BO8lsbpBapaGMOtWRDd
y/CqWsuJqVl+QjFDChdJ2hR673w965yHziFjfXQjs9dlpEp33GSUDrSxwbhrVOBjurIeyQQIFfj8
JVKvkzMdzGIXIjfNoPv2xTN+v9FE+Us+mPtK0qLu0Xki9TIKm7bmXpejDM8gpF4CWel5KrLY9K1p
7a7FnBvukqj56x9ARd9GI3GA0XMo1tnF0JDm9+vi8mlkFeulUk1oRd2i9AC+RzhgWXGqvlg1h9fR
J7xCv3ClCqfQOkHXHc3kJWviSnZHjJBrOPtVy0LwMStoVGKA99t7Uof3n8sHjhKyH0Q50glz3hyW
ljlEyUZqbd8aQVPQK3sp8w+NjJUMPlAbItDF5SYWIZVLQW4K4sVnIRaBPiOhTbK5v2p5VKVAMl4e
E74lkBMl+R9SkUZR3Do4APW6qiymeIymxKCUd6HfCEF2X1WmoYOoXErhqwPMq3m4wAbnG90ih54b
mi3Lz7Nwt5IpJ7bD6RXHbS336jiOWxF0R9t3tQjfFfkPhz8zo1spKsEjjm9rOjKBXIIj+SDmltVp
56tvvuu7KnloaVq7SyGTE+94qtbM2pseFsAhkcw5V9m+LBUkLc4yLL5H0dUwevaoyDe0EgDic2EF
yVKX8GF0DsiJaKrAmuPhrUex/MJxW+JmLNOjBE9xSSQMQVK7zu4qo7jHAjONZLujZmCgtiPYuuxe
cGJp5GtgAg9kT47D4QRNhK94fvnySIwrfHa+XwyPlISDi4STRE/fYh5xKhGRpz+V+XBbqofIE6V7
D9rS0DRm9gL31lBn2rbMIxuOjNmgSJNJr85+Ws/EVDce+LAyG4Ojj/91ZDSlv8AMKL7g82xKHt9G
MotyX3WFtjjnE2xTy8BNKtrweuvQ16SRQnZNTkbEuP2f3bSyNvEIablajNhzSWAL4qxjFsGnnvwg
byXHb0CKeO2NnTMH3vqKuL5K8+rROdUDGjYJ8SfG6pBdzbsC4Ngm1Km7QSDlPg58v4H0pxFfFhkL
B/ApzqdK/k4q/DxdnrGw2uw9/PwfamfZBI3avKt8a5+gKS9DZLaRU3en3Byv4RG6udSZaGvEJ9ip
3cglxJ98ahNtiLPvbCYbiS70KM10S4/UtXr9W3xYuNgDD/xWMmnZTVLuln98vuiM1cwBowq0T/m+
ySkmc6HpBWM9IxHR21r/rXhLFIUHgtGjqh0RUlUNAZTPZlXXKvtFXfTbJy/qUwt0MDc9saHj6FlW
ECfPdwpF94UY1lYd04gEkrd62rQTbfd8G/hSX3Xi2xyeMjvJ25E8nZd+XJXrJcUw4gpQvEPBxr0N
TRxs//62IF9FOL0TuJuspCt55Ly6BZaE3fDaNV8QXixzz+9Fot3KrEjhNPFbDAXB/xJ/2nB5AgW1
aOUdleVheJGwsNu7lFRc23lHn0mOVT4aSg7BThWZ+D7DFha1zmOBSaB+6i2uUsCitskxw65x9cVO
l7mgI7vg8XX0wp6QXlLbX/xS6k20SZCkQ6V8ik9BTDupFMWZo4/4QjFnWQAG4H8CXpL/2eeJ4vWh
dK1X/PrHf0+N+eVE5goWhI44KY/3v6wMdmbQaZtOVnjPkXeyYJbYmtYqHa4GBzFLgocCsqNxPCHa
NoYYuTceztoEXuAlalcgKv4+3TNJBid1r5q66M1B9KWt7dsT23rYqXDvaod6pQ+A9n7uX101UEz6
rqpi6tQM3Z6OhUybaeK0zBKnbEc7GUyUbNBmSc/WtSTHo5D3NbgdUJgddJNHJyYhN8OHVwcbD+Mr
Q/zteXoEMynjSTRoNVexX96jgZoGeHzgCMHePe7MQ5mrRlvikQiUQwuEdK74lfkx/Qr9WFK81ee1
aFyrnnx142Vvz2pAIpHmEI/fFCCIbAbiCLsdMQ75Aq64mJ2cR7HK1T/VVdaqYRDNjQ+B2yznL1ul
O7javjPG2SNtXvGoCBWBY0l0hnJmVYg5mSYfwGFfA4jTVzlAX5S5JsEDAGDCezLyL8UJV0Jn5CSW
P0z0COUUsFWlRik6Y2MbJMWqZOAa/AFNJ6tS8vAljlPJ0OGGbMUCHYT7FhNQbeQ4IAkuiob9NFwP
PtzZ/5BNydpZAKtlTZHfAacBy/Ih1Ukg/3G4K8o3CU38e8n4lw4knxJhcZNtuMvKvzRS1JjGfHwX
2Al0rxdAv5cMG5SDuTqxgEPQGNTzzGxwt0M5+SDQ9OhmeubBgoGbrIqS9+NL1LTEriOSwH5rahMw
iWDSqVepEsd6Wr/8esSvsA55FKQMRSHqQYSFW31245gxW1czzLA4HXARrOTL9Ux30QJSZAgvtCY2
I61Nif5S3qvLv1Q5Q6tcjLy67qqDTPpmkuOirIluug2buyBM9I++NQDZiHqu8KpUP9w7XZ+m8Ak2
2ErNq8mhiqJZKV7KUNT+okm+f2EqV7N4q6RAK4RZnCJgT+rw6obh9NKgYe9hDltFhNsCA3TOyG5M
YzZ70wqCV2QrU87jDe1Vx98ZPzRmxrhUzQVrPRj8YI+2wWEBxJOd1HFDExPEtgXd6KrkNemzK87A
7ZgkIackBfa2wPMWfNWMsu83nicAxWs26za6KEm5ZRYD5kQh3LKb3/WcWZzZ32pe4ec4wY9pYSPJ
Oh/eJYAFW+IMJ9o8WikZyhjnIXRMnkCzgi6Xlc3o4dAgjh3wCfQ3qVryU1LJ+paG4h6ugX49G1Vs
+6liBE+h4bJzEMnhPTSybzst2eBaZROkmhQE+7tMZm5wHOR7oC18t2W6wRrHTs7UGzlgbzu8P5Bc
TurfUtHUJRUuKlaluIXSJFZ0TBaFp0PL69jv9C8r2tkLVKsjyaiM8ii4gLZjga1FnuGCiD7HNqPK
nsxYKG4EHqaWXnUjKU/vujkxQhaJh0vMVVps8MVeQU7+NMBMQHCLG/T2wVEfWA3gL18JtJQoK+3W
RdwKtSdT+uzVN/TaavT1cPw+eFWPp4YOTOf3TpoBywrDdknrrQ6ZJYPz0KDfNCiUnWL/0yjZdqCw
3Z/WJuGGCtkPTxA+1Ax0uwyDGZ7Zol3CDgcbS1FOaKQTcvw3VMyc0l9tRTMD09/VRTJVJWK9lwEF
5xC5xwK8Ygbv1qlkA937miC5dYSK5U2VhVa2ldg/LB6pgzzHvrl5jfktxTT4zm0459qvTgyvgc6E
1Cq+Zj4AUbgxRDZt/3qqktKhbQKh4sqmq1z2+wrYCiz1XDeRlBCk5MVKQxd8VJgPG8JH/RcrL9UG
1pzQZWKg2rR/7+YxOqKY3ukn7/bLLh9NEUHAZKnSNVOAGfCTNeblukxZ90mRkasxbFkqVwz9uZzJ
gpBM5azDDepBMHTyeLQ1HpQ0fDh5vJnvt/U890XHWcPwmBHSgXiArcUFB+fSuk8TezPH5C9UBlLn
CqPJHOpPzkgpfYEG1PsJRt1wm5Ej1BTyLHl5CtE8r9qtbLKKzhFHmn13m3ve/uSVNYEdZP/Kfdpj
iz5Jsws/EuuGxLExA1wRvy+FuHnOWxx63YgYHTQHQhgxBVxI0LwseM0SDifkUvO+3kMUDQHZECP4
B+ZRkhXKv5INVTPcxxx86lYu/mvx2nL/jR2AlYhcNxxNTptUD3DoqfunwImzB2nTugT6CRl7T4VX
6pKzplouBcRzQEQG3X/NrmwxdS0/fpJE2wh820Hm+LDKOnqWycx8PECewqoZ0Ngh866CLlzPsAWn
CvRofRYacR01HfqA5nb7On7dSigG4cknojy0fdbhAkBHAptqFqZ1+8uQw63xA9crE0FgcNgviGLE
V8dcG431XpysAW9LBRoafAT3izP23yI9fWOns0qL37Z4hQqx4K0vPZOjBIp8KEDZXj9nCimm69Yg
j+Uk6G3YrXHCOZvKyWqZTlf+W5b5M1DN/j34wWoW+qS4cUUjbfyjmq2Y8W7eIMCvtKoBBUhjhhGp
Y5srEkfJ96jwMHLZBkQ/7UFEcYMmGOWa0tt/U7UERSoY4dHPBQPrvpebEHVT5zGLeWWAk5pypOGV
SXTbn+xDtCrBfzDkHSYAuQlw+z3dawCCuYk+iLRVK/HBFb7cbWQrkjkUMjyjrRKPN4zI/2z19m4E
c7Zm7bVR0ljD2GdPS5/78VyoBmA88n/WTpnCzCwvuGwZsAQFFgdg8wMO1ahHW5e3CF5gS6wylFj1
9nHGIueVIYgulV4zqGYf22f6u3ZFtKr0W4xep/NEAGD5Nqtm+skOLwSeXdMAVNeyVoYklIpNtzly
cKJ9p5L98urR47MAmucR3+l1etyT3svSh0aotc9e9oF6b9CvifPc1jd69z535MfURffqhLmpgXhU
cFaEZbBhi1sU2GrMpH0XDXQzqwM7f5w2QK1ykT79tXLt3WgM/DDYeLLxhe1AoH1Yza94RKr1oYoO
ZGzZxge5m/LtlLvCh4NJIa+wwTyQugQmwLywbQbyz9hcDLBma2uSTLEnVjdjkVAPqHEvCRaEiftp
2A1AC+1yIluW8j+tfdoaKWZsjXhtnnVYzeA8RqzxKR78iga7Gi0e6h63OmdKFPtxtO6owps7wrfI
chQeZ6lsIT9f3bcAlkeFcwYjAkeIE33vdmHJpIoX9yeQEhKiV7AAHY8T6Tj9qBsiDnBa0Bl+zRhR
aiNkm9E7wTFKHz2gsWpho16RCt9vzd27wOH0g1chxDdIfP1Ids6+70mXuaKFoKIpDUW+oV2OyfKM
IkNJtymBb2nZMzjZOgCL/fvVwT1Hr02goRp9StpC5/c5jtjyZRfN/6JrjiYAtffpFtR3X5iiPOwU
Svm6T9GxczRorIEDczCvQXTUKmWMgs5+vmpmWl0gVPUuwGrgijToZJyPbpDgJxj21cBSriZQcjfP
cEgrxM9CnK1VYqhaK1JaLts8KhcQ9ccP/6VD7ajjc4HRmiuJ1KQ4vDXtQiVLDTm0lkeBH5M0/Aea
//IrlXJUNyq+F+5KxyAFs9sdtyo2oA8eXzgIM3LI/QtwOKxbZYJU1z4GkS67LeNQTnbpxtRIyKZ0
7rMRv6XuMijozC+E9VcMlitculR2G7oPlBMwBkLREonzT6dLL2Ctq2/HAPyXBA39rZ5Vcp0CnC16
55tL0xhaFcWvbJB7uGE4GIcI9AiL0SahUBmGKVwMSAtDPCweZ//oNQXQgJapVCHnwWDn3MziSK6b
DaurZxws9pqYMQalb++mDNI3a/6yp/gy/KsXQVxhapvH0i1TPZK1AiNPFMi3WJ5kcYTQxLnJ5kpL
jWbysdF87njuDa7ezltzOIjbJrmueACLrHOHf6xRcVgPTfXZy9hrSr5TAwiEiviTyHsMqsVfrsqO
cfdqMWZnQA6e1QtcUSx86ymZ1kvdOv1A876TRM5qOlst5UAweZieQL4FrNJXdTcRWiWTNOoGcQtF
yGmjcaToSZFwNWifUQS3RlICnwu9+bfU6OSJhKgZdk1ozP5TwFOKVdD8AjB6DYrvB4mWeNoGr0/f
0jKZfI9GTFnqs5/Q4+GBsduMBIG3RHIQ797yhEJ5lzMVT5AoWQ3aBPBwSQ+gwLStYK8eQLmwVFTM
KVY1ewbYyK8plnfBaIxPPPEUMpvXhBuCrXGoCJc0WEfXsMfa06xer2V31OoFTpVX9Ub7Qt7/VVkA
EliLDlf810VNG7lh527UQhQKfXHqkeQzy9zS1UFiprconyIEhir326NsqAxi0SjzpQhFWwhoadqX
MWJ3egmE2MJcUvtvPNO04eZsbi1zKhYR1XFpiae0qqfHHELVx2qlvAezYcODgvT9hI+C2V8Uu9qG
qV5gwr7RlU+T5f8Kn/Pj+TMydUOqpZtcVpPcOY2V/t09Y69lfiPOM5c9dMSQfSUiTAWvxZdHQzRP
Tr05en1B8F2fo5qyXm6VtiXybc+2A3t07sc/gQamYW6KhvdhY8Gp31fv/FvFHlcOf9tybwxDbMS2
BU+vFjl39xhVs7v7Uv5Y7cTQlWxC+yIiSWUs8Hg1H6a4oIgYNZy1RHMbeAY0tYrE8Cbs+YQaP35X
DDaQBzkVXy1+qk9Ypxp2wXfQv+t9Sd0l4GFjP+NVsy04Tzda4TW1CuD5Qwbpl8F1Mwi3E1mVk4nI
nbtbCTL/dnXFQCkYyV2qVqYnv4VQi+RmRAsGJ88j+L/nnySZhAcaN4UrGmMYAXm9on5ZFFymdXtC
Ga6jSFiRljX7OdD8YQPJsnt095kWFUaPpaJHmdrFnkFPvwJvosW8yZxNAwplq8b7ssqmU7O1x96z
QX4Hw3AnycmplpWycZH9kdiR9kFH3h+UtvuuKMG7wcGauso9LAEsoVs7SSEqEowWuQvnZeoGW+40
p1ljahRrv971SHtzxoXjnaXMRdb7ABNc6XJGAmkzfUQ3JtJ8KAO/xy64FbahLDgLr5IdTRCVAXRC
3Vhf18uBox+lki9EbsvKODgOnBtjADt1ZxziNZh9nslsNfZtPS4ZvYXcb4VkpJyJWYbBYwye72HA
R9qph3uvJCewfX5GDo8MceVpA43YcUUk9TqihNU2HBJIIcsXVMZIHAMS1INbPQTfJgtszdQn5vh9
DgBq6c78STV/p1eP9WToRySlfTjkp9KeLicrPL3duKcDDsAXLSGvYEvO2yJ4UFP3RfpZnmCeMqA5
SBfINhSLB50g73jsYvyy3fduRO82YkvEZ4lLOQfVJswJ2Ci1+DUhOLfSeJiCxInZsjpu6Ba77Tt9
r6bnSVUHN4yhih38Z0Vop0UZ55/tra4LwXMARJHMc4ucd609OmHfbN4P1QDqwz/4wUSxeCjpHVlh
UTJFbsaUcXIguC/nJAYULqWKsc6qaBWWpV5t9Bpeb+lmtTVBGIlEGJQiQwCXC6rKglYbvPurlXt9
z4ahYehoI98b/3KkEAWjjBvY9c5umvrW2PArGV6zpvbetmyoWni+6QkGvHYxe0FRG+pmcnFPUuMf
xIckVKgFHkI1yqgaWLe+nk3D4gVrgkujkGk4Y+E3QwkErDv2RULohM74bA5EBGbENIGS+rm8suu5
u8NERH5Ewzx3f9DDbl7427F+uUMSPQG/bl6nqR3fbe5cWRwvJTVEiW2o3N5gLcBh5xy3WbB18xlT
gD+s5vehn3wC+anGLbiVV51JnBWIS5W58Cnh+1LT4IxzIyPXDxGlxhKrEMmUw7XxN26mJwiRhar1
qu9r9zcMTMZHOwzvN1Bli6wLm1ulrBkUEfne08KPQMZl3MX/zV0AQBDElnwJglzdSLa/AbUYfgId
PItSjCh8DDCnkzpSP2fsRa87gCaGQbD46d2JlWz80vRfvi2Jm9DcyrFbXp+YQJqxEVBjlseM2019
nZrQvaDX4/+JrwXPtBfZuHh/qKjBUI3hQ9Y62PspL8z9pF+quNkdPHG7dKhwWGVmX7fqoP7RXQuG
4oE9phuXE4yOtC+rDYJvwGK/zt0oUvC+uK1OE01/D5iRZN16KwEqbGdvFIcEqGrh3ObSBuenMQq+
/IGecuE1jYUFh/aVWUoei0cyev2F+551mFBKYBJVjFAngbETrK0uhEC1fzmxRcxOn4nqvYHen2fM
TUpC0kEYD4QNpwltem/yDk2esMh47fMpSvE443CCyiPmtUe5mqB1zq29uwu2w+x/yNak5rP5ju0F
JKln/nyThBWGo4G7SSQ54GmYWT9q9J+6j0wSTQRjx2H4cbQbEOkKz1mrqVcI24Yu5ucBro2yvpr/
DLid2vUXz5zQv7QvGDOQ0ppFGCW9qqbkfkot2e34afS4VZepqq53yuJUQMZYPVACcaHrqzTPt09Q
7CxOzIW8tqYM3OvcR0GOe6AsZXu59rrBEJIAOEoCBmnTc1I5ZW9kbqc2H3+CIHnaPHUZIt6URJoc
xjJlhhytGeFfCwMEoZesUZBSLx3z704J8YGkId6nZLcOMsBYWkRKVGK2RtSJR9OgbTj5y5WNTomV
NT5WO/losyAlFvqpMZPr3wCCblDjPlQYH/3BGNcc0RTZHlfRnPzlKrTS+EP2oFs9OEnxwzR9Urtl
vVxibhGwxqsgS48xFFGsEMZI16lq4chw6Q/qBg1NJ1Ff0ByL0D1Rl/ln6S8Nu7rJvuf4zDcI7wz9
oGJLTybdPdvoH5iYuKu5rX7i/bCtZBAA3TIBLCL99QIIM+PT+bkQeSk9n4TGu2dvxrITV1W6V4uM
8/irX8SzBf4T1cPIOi3zm3jrlIcXVVawoWPTEIi10/V9dU6GncRzjUkINdfAK8fzqRPisZ5AWtng
o8fFxAWjghh9DGeFVe7mNy/lvy79vEBhOQn4BRi6D+bULsZ8AoQTSTJQx2FAJFRWrhST/78fGXZj
PyaZW6eU8jKTzCi2QJ7TE+9DB4jP2zIOseunXT/ta7xqrbQK3zw3ZRDQscl+tYOlzUSVzkySe+hS
8Qltl4MGxXcSGTSBJRx5jS/GQmGhXkFVJsdgyJqLYmAkejApMXRrRIB3ttEQcTMDMc1e8bObv5HN
uPDECV4Ge6dBh0pt15VETpyKXuyVybScNZYvbW3JZNVZZ0JyGUJljtA6NCzl9ltE1cxHwnYEilSG
rlZusPO0Aj4njcO8KZrrA2wX40/nZCYcNXPmQ8kJmnATmW87CqJ/u1EQcDhTsjYjDMpbLjFJWjiK
t3pU9v6ukrI9XiiXMvDY+aw3WkBhOKDlvVhMTe7jwXfPJnr1Y0idkCZEcu129fSCIpREYQjvfiAs
oppfxjpwbjsnVLJIc5mPkObeDPr88f6ZLtJYFH097TRo7XojATOM+6Thtdxfgw+rO9N4V7U6fzeC
dkYyx0DI+0lnSnU572Dm8wUrfuZDg25NQpxLVsdy4hbr0Y+x0Y05VlRzb1Es04IybBylys4pNzuq
9lAy8JwShAifdO/dEqttBfKBFC56dLV8WcHT5u7zOSAiUg1rba37EPwJTbr9zj0xQ9Wy0e+fXg26
aXfise/BFeQ4dBQT/qtk3kbOnpK4F0cICntSw5LaGDJYOQpDMH4r3kaj/2CZqrkpk2YQbDIwv6eK
yxwzvXtoZzbNWSnFC2BiS3w4DSL+6YkdumMRo0q33EUrvwAaceFat5Mz9/hkip6pBu0Dhb8L/Dix
WW/lJxCa2JPUQJgZDzDrZX5SKA77DDAgmgYJw/hoP4RiiUrdl0Bt18xV55i/Bz+R9TMLSv3CufhK
igQNdX+ZQ903FjlfEVjXURg6eFExsWazG1ZhE71yFJNJRnq7NA3EPlKbZb58BQCp3nDsep7d2Kgc
sgnJVDDSgvtiwOu9oVc1GtrYVwFo6tpiQu0loU8FE2twUaL4rViS+q6uEscUpXTEXkFkHunVHyOU
RXJv1gNAF613vZgiLFKODV9mDDGo0wMtajzPkqRV1QCuqXaoj92YjMkls4CJVsz5zmttmfcVXX1S
hLkDzPznqW0YWfJJbzslcelT625bniIo4wstTIh5nZ7vJjjN6l3wGUIs7bHqShPkw9d0Er8EXVME
3FfkG2TC8OYW6qmOk4ttXptJNzbloPKrzMYcFyeKXPSQBL3kuy9eNfbqIv1GX6AnZnK2ko1Optrb
ILZlECpXQHLQ5Zma9Dvoz9W8Ha1h0mihBOasQoPzip1kodiThc/z6Y0neBsz6Bm0FcgMzV/kKfCy
MlyT8mp7jZubdZVqbfwTpfzzf03mAPTSWUenlAbMfLvimoJ1QddZcZ4PrbRRmkYS3+9wNTfu3yP5
blQ6csW5+bIROvnkUM1hrObrhJeD71sG9e8+ppqCNjOUXYqOjAJvBOKpYMX3/Oz3/sUO6VWeSI5Y
wtut7sBr8gtEDrZ9spIBPV7ZHUou26Y3R7XpK0fz9xHv6NL1A0uEQ8JpXfqplz9LzRrnnvEqtPzR
A9D2tucW4OlxhfRrwiSaJz3K94dcP+hepK/nd+nSin9GLr/vI8XRcpXRr3ktsboUhtjX6UhkxQn7
FcvTHEvol/lssyNU4XOSKa5dmxIiL5tk9UfJTDRO2z698eb+HmNZVjKuCPkFErQ03bcdIGEsYStA
3wRDx7hlfhcoKHmev5b5Ut0g7MrKpUEq0Fljpz1L7W+/PZqDktvIC2K3W7lkQ78M0/rSaZ7X3C6e
cOCgFAJBqXgYTJiT5YFAbFQ/OD55r1VjWUAg/rBeEaOqrYMgBLrLaJ5BJ91ZGDzNTvWB3i9Rc8Sf
mjFm+58cIgvr6RnrZPYFVcfyhhIBuJdrltQmb4OX2KZ7fO4BNPdb8HTzQ4NmDR4Evi+pk5ZVNcMg
FsqHmYNGBqnXFk2raxUxpn/DvmydJaXJRDKFlbRu8I8EyLPn1sYpI5Wpib+FjMQLaYlcBPuJRf7C
1sedGEP6suMje6BTf4pP2Oo5r79GolvAIYq4GVEk88QGWof8LYjYRhfIqmRCdES2jIsY2gWOn+nj
rQaYX4/Lk5iEevMhVJghA4lI0B5nvf7qvemUpJJFjaXyahgW0gE/BFk7W72148N2waJpvlxeiJzO
+A9iDjx0IeaeCe9tFi6D+c//fnWeJ6gAjynsdlPOTvslLn3kbDFB5Pnom9AgGcaj6dmHGpAsKYqc
1FKypJadZ7xJ02/9EB1nO6jGCeW812wsbyEZQojpGl+q2a6bOH8mqbYTAg0LMHv94MKHv2pCUp9h
4bygy065OV6ttUOpR0ljMhK4dIjoXcZagi+LbNZOrQhjJiPc4ls4sQSECbZKBce6gvst2UNxUa8Z
sGXtDR6vuxi7CToQVdwJAS6F9SPy7cXP9Hm2bzI6UvHQAE0w6DUhhqr+dEQOr7YvcikSSr8wq/xB
haJrCVmHQBcfERPhwvxBWbxctpb3AWb75qHFxZgz3YT6UPchGNNFGwaO6kHmBsOoIzPY2VbK9/kr
AUgaQc6DzlYOLG5hBWuPiCLsSBYlg9Z83oQtFHw2bV9vCNYH/JYWgee9d2ToLjAvGI1ta7iKOro5
44jgmFufkz4eU2HmVBp8lUhwuREnMF3adaIijFNVRHPpRphLjUGj26XdxZLHLf+NowGm5xWDeOs4
QCL2hlgzkBJI631aWPv6ZzEjU4K9nPkV6GXFQa4C//pZPYv3SuKeHcfzLhwD8UkQBvDPt23ezFfW
TtDJGJC7WqkW4aXZpSh1ofSTBgT8LtY3xNf9ebd8rLAIk4RCSvrmSyy6dt65bHLoVTapxyNQ+93X
sn5EyOtjfRUVa3zUfNORaSPhCzUAgh/CpzEtMg9P3xBaeUta29ocdUXoiJt8FubZgDKgRDYFVChY
bupRnyw6VPb9sIYM7XiT/n3e/UNaG59L1Y5yCmVbulkA0jjYGD7vKx4fXfDBsWXkFsh53OJvSX+D
5q0qrQjNdyOkVIZ0WnG1YBf2zg7kuIg+qbbVIEmhEa9Rrwiq60HPdIozEVJX0hvxglHJfn7pKsnd
xrq6ZByuTYZzV7NHoFyz51wn/VMXIejm593dZ8xUq/ca/qUvk8xK3aVvNt9L8qkVQEMWcB9U1Ud5
7s+D5Q9YWrq1/nYKbfJqWJ+zvt5mX5wMxsZQruWQkhqf75j+gfcmsg2VxTTGyEPX6XUXu8Lk+IJw
yNLRMOQUzF2oJr7ND4GHsKIDz/jlTjozD+NztzN6WF6TpzLAO09rmSjUBEOIZ/FSQ+8iXTPVWF8I
kmOGZ8YckDvtmbb3hJ1b4c6Gq2+z59MHfv2YObS/BumiZkna/pL22XxRtt17YzAd8Vv71PU4rTrO
d69SoZgDw4jgYmC7fh8x4Q0TdNS1MoIrM9IKjk2JsxDiyorJdGtVpYHVuiSJDrxnl/T0TmcVuefl
pVfjiqi5Ov0d7QtmEvqir+3kNLaJrfG2JSWcqQcVWSiBlsAt7tidPGbUUJ8kBLYPF9r+4IYml754
PWvEHCzP4Utq9dzKThfwx6YzYWzbOUPHHCd6wUeqn6JoQYRRrRh9pvQDE+WkJbpYh/HAaUp9cB60
K5BOVwZlXRxGHlzMB9DUwPhYiTgONzucc39EepPgllYGolxv8WT1UEM1wcGO3ZfyMucv2XAREUME
qw45YEdrvogR6x+2VPpbttwaXqEj7y/bWp2bVLnV9CIsyTzz3N3wZ0i+GUcJHFxA9UrRv3lpOB71
4ohYe7SwdpnrrnSlzua69qD9U0pLykCSTCLLCYYW2tNcuRcoNFZkcLjBPG2WgBQLNiqoBb+5ewTF
fbIO/I99bwXt4qX07la3vmXGmeN5hk9GW/b/zdzqN6QoImELFMmmqARyonZo3tt8M28KAHOWK4gc
uFgrViaG2ZruxN/HGXmDxaRPg7QISiRYjLEZ2loJ5w0LCJNHFQX+WBR8EFMOzIIeS/ZE6tDYQGaG
WvH04fUXf4gd0sE28pmoKHpnYUC4i87YI28qSreWiTt1AHXwcYvk047do2pwaFCfK9J8XzYzgZ5H
bCRRmmwFsUjbEoaPP5wsPDdYgWpwlf7d2BxjgrZjlkShX9rKrce/HNTfymezLw9F3EyOGdduXoOa
KJyTZNuWRrlb1mkEPvPr2ZZV6gwVASCYPPPoZYIJhp0B+Jxnx4AERlZ0g93VNYlf84A6SFkzXZzB
2xsqUIx+viijbKN7Zb76VOTMVGcSLr3mMQ4akMefQCrQ+x6gOJ2ciRGzPaIc0UyGxN85+V38lMhw
TSWH+8Z7ZIidfH7UBg3MHRqhPkyJx5CvYhwheBoieJYb9ksx3hSHZNVVK/XbQQDkQfpKooDGAkuH
HV+n2QYpJS3vrVXR6b3fgVwB0+9xfqoLqicmD74odzDZsS4n4BJcqK4xm1oVjBUovGHsO2AM143D
aLwMxTdnQR6YDLH44UL55qpgz2QGHEV8nKLQ1UU+VonM1L5jue/PUasqW+uETwpG0d+7RO9fxiPy
dS7dsFWAIEH4BUXCAwANGFzxYeAXpQphYCaEu3D+DIQyhB+3nZJRFIaTDsngt0JcXCOu0jzSY4Di
WAz1Q6meosRFlBjJeTn8JciPj0UdG8PGevvrRSbzrS3TGK6KYx2j/64CIVoHAQjF/hRd8bKtAOzx
pJQJupB+KX6RTvVzUztuVpSRzW0vexVQ9kNKzIENLHV3g77kbyA8KTL5gb4ySXkpjbGcDhRg2cTa
OOG5MJ36y8s4D+LBm0xjCDjVQsyTLkhg2+HrKIGq8K2jUpfEFXWJZxDdCBN+OT+eZSm3MQ4KV2R3
Jveb/9kyK9Emkbml4pGHRz/n+NfI/SK6A/9mt5zRhUNGFWBP1QEIDpl4Kjqc9qLVJGVlphjjBtvu
7T4711IjDnVi//moT26m9jHUfPvIepZ0lCMP3jPCkY66crfRywZEwBZgsGJ6C2b4VstspuP6AeFn
/iOTxeMezpj8NdA08Cwal2V5rYe6suq/+n47jx1HBOyUzhC3s6Pf8j11E44NEC0C09ddt4LP4JIc
jEy5xje0aALpswlTgidUU9c6/AMGVPap0l2b0RRPJ73zq4K9CmXiN98oqrDmco1eSBYJAc5UNxdf
Unmr0ZxBuDw0Iij5rmZvSqXz0PSQmok4EmM1avpcG8pi7GaZgC9HkLYpbYxxPHSP8kpYDSbqsHa0
ff9c2cmyOetmtbGARED4y8BCi5/PBEzd0kMqItHUfLWx6zJdTWrBX46EfLwuHCkH0l986CmgxGCm
q3hZhQftiw/vys5MUDUjHr4UW3j1XnaTLUqhVb3+asfXpYZp9Hc+UzNB0FZRNtTt9olrk8MckX9r
K3J21TJ67nV+q+OlutIHUBXeV48t5/stUi+irGChrBQp0r3sbQjqMyaN59p02+eGvW8pEseBQyLP
DIqFgEvIHexittamuOFueRcmBJuZ3dz1DjqrD1JYSSob6o251KUnMXIb3ynI3VJD9gxZ9GY8CtE0
M8fwg/PCttKPEDTX3YTfSGhfTONNBUSHuvBVkOyjHoYmFQs7tiWd0AonvnTnNkF6L1nGn7I8MOhS
tCcntY7c1s9sfsXBSqBbVH9mC1+HgVPF9UY2sQDsJkikklvHtqGNd/SywWZFKAIC/Xd1tmb8sOho
a1DGRTMim/y2++8JhwIxnMDQaLyYAzIpKxD8baCfbIlOjMwEJq3prwyj1paLcJVEcTkM3LdKoqjB
pNjD+IRknC6/y69HnB3fC/eL2qom9m4z2yjeFZx20qJolWVKuMmV9kkXgPJSXIdSTZPxfu2mYVE5
mF49InbEhN+6Qtq4rNTeS4fCpU4yYRCLkxmxSP7SYogPVKOncZ4z46GXoR2KmW4lIobiCHgqxtBi
Uluf83hjTGy4EHOFAVrlw+y4hKmgnzfiMTYY7Fu/8rwqA1MlENIcE6oUGgFblcl2f+DjyljPBJre
nFXk5pt+iKbwwpIAHuVB+At6mX9yycRT3KPlRg0o9DYRENgihPzHrIdhYOocOmd9EM3AYptg8wVt
PQpqm//KkcyW47sdcV2tV1lnYu8rXWeS1nUI8eUVC5jM6envdo6jLeCJRYMOG7CIw4O33aPT59TD
FRsaB0lXj/o5zzIFDmWiTesVNiwAIpBf9TPskBgT8nfQJsYM7mBomA+6X0cHlUfAZ59Ex/hT8SDP
OfDMC44gES9IVHbdbnubYAOke+LTf6o87NY40MyfhrJ7Vfmpbt9tvKrg8Hcbn9RS1W7rNY4SqOUm
CGKJkmSO6U1FHgyl58TSqj8SnzZGyWlp2VDkVzM6+NbYg6dG6yci56D4avMYE/n1X5U7QUWJjaVm
7Rh03QYgnX90oltrZzhKBHkXLKZHlgmdONxNYLGw8fQemFcEjBdp/3Qc+sl4hOqq+blVYx6VjOlm
+3nAosqUDydBxM+8Nmv17TrW2sz8cKDUoyH88BehxHaEwh371+ZfVOPI2O5BfBhKpnQfacMHbPte
iQlU0Ej+uWIogG6jp4yxMmLFZlehDds7ZhF3knj+RBBDDv3ZhgTTvm2xK45U/LtiUZJeRkgLQ/Hs
uPQjSu6eA08hpkmllY++SUJKrfNmq/I/X4X1KqDWst9trKBp1jPtgS7V2PtWVoALbANnLZSPySNI
ycSmwojxgw6G4f1rmIQ3hBVfBWuRq1xbsEUOZ8+bkW96kOlloJdzXTAFaA69SWrZpqppy0BX6uq/
odl9dD474wDQbH/zfthcTXQijxnxFZXmBbyajkgi0XQi1XjbPKhGg9tL6rvdRpciHfOhY4nzxCmg
DCq88B7naS1hcxYoRSVYc/tzvjK/fDfbLYUW3aVeKy03Nu3isn17C7OWipD5TuGAD8rsgMY3yxG0
jAfUFrAytzVJJzGS0NgJkhDb31eiBQVd8aym1wkF/YMS6XvZzqcVtyCIuaOeva6Xq2SZ3AVlBujk
kIivA5RKWZe48VVNE5HLXNrGBjmG/fjryLHWbVObqakhVzVKcJQm8EN0SCBzCUfJphnmb+ikXjs1
XdVDLi3mVUaopE9Euk3dimR+kJkmd7VunHnZwKM9tjCzR0RuvRR0LmrIaSh/HBtd4kFbeKJPRcbo
Ckem7mFolLYeddZvbCyq3tC3ZPE3+o+BSFwrAU8hDFoHM5kBxF8vsICLwmoOaxL1Z8Z3Q9ab2WHn
ftruXpQKCVZ6vAHOH9tPmhwGku+B86BiAx6lX5Yp4QkV1p6XUnfayd6nNYie0vsbXnGYRFNdNcBG
MimCJ3afOcSiRiPHzIGL1TCntgNxucc1VGEi/tJdKJ3rsxuCm5Rf1sIYXPd08kfzWeisHBbhn1+x
1XgXJBtxaiOgEuQ3sq12p1o5toH4Jv4O9d5GfXrrUABJaeJhBaczILJR03dInSLy9vqMeWEjYUbo
WlHrWQqAp8hqFuCr2uG2T9aaTlJGZhmuV7G7BMaleB6CwU5FPlcEQUln3LSb+WAZ9j1+8w/4GsxL
oCuqXSs4CLLF3mBjG0MIxjTMSgVkLl8x4FV4g920ab7oe2umZEmzhW3pKFb21TTLxmbeIWXPCGNf
wMR57mJT7cEjsaKhiU/JbUGglfty0SpkZcCSSSrpo47NI/bGZehDdfbmtSPxLczmX3lzmSoSjsV5
21sAuf1Yw9sQp4maqDJsjzvf4XkV8ahM08t84Ga9b7DJkuSFookOgRqgoZKapMd3PYONgIREU1dQ
2ugjEzg/OgTTmsKV0DpEQcyMvimoVQi+jVkmTwg4rKdbjyk551mHrw/Y7CBQUdZElBeAB88phJKy
/69hbf66Y5FWb/lx0/+kyfMinz7MOBYlb6Mb7mlidDRot5Bj6Un+P7BiGr2SVfhy9CdO2pqGTGiW
2yFWViWkLPvaS+BCL1dyedF6R/S3d0+MxisRtTE0Pc73zTHDMhYR9GSSe/RGQk/5avCKYJqtqX9r
7Gvd3c/neMpHl34OhyVIqkRnsSW9CUxYvk4I8hhK5GtmO9soK7JuPCMkF6cyMYizhZayfAwN5PUu
Zb479iI4UtXkVDMgmRp2gBOpbx7WxHLGAAIvUu2erqqombAtKKaCNZ9BniBcr2tTaZP02mwfoKHB
C8LJ9gOcuvS9rO0uOS79SSuu6daxuvUE5MVDB61TIA65W65zuemK8ja8a0kMwviJoDinJyw1QUA1
NoM4q0HHDF2NSt1jd0L8uhX5BjsUg6ABTe3+ObeU13iAq8tBmfpKFcEwxjTv4Gm3e0vjMNfK5H4r
tjvggqLh4/m5Q8HTh3e9Um5JMy1TNKmEpocp1vuAP1PeuxZlWUktPjnm6xpEt6FmDGoZ9+uXZfuO
JUwjOlQh4QUOhSAtOb/frb+H2MikAvzwrtwNXpjIqzCY/EzQAj16BcvAVAusaQ/qfD9gKM8hBY3v
QLUm3WW5iL3JAlJD07kYB0RZ2t6R9w5Equ5Zbdr+WA7X0MqHnhXIesonPTHyt+wpZFoZU7kjEUnb
fBzm5OfP8mqazMwe/GC1aPh7QmHI+NU5DR0RORyVcV/F18EJR+x1mg3cpArStZoAVikNXH0EzVdY
HqXjZ03nfXwCv7+RMn84TDdwUgYNHFsr6/XDiLVeApZTGS3q5xgP6E3RxIvrqzogTEltnkMiQTtT
w0reXpJA6Vr3dMszRqEbuqyu0jCTnxK8IoOx/AlwtgUXpDYd9pplhBJje/YuNLOVSISBc1yfe4Jw
bTCkW3xh2K2mXiBbG6LnevtdLeR7li9fBV6ox5Itsqk1KDzEoSd4GM1/gNLFrLXuHFxkDlpABjJ7
rwKkWuj0oWcwltcBld0pNGoRJXjLGla8oWw9mFnrGDVyd3978MbaBSk9esVdQydiPqGoAXw8Eh9A
US9LMvcT40MOYgxC6O095yUxcsvDjYWivPWOIoYBXqaBgtdZGFC1mtiftFf9h8VvwMHerqVRgqEC
zyJlwPZf7vU3fboPhovPGFk/CqgLuv+EG570GL/egzUWV+mwPH4UOtb/rhC2nK0y4Y5x2aM+x3cQ
CAYcctlub0NuI3m3K6VI8H8PFIVLH5X7ED6O11NwVXYi01/trwtYmjCmZ5CQEzA+1BR65mOjTgUL
TCxsihHjiNLsK/uPMW5aTTqh+Mi85GfOO6ksiRrEO26sptwvW5jbzC73ngsW2J43IgGt/jJMCPq1
ArCdfE7INJxkNNYbCmIV+ZfNuMyWMlR4RATtgkTNc9MhOBtOu9S2fWM929oaaI1irO87KUmCiP4V
z/I/D43VlnB08rNoKg4BD3MUBfWkIzLs3dCOP2Q3HxAlS6qz6IT+bLRBhPlld4Ur6jDLuXRPXR2j
UDFM06JOn4w0xtpY4EwehB7/xBUtVRaf+pA8K+Nk99r3Ccgj0cOTOpFE+6Qd5cscgdv0abE/NWM/
DZd8i1mOAQZhmWaC2YeuXg/TfJRWWwzs9qdf3te8Oc4GWO3j1d0iWPJP5b32RHDImpnjnCLsIqOp
gGxR3YIUGPtVcFKW0YfDfkvDd6pZ3AhCjtsXSy2L1wXNj4CQoKSqI7Pg+S5OixlF0yqvEGlumtu9
Tjd5Cd5Tbst5CZ4P8xczP4F0GpaMgjWzICEWdpZzfmB3v2R4WwdCsneDiDEcTSbNNKJET18m7GmJ
ZsciwhExV7qrymzL+AHTryHloBXojn7q4evBbY3W9eSqBfELA2rW8P4HW4DAmAXsXEqZKoDmVOSv
ynyMvtLIXD0gBcMVPBB8skCbo3X94lrYAC3sVTtdusQEK2Pa3TkSfH+mZoK2nbEExfJrvMZ+eXiM
W6YJGe2gqmK1XMxOS2jl8gJMd57svZEIj0k76mlhXJQJpWpWfXAgxwROzHb422pNi4jJ9vDGZ6AE
lN9/dz1dpwlM7ZH/j4WekuGJnEFnz5vCmXDO+UlE4SjcqAIwn3lq5owHFmMAXWHN8PodJnXe70QU
AejWcQRd/QnwhRvKbxODdL9E42zYj9kMD3HtW7dAZf2ZdBLjB5Rwl/PresubP+2LhF0oY8rrar/0
bzc4rxrccITxipnHAF2w7qDtig0XklagmA/tBH+2JsU1zFzBYGu5D3fgxIZG5YYLcKel/lsZwvxq
qtcowr699oFWyISpS9U+v7lhZAfEmDInixParGkIoRCf3uIy8FpLumotq0J5QQw2ObIyAd3JkoSF
3njI1DINwZleyib81CxbbBgA8MsDiJ8o2RHVFntOeUsvyyxYIFZW0uh9zkBgHmDg9jcWbhRXs0qF
xbvtTwpGa8uJ81tHL9DwlMXsehbllC01JNcfE5XlUOOyHpogdGOn0efzlnTLRh0mFbMHJmB2KsUQ
4VTuVLK2QnOALRuAo7vvJfGzdvZCbuiQeGTrq7Hkz6EnkeYNqFpdR0bO73BvDfsxPWLUL2OvQWlJ
e4zbOAck+j3ELR0AVBqbFFAsqQJOF9x0EIxS/1Tg7zkhf18cD+8ZMyLUC5v8hQo812e+F9DHfik/
Q1k0QPsx4YnIWcoCDtECckG6ci+Ky3ga8ZoDnDgBrvHMg/+SQJ2k5Uhmv7Vp0ZQa4u2TZTxoNaNm
tzkPx/tVwyek98RDiIj5IjwhPPK2PZsnmpPPPnBhiCWzT2Ca6TfLtpMxBlgFAryejZxOV1sAN8TN
mOLiGYbFXb7vcyusz925RbRw7Md8rwK5qNOE28ra9or7mTjCR/k2FzeMEOKWi2IclR5fzIjWS1oM
0glq+h3ZmOeygp/eMZ3/idoFUCtg4DYp1hML5LdP5PWIXXqIkiJHHb08H7vJO866t+rcHDEbwPfm
KsS3l3SNQ6iV15yrWfUsl0TkInB1Q8YfZEOcrr949NMjV3bBVrc8/GRWZ/teZs72AJVjJf8wVAx8
hmn4EcFLIRonwmg2lqNGHNYmSy9Fj3q2lgoA2IQj7tNXKUkXx29O42Y8Ecn4DeEs7f9G3Ina/KHe
E3EPovpBb7eMqe88V67hf+e6KwpWr8W4L2CbOkf3X2VYpsmnyPhJtcDpMJsb/DwRlxlpl5Mu4SpN
B+6WPVtj7F3uyfWAY1uJCpOEokJM8ZzH0yfmOo44RIZwFmC6js6dmmXNas92JJJNVbK0o+RKt3sg
jG645RJAyQCM/0+Vf7RmPBDWj8IvUyBxi9AAmpvHEBwc7UE+Cnj8Nh5fdDr+Kj+Jn+9YiINmSgKT
C8OHIvmUeXOQc8QY75hReH6rMNGFPztkFFngcfjW8YXV3jpMaX+70bOLW1Axhsfwy8muVUBdkxsq
NRqNN9M3mbVFdoWqPG1o7RznbP08LKrmLN8fq+N9UnoGNazOZgtTduegttJGh8Rlhves0oARW02F
BiCTSmazzKU7o+FufxzZG2IHwA/6p2kbLwm0pjjZk4jRIvc64DVQ5IEY7lWto67C4H4CJ8SmY0u0
+6HbrUn26x7tuc5zKxsReWN3dI+e+yDRURV2nT2StZVITY0VYbtu05wWkd8lSCbHzp3JTKgIaNfC
4n0+OhL+II5s1y9yIAGfcFxp8WrV8RDlneAATJY8q2D/TMMD8sBRrn4buszSai+w/k32/B6nLIVI
C+dTru5kVhlzXRqoY5qdfuUsOQHvPfxw6FZc7CNG+oL62xnNVJ8/HlV1uS0vpJ6XftOmPWFIWtHB
1wzZo6ofAr2AOl7KVw35ZDTVzCphv6loKYpM2YqkUnGoJo8veL4aygXdfEwHiGlgwMdxVfXpM6bo
8d0lyHd1hTlMDt3+E8tTPsoZA7OWFIZ8byXIIwji3Kidl+Onz3EgZoXm1vn/caiRxYQFR090XQNj
oRe2uIkL2LaXBjW3YlFxrGldRStHZVxZ0uh3kpR4Uwg/YNoxre8hAYS7bMm51SzFxOw5e1fZowfc
BoZqBaA4mz/bGRSJvZrr8yyP0dL+Hg7mBF9qvDhRn5ltVn9ShFJ7BlDzviD4cDuT82wP8qZRqB0n
TK5fmuBuxpdd/HkPwmI+5QlzCYMpxFlzJoX0kjbisX6BYE5AUEFd6NZZI8SVnsPMAVvi0DOpTADj
8DN3tmtJ9UDmmCHcOQ0vKKIwncucP7fLATex09uRI9V0vYmvlXsUyLI1PqRu6GI8btRnML14f7uD
TJTfD8Z0sltN0Ou6E5Pi/5KPRkroeQmkzOc/sDZIUaHAbbE6V8/QpjEiDTwfYyfdxzO0d0OgsWN7
jT64dNM2zNGgloLwc5m0oGqCaqDrnNDWTuUoIqSAdhokQsULSc34p4xdKTf1ykfiM47E3GPPbXIZ
QbooE6ZNCS1FGsgWnnzGuM46XZe6oO/+HyB/xc3BbnQoojstNRAqoy/rMn3JpQFOR16mv7aeYRZp
ZNvfIxCTqYnPY3i/eORMOjKcSkl9Y27EuBu3TFXHLZKlnv9E7IPn7zq5n4y1IIBErsqhQNeIeKah
VJygDV7Glouq0091NfV71gScaddGa1tdHgn6hOFEvH+Yvn5dHhEsglIFcm5O7VczZVT8UQjCarW6
5Ent5eJodqrarXulTrqmP3Oskzt16QXTnCz6BmZXvOzYBYmsOySYxXy1xYHU3r5bmkE2jFrH4ghS
tLPPUuvwDIfI54o9olwcFSD7cniHv9RoSZoUrHOnQxmh8LeTS9to/4VkGN016AmKDPtRtqPD7Dt+
KVL5rpD/pBQ4jG3fjIWUXDsdpdDVQiCGxuj233vHpmXtEIlSxjBYGEjrKQFzVZhT/0m/G7bEWKvQ
9XEXIckg5goXrNgEVYB/5hSJlCswHT2a8fWEiiCAyiexwNIf1fTxTUGFesL+hZfGx8+iCmFoK3zz
+8EZKJBTjeHc2evR9b3X95kAcHSivsn8zzjBd3fXkqkveM4CrE/cxC4uWplG0PUMEAmwKJWVnxop
WU/lrr5GU0RtVcUjPXUeyDWF7GVVI+Fzw4Py0E2VYZenEffF53ukw7q2uUcbXbFWOxUUPdb+EdwH
6CWszgoEw7jXwRHHlErwDOdsWmbqgwwbMkAUgejzckWSzY2SoYip5nVH975gj3u6V5hNa4fuGnv6
YrIHcbOBiTEWBuDAJUSygZQddBZD7EjpVvoCNWEO2CApE7wFwLoqDmnnmOE4BvXRFP63ZWuZUF06
MGhJipkQeqQD1eJViEAOolQZkBSqzr11IiqMsJkI7AZz6zAQTHlMmlCNSK9tN5ejLO8d13J44DPH
fbKYdx/T1m4XvwccDetUYvycT9ArV24FyKkOi4/Tw5ZIO2hThL2clZwarUIoEViQPnFQYpxWlJ4Q
YiROLI9nKr8n3P3MB6f3P24GHPl99A1TE9JHapgN3StE2BJTQJW80XSwgHpfGgaH7KJ0ye554NSc
HMHNKzZUuTuUAEiBpaMMlix4ks426xa5/vZF45Y5joiujkw+tGb6BeT+ZP2wKEZAePeDdV79fPDg
09XBfxGyvvYXL1iv0m866jijS3E3g8oZzl1iVZSs2qy9gy18H54xbiN1d4ksCRxwmkDEphxWJkcc
MdWXYBm3w5CsW9Fsp5e0mQhmBqSTqNKAKgCFJXozw13Ogd4Ce58RzB4FbZH9vtMvQXJgbQM9Ij39
iXLDnaiXUFOj19bvG0LaFHefQznd6S7lr01zGGSrEAd95uld2U/2clqjmP6nWPU998r8/KzDxKDb
ECJoJraZcoI/Mp4Y6KcWgpLZENuNikfnTCKOygr0OwkLyV3tZToevLS51NfBsHWFYalhXQFIgl+E
M7BCdf4P8n+S6OwC+oEYwYmt/AfVMaHBnw3wp7zYEtkwmjMY9puXZr/rRKvHrUYdedp/TbjZoCkz
nW0pTOeKaWSIseZwcRNJWXbXC+QzRg/SOni9ld/UOwfuYgcsazE0cjGP5Gm8MEAvByl1SzcyuqPx
LWwWo3JJMzGrLDo6GQdgqGAxT0DhrOMrPqBAFhToiRRAtL15AY2HioiadTxEewaBKeh/niQCSzt7
2DRNiSs2L8cIItcAkFZah6vZL1VOqvt+OwqmwnOR2pPCu9PCic53cyU/v9zyQKzFmlK9bHScbweP
Mk9fMueG9hagh53LrCyacaXEpUDlIJrNLGbRX+Bjn/slUELpt3+HQcMTXeQjR3Klu6874S5tQbdW
9tgjVSkMGzWaiopIXCY4rEMoKq9dHIvIZF6wnKZ/XpLjoulW1kMes/zxwsaQqDqZH98X6Z2/6eOR
wydVqgaKcCf2FUPSqu9pctgmhQog9zc4X0WnvYXor4YYGkFwxwrpLeAOYDYjFpCb1y0C7msSYYKh
M01i+MHO9mEMJSgeb0LGjLhkq5qcQBaRM8QDVH/rk8oSReIq4eH4DU7zxPe/h4sUPGfGM3Y+3r5f
3UztWBAeIYyjNnJxDcjC5Xhb0DdXJgyUxnm9IK/j99Or/NqBIxwy6VAZ5V5ByhGDT53gmifpbuZg
fLJ3j5jvGwwGE6UBqRZtq/Of3q6pttwQA/UjKZ8++5wWcYhBRACqnbdo474sSKs0JbBZtOeKTSNd
evloUml9folMdjCtyuhF+6bYjTniwZPN5EJVoGWbHtnb1LE8a1s0kWSXnSdq+iCZV5E4fzTeyLch
gqOtmYjb7eccbtPqOwSYmj01yG9kWzBq7JHAgElwtjUbbTNIih4FUDbqCyTk6Cp6VWXUgzPP8mOp
bW7oN5Z8I6CWAdMcSBDt9GFyfnADgMHJ8GAXm4XlorHkNiZyfhpM9H4dexVZwTQukjjBCDovRVsm
P/5ZYkGbcjOu5wWploIj76mZPweKLvCWpczIqimNjE8xtVv+bkzJ3VJLrrYVJvpBjS71qsYW2GTc
7KX+Qj+pfYyeWkm5UU2hkgIbw4ph5Aa6cln4aPaq01x/k5N16LHrd5Ic7ClaoNACtOFiJ9pgQgxR
mNl1OkBTYhv/bINRYuugGES8SW08imDme7TTEqMjUShI5AZD86rbR+muPK4qLu0z8UvKOZ+oua3n
hgf94OqWMlCGAYQ3eEECm+FSo/1579sKstsqXhs/FiYNkXp/P3HE8+cmyfdqhV13sI1u42AaXRG2
nOKZReU5+QpVZvCIhfgqeAU70465p4SgYIiNxtwv3BCeLJgzMs/INCH1cbRcumYwef8ymO9DDnbV
nUtJbCHNI+81SGwURn9f/47HuHRYL8bHXuNdFoSbDzFXKX5gd7vptJTWbHfBPFnYNUbZ2qqxSCT+
YOqhLloHTh/DIwxqEwjXkoSVS4ky/iOzrFbPGHLU13ltEr1YPJuQeQmjdyVhkTWnSTZa+CDs+pcg
Z2fou8v4D92LOz/bpKOVrlDUCUET32TeZKGekSVaT7k6JpS2lp6AqLw1J792FIlMqP2gvitWlF4p
DVw1d8rsl6CkzfkNYO/XDieOZ/1xBG4hQvybcbkXQFpkBeKT/ahGL3KTsJQ/2ghg0Xi+rHsVv7oU
tMNXwsUq0sjH7/mG7VwXaBte80jR5g0r2zSZqAxb1oFt4cZvQjn+fJN7vKHGei/G/EFghJCZD6MG
d5l864pa2N/guiXLVZqQtAKZe9/NVHNSe0d9Pqn5Wxf2ulydBY117eluxnry/jY2KQy5vEAZqSO9
gTLi+0wQsFwhBK0P9Xz2GCxrg0Ha5QJmdWrl8+XKkGVIRDE3Pcx8stQlnAdCaRkqshfEqQdVne4M
XRUW55D0yhAjadqBeLGp3zO9n5GRDC33vRSF/aSH80WsUFJn8TKcK+9BKWeBBFxl47DDXLwZkdAL
b/yJjw4l8vOO2cCM9RBeFIVoYsdRYILmP3yVn8j1Z7+Q2Hk/7v18wFktOqM3FDmKbu0rCQM8oLHE
QF3xTwBsCisQ18HzyzXR0+gOe8yucqU6Vn/EwGi68L2xaeBf6rGGdW1v2zyII0i4rAE9QQDuzGWv
zHzXG2tGeMjHGK+v4qCg+NzmlPJfbUZLuVTz19Oo62jXKe2oCYFUmQ5sy/jiIIihqxYyigCGGzA0
BXET970aSU8wKs83BbTH7ezhjDil04LmK/mvOKBrr7LDxdEvPNwoOUUPKIlOOXtMjHofx4AGGa0J
Zu1S938x7pvj+WDphCAK7rgMrKwRKhtZERvw+13hfTQrnin29fk4asw5kftoHwtbY9WDI7RCEKKp
PiPMwkxZ+e+D06DeR8LFQZnhmtjHhz1LxHNxoSvANK96RWFC/GPe8E2TdJPyuEnhTdjeLYL/poZS
AYLmh96iwQ2h0RbDMSUo2ljFTzS4dvlr5XIyNueM3TosRjhUOU6La//WUr9yCB+J39u/mMIN9Bhz
XXyyMyJISscJCtq8kWMUOQT/2mstDrhPz7Nsicq/esum07E8RNsGnkGAkS01Gl/nw8DUlQlNeBci
NKrbhUZGfse+fQJJkJgkdwtlOJdVUq+xrGDIWptmOuIle5VlRdNBpYpkRds74xnVfVZsndfW12Qb
sd5YnATsDL54IN/7xgbJ+QKA7dXHWT+PvcYD7uA4aJhp1gqbS5/bDSL5K5J6Y70d5JZx14e1xyKT
M62gG89YRfDUmEpXLf+SfMhGJauAHtc7yupXgrA/rSsHtG1zNmSqUogx+YqOkiNQL2r7fWnv1/3q
+PC2LuzrvwzcLdR/14c4hOZJQ1ULliCUDiEmvGmRh2qS0CufHC2ffIcdHDR6w8KwAt+H9Aj+t4cu
HCr7cgK8mAN4+x5FITBzWn3LY/C4NuVsjxXGVcDnc0RfzGKuEO12JkXHn2Guy8vdH1+ckl2TsbXX
lEGHVfjKAqNEkKe7Fv4gpOMrfxpz/v0GtBqscrq6EKlMgJtAau+wFGAzyqLM/+wVUqerq4j0Iyda
ImlhbU8ZGSkJzmRiuTaOHUHsh1UVTlD9l5XaXTZpHdcwbHX+fjerYvcALJswQ00MQ1cl2SeFvQLY
HvqBsY4iSwExeWHRBfnNIoh2j7i0Aiq0S98x93KRyK7rcsZPG4quB6qg7Mbq2jp79XTMNi3KoWWR
k3liVUzftgGqhBRpbCfoOU+hVq5gOcnoNtJbH+xAFcCWbdfdHRz18bmxjyTGpftRQhkq2GeLzyaE
ACiqxvlSVz1GDFD6S7gfByGMpeTLlOmrYKfjffUqsBQqE9fynw6gM5ZfqOCR9mmvVPLeeH0BPRwy
KwM5YBXSbl813Wl4J8NUTkjwGwH2fmJMbZKR4SVUyGsPfPjGcAB7VsHO4TgKoVggEfakUiBbAVK6
pfFXnxEhnBH7yNW/Ux/3OalSpfPcQNWAeRKgBAr9bvkj/hBh7StsnLTpG6FFX8Q5sQYtPIduN2vF
+Ypxt9hwWS2AYlIR0aE/wdzV5XdSjtXIXdWk3Yhz4nYKgnfBCECBhGPZ8Y184gub1rtVp1eX/BUy
jE7cs+4uDuSiXoofD1Oo2r4Ge+cBeZX7V3QM6aST3J4o8YavpiAJslCxnPQZ/utpo7M7DCxRMvYT
yWDBXrfw/iWRZxZNlSNbJsmTWDelq4PZ1DqrQ9u2sAa3VP0CBkshdUBfJq1DV7q8YDodcVDVQeaV
7TnBNlivE9LsPY7SwynHHPkG7hEXlzFLR3Y4Pcp3FjV6t/1r8QHSgZkyzq5P53xOQJMhBOiSuA/V
jubqDxprVvtZIlpf8x+VpjID3m2YxXwYWhp3wB3q+70H1mkWLPb5byP08K7HXJQ566nVS6RQA9tm
WTtyWKFkhAKpET3eQKX9Vigy0kkraAJ/DYsDOZzGCHSGY1ttrqPxQiK+guPJ+jCCZp/uJMYQ65gX
cc+ZefyUhT64pO8CBQHAXt7bretIGLQ05aCK9oNE4zR1uFxiiHZr+fr0qHo0O92S1OkAPaDu2vTf
Pw4s+ngW7ODF52iZSx8+6aab3j5kU4U+ydYLK4EC0pn8OslRckwxuwNVJ1P8io3LeZtsaMRMb3N2
PCVlnw7Q/+hQ+OkytcJXXls1LLjLO5UiCbCRM3kWdJQwPsI0CwUApOaGrGY0zNozXVtv/gqQgUYm
Q/FQ/XgnJrmWRDcaOR5g1TFUckBKKidVU322BN7SOOBMQ+QoJ/sdLY2sP+dU0ny96AY8MHEZgSvT
oLnht0iZ2PFl0+ZHNjMAPAN80iQ/ks7mUTLu+wWBw57XvTtqdTZxnKzg/BRkaJUy54bjruQTKJ8s
nRldI9kE9+BIYjbUwzBRgBbzeGT8C7YHrzY5D4GkgITBc2D0YUiUsTnbgJhvZ3ItwhagUIFEuQXb
n7ZeeaxDHxBwA9cFktdtJy1u8dPVcq2zWuxh5uSvq58/L0/m9xu43t7KW2jXHb7UnYBgV9GvFdKI
lrCojviRKfXSsvbugf5K0INq0gmaOyrQBVqQjcqmXsck/716IlnZC5AAHki8sLn6uLVuphWwwvA5
Z5dhuMWdyBJ3M6Q/qDJ2aDYKe2LfWRubC1cRgvsAtOafVXJVkOtp0qlrTXzyhfhDDw8hwoSe9NaF
52W9Ms0M0ScoBePETitjSvNnAAD3oInv6T/ftgnIys7v04ZPpL9ciIAKz45TyNz+C+wCNNOIXGde
mOYL5I+4oKLO7kSJSglp6MZkQlQBefJilqN5zEbfjRB+vd2VzwwkO7hK69yQyhSvUmsyrwXyytqX
0TtG58DSJpxMrWBXOUr6W8KEVKnOi8PlYAb02vPRzg1gSBSLJrvAsWBkjxn4MAMKfqdmKyT61bDE
d3jaJaERiveVAN+lG/c6U7ZsCyVIdXJ6f3gVM/DW5uNsNOP3kp84phtamNtGO4yUjkTinLRtq70k
4yH6ODQZVfJqJ+qjqqwhZl6Jro4P4gnnl0nBKPIlcLIzZY4Vj7QxbxYe2cJAS+KwPwzCf8HyooMY
grNzcu2yNFtdhnMxQqTTI6i7CHS+gwndTsXVhrOyBxuklqLICXyUKJByHvEKIjex7FOSNI4bOI5a
SEmEscE/s9ClLiK+55PEum+aZ7f6zT5TsDa9vPqr5swzYcGmSH6SJwJFbg6U4/7eJZ4GorEA6Axk
iYN5riM8NRtC8NwBIvHhnjR/ho+5zzEM8X+JI6u+VAuBtiqu9/6ib73k38jEqzveBsaehvwzBpPY
SlYzH8BOUPYboQqqquEBk3uGLjmZZL8jHzFM/eWKNXD09tvXJhDHE5Yfk07sBN8JYc9HouYgYnnF
+dWs69MEvCQVFOFS0YK+QKTWSjcEX5sEsqDuDSClzGe2ed9GsK5HX/NtEK4F84y+w8l1Zl8wk9VM
OYpEseQsqMyRru4F2cZ5eeYB5SPnohJOVdU9g/bCe1kiQ45y7NJ8T13/GPnoT3hhTEkyBr2qWx1I
eVB6aOAa27d3TDj+2HpbpoMgw+9mxjDLHP5HDDPZm06Gg+gK2Uf5ZP2SFLmYMzdPZ5aR1rP6Fgj3
Fig90DNADgw89Ot7SB/jxZbF4VQa/TVGjEe5xYdXRytCIBgpwjY94tanc4akiIDyxnPYl7iLmlA7
LyztS3Ew2LbaH3IWTE6414ci82vZyq/BWl6+awhqCtShOSZUsBXoXtki8ioYfEGO/W0k8BBTMMr1
HwvuMVSN13dFRVNrQOtgPgsbRFV27G6iTghhuL5u24yd70lHbrFm+AWP0zIz+QdVLsATD72/rfL0
3exc8eRlta36R2iODA/RwMn9tdFOlgNOEHlzOfwKr+5dCSh/MAEpOn1rhbGMAd1g4PueA8WXoMkX
7b9K/7AkXKmKoqadV25BA7o9Zg4TINovVkt4LqCkGvJIyHzdoV9aP4VgMdAlagQ/CzfZgjJYyL+F
M2Ay2YAMf/IQyjsY8wf0uFrzmBuvRZNxUINZhyh6Ebsf0fcS1MNOabCmBxnfJwRYUG/kJlH1BAdB
s9NIEyH9RurfRxMfivOoAMd/kaqP7iTeuKfOo0JSlf3MGzYj3t03IDpKn1NlX7DNELWwQBBgXigQ
GN2SUmAhd3e1I6aQBsr5RpKdhmnc4mN+GgsFWkF/LGPBd+1nIpDSEhpKHD5ycCUy5PGW1AvbqjQe
ZImiR14ILZTaq8Kp81cpf1w5U+qnAbL3yTZwxY4s8lKqLUrrT75kM2DlLQxpumNqGpvSxIMGceUt
U50C6mJKpahhFW3rqdl03GIND6F2IFRItMqGssZOKrhavj0cBjoIAilnsSOzg+SrCyFf73toBge+
ueBje6Qgd90QFmu2HVV/5dT98/MN6BuR7SE4gwRt3cuygPtO2iZKtzPChiYke4Mz22jYgVuA1Yfh
ZxFzhgfbXWwfzJM4Kx2pHQIgAooETloXkwQWBZc7HLyMfgaFeLBL0Q9Kiket47m068/t7YKTC98d
kKtDgMlB8RNnBX8nB/inhCboLEv2vYGOwhS88k7EoHDeoIP8qahpPhl18ynWPtkA0R/wZfeeLgiO
2QzVoMMxkFyWKZVcC+GWju+hdombs9PphoiGvnqSinPxzlHUTh0thumGoYrsbJOfkeMKEx7mY3dT
HPCO+Pu7+Lk7S8QN/YEaqfT/fzy+bu0mojH4YhPDZz125tI61xcO//iHXKOnfQbAerI1lgvjBTY5
umaLfBbaW3IARDjVEfMx4mvj5jWIGWIY54ZcYY32wG0d9kCVAF14A+eJog6qhV4lLmhtFAF8C01z
IisW9ye5VABcI+oaLT8EBjFFD3b+JRn0b9YiOL0TCc9Z0XjuXy81XatKbKisj++Ku1An6FpzbM3R
r9BDDXr9SNf3IG50gF21rfYfzJtDWsHvlsknQFSf/eQKbVQxzlCUm0aUAa5es2XJc9xLnTcJePXS
fyKgtlVYZi9W+o6KhpRRRa+R/ZCCrNTWDgFNQs1mkWAbQq6KtNgqJscs3nAaBziYhSXn+oUAoMmc
qN+RKjlvKlx0lqpSzSloOJk9lNQkXaP4efeoIwFln+6L9AZfZCUe2a96mfP7qL1migr834m6shoO
9LdB3GWgqRBfUBAjZOOKEYqWMSCEQLAk2m5H5zHCaIC5tMPeS8WZ4WnTyCSkCforSoYmZSPZjOCG
tOkToSMaoxVfVBgkJ30+Hf5Q3vcKXbWaNqIBR1AYTBRK+ZPLrGmXqUXaiOZZp9cnfb3QPhrm5JrZ
kwQbJlxqShpElrH/j0bLkJkBGUMlSOwg4LZZKRyChRbOoPI+Zq16hwI6KkCQb7Ziy9UNOYnF+qfC
uiusMoCdcobgHe1La8t7W7Vz2wdDN16/xRexefnbFITj4okYk1hmgRvgxMR4cTL6JgllbsiZm2oB
r/HsB+PV2vMhSZr99eTTl8uGxs931h2w2XH5CABUtTGXl5lUbVTVi4c0Ld/WfXhUMJmuPH2c8/VF
r1UIUN3IZ5vOCUs+LmI6QLrXAUPfa11ejXeJTvUmNG/G8hZVnp67OuCyOLx3eXyt08DfIaH/Qys7
uNSkYzla9kRAAAg1TVtKBGGdf7e72tooJgmVj0PuFtMSRSBlbSPcffPhh1C0/uTHT7mO4mQsScpX
JNZZuCm4b81sWuTQKNCo1JmcsMIluitwFKJ7wFkTD9cbE5K1eOGdjioBzZz/cgHzO4xSqlZuUyZh
vpsMO24wajGnSTyB/dweWZaEMVVun13WscFp23RAiYYKZtd/bhZ6d0HiRnewKbHiu0FUfQOxJovv
CSd+D+t6iYUbC7y0nsCXuRjA6ahcvyoi2Epa+aNgpvNiqYNFyfFxlEQs/ZqbQs2jzZu9p3C5Bz4m
xPzYv4RvOWnaFCSjfrdkoEE0SLwMeUUfZMB7XFcTKcGaor1KHVY0dX0CAmmjbaO3Gtd6xO5OeDbD
udmFj3c1yFVtoibKfCpvrWJX7+zaymsDSyZNAp1o8NFaoNvb4cNrmKZ35xKEryhL6SMLBV/WM3P3
7S8Gg4LluYnQYYZO1L8F5OVcENJ6B5qkIb9uOcZIbezN1cSvQpSGHv306deg6iTRCM2TxWZcDFQG
RHV/TxXHjCENCbQieqWvFmIQOFgHCniscDvEqMEfBgK4ntWnkSmY0qGquvnK5QV0ANS2cnNVFU80
LUVBo530w4SvznYwhZZ/EsdKVafFS5ckgbio0zhmu12kAXsdU8fJnwFyinlDDauFXz9LjEPavkC9
lG/4jJFN8cFSUOybUAfglcU8P16OJBlxMuZ0ab2/o6IaIF3ywiQphDdNZdQh4wJ4InC3O1w4TM1H
VjF1PzKRJVRD/2F1GCJQYGWl8NTb0KvDZfYFyV1wdwcquiKtsa3QVUKHCMOw84ey+IuqKiZ77waV
+dvJLveu4dSQmesnjzJOiZ2d2PYkUtpBmx8ADzKePL0h/KoUULTRKxiOpZREb+6KwWOuBdxMFGgq
cMvJiC8VkKOWPMF83yIdTPF+ls3abEtCXuZMhzsLGY4kIfTMnZ0iCnc6knEOYBqhES4jFo/juLqW
yCoEfg13hb5sfbTDX3bGRBJ2xeMsJ5yyUiYOcyCAPmxKqY+CGJajS9BhGUfi4GB4hr72I+k+1DAs
SCxj6k1qWnBqQnR55x3kudx9DV/8ZOp5I1W36Crn7rJrWt0gfu5o7u4fJ64B4hClUAKqU6uQwzO0
8viT5omDwq1mRtVl6uiC3oeDFifhc4qOQINDzo1BIw4H8F/gAYBhnx5MEG7tWaoWYjj0Ok+fAxNl
YoW/lXDP595KGDcLjEAFAIg8f1/zkbh4YXPtMPex665w/0IzqXEQ+Xov7slHxdsUiG+u7F2TogL4
MFGk6timjhrZbWslfc2q9vXQQs9ctxN9D0QBrYd95TYRCL65GcuZvPif8+XAd3m1VI7Zx0mdIhPZ
RLu1drramNa4OXITEpdLgkoQGqYEL1y5nfYYclIZE20dcw6XStt/HNmQwI2iqyXGYa1UNPvs5C8G
pXQxO/AYtN7JTs8tJbTJ7/oW+8aCdvqam1IVuxjdWjSJrbTB/vO0hx/j5pIxCOnT404tEeQ8YRHo
brTYLhz9KzRLCRkMgrWFyNbtvZ953zd/enYBmDj7CKxp/3BqD5l/uxuyGtYnHs5gU4IHDfiFSxcR
zkGDxdW2CxG6p9h7mEOpttQLO5vkAFEfSe6lcH/o5+pcvaNjWGFB9LsCLV0PSbZpDGSd3kwiAdAS
OGzVjGE8OPL/oHwwl7R7+4Ux0XHjpFK/F/3k9mzw8nuwszzZ8XSs1mpzFjLJrMoYyCNN5VFFLzLj
T7La+pe5MC0PIVGyUWN6QTKqKZpprCvNlw7s351GBr9WAYFx7VFXF+5tdcyLPszUiCp5rjCTHZUH
y4Jj67HqrVLbx41EmJwFQ3Ie7nNB17ODabV46F3G7h7OoIDXeVveLsY8OYomHqpV+7tDyxioORu1
LcFazOKZDSdQI8sBCcEcA0miz/iRZ49hTpMVBcKYvEGAMMbIrIuWTbAI1mD15paOz4c8yK4mKzeZ
R023A9hLopst90Fs3ad+fIFeis5Vv0VWXqvUbIQWT1R09MeirM0FgoXTK8gMio8wjszIgmrU2i64
HQAkiUdk0BrGY1ABpDkNH2qgB9Rmj4iFbixFKB5k4jlKdxVhabbvb8HXHAzGG9kGWOscOAx9bMqh
IXoSbtkTli5/cMyRZSU3DDy2OgeprIXJSQtk94B4zbi5HC5tni//CokP4ccBoozuMvQt17ECWoIl
0icTeOYx/cjmuRQTn8ksKkETu8joW/kO/yrj5hdN20/G538p7Kj2wm/vG2b1llmIIu+qnCLXKvPC
3v1l2DbJLRVmfu7sHeYQim6uReWfA91Z3xRCfnYbsz1S69/BqJR8u13Hri34BAW0vKdNte9469GD
HicvWVXfbZtPI0ikQKn7dyFjLwtEb1T67DGd7KDO/g1nUuAz4XaHRIPdbFlg9yK+eFQWL6L8M4y4
kAGu6iz9fzxaDffj+6z8xCnVRZpy/Nrmcw+fQ3OxSdgFOK0KcEBXj6Uo2dJw0K+/mRKQKhOKmhLy
a+84MtPp2XXO4EH7FpcmwrFqQJT8qF/Sk2V8Nn2hIQ0sOw5Cw0GIU30pMHViEoFqBbrFHBFFewm0
rK1YE8KEwINU0jEESQSzT5Eq+NPPwP7Y4VICzcsUSwaW2pG+yGoqGAaXfHaIkKXLHNXevEFdiPi6
9tyMGbOfTCS7t8KndK0E4cS4Z4T9xdGb4T1Q4Fd918yYvdWWOAjEUsP5gWYZ/vplm1Ac897QrEZP
ZTsWui/c0fn4HJS+aqPzbvogEQ/DEQP8yk2cSCveD8LAS5HTuRDx3HIrDbM1I1UG1mGGtRuz6RAm
1sZhCi8N1+86CcMsREAtA3ZRU3yXt03jZHwZkJdPI+LsLaHusua2kwKfcOSb3JW8bj4gjaFuttCa
loZgFD+IvnKvqW/TD2vsaeNdrjo5JZ6XYwH5iOgd3RSHbmWcgIWe/3HkIXiyMB8CD6Q3PuCDZmlz
frvpFVAL8waxwaiJPK8BpwIOOkJoeO5IBSbxo8EWkDUNUebX9X8z+5dC78Xja4aDRErWa4ktqV38
356A0SRoJEf3q2sh7d6Ceoyq++CcE1NkOWLhMp2GP/AXLZ4a5Ps7/pXQvjGIFMhtqmNJFlyXgPnH
9CSSc5bANWbCbSXeQeKjBo80YwNnmgS5Dc1Igv+kAjcrDSNG9trnD96zUUOOmGKqj/ytrgpesJEz
FmwGXMYUOwueHESNeqF2sB76g9lxd28hoKp8HfesHMy9JjwXwd87oGlRSGJbzl2FwyHNsTnh0x+Q
jg2UbXgubEMhfhyfo/bkV+epwQIadwmBaJ11YA+vsSa1ZyBtfjRzNl3Ws/CTvmb3UlZf+B3taiZL
Kvc1cjDfwxb1cBD3L2Bj1yQZh62aCHQpV7HLXQdrZMvBHU5T4r+O+zwyYzD5qKLhE6DmGrLNXnLW
VVnwx18xLt7cSzRCTSyG9JCMHWynbQczrsUnbaXm9WnRv8JpkJ0lM6I1xoiZLHroGfnpOqxoAej8
4alDtEI/JoWOrovbZh+3F1RSa4eC5zXEqPQW94FOjjmZViEo4sLQ1/4nWWfPMhLZREOn9kgJoyP2
usupB3za5WspEk/srtDHPccRtvzK4fYCc/puP+htuoXbhOx1VO5zWD+HI4cyhkGPTlpMLNNwb9QY
ot0M8uWJ4mIcY2Y1iVFvjvHSDloSG8nrB4wQP2OUxQ98hf+itBctJ/e443h0fdDy3z5gEOdpdkzS
9J3taLrd8D1Nc8wj58xZ9vO6dMg7hUb2FAH1P7/sQn5XitjrfMF+fgSotG0HjSFqk7s+UQJXC3JE
atdqXotDCfb6zkJktbOftMAqKPcfgdg51S8AIc6yvfRjlnbOE0K+GjqPa1ml2x3FFP1G9790VZ2r
IoUMe5ZqlQo0Tq0ztAw9ir9rzZvFzrNqn01DZGydB1VW/T8DvHXil+oB+BELh9exUbPdBEKJGd1w
uudILh8z12P35bJ+tT9h1M35xIGQqh0x1ErVXC9bqn6kECQRAA/asnftZoMtyq1TgW92AK+fDDRX
F72Nue0OAcDwbWMYxYSOkYbDti5xv9MDxDa48vd65Q6E/1mSyHgkeRwgCbEek/MXhJ3voiEIpaXH
c5NU+2ZnNADCpYpCJ7ykUW51J5PZ04+kFqZLO2ecoYDO3aPxTplr2zSsDrjir8gYNuhpxY8SLZ4m
fjlXjP2xX9sSwYivJaz8LedHfufQ/cBvwnwJwcjR0j5ak8cl7uiewwTxukUkKuhyOa7JAIL7h1fI
QWW8NJSpJCeNwLfut1aL8szmkQz1t2InHHSG54RzPBeM9v8pLlDgbUV/8XzJJM1UVT6SaONHdZ4d
nz+nnWr73pab33mLgSj4lBIh8fGM7YTWf2tRPYOomkKuJkupgMBn7e/EqGxxLXv954P7402RY3SE
yriFggrCBxJ03/mjeWEEWfdBhBvyiKjH5P3fKzda03da2JVddUXSnmGveGQ1oHZJiBXlbH3jJE9y
ykhoq7cDsrjIgv5mUqy/ssrYPHNcFQ5/xsNAKe2rUe8x8MZEhchHv2MQ1RwJv65Rosnvx8BoItBm
uPoE9hlJ7w1cFkLYhOI+fLHGsTVGEj5rUadvuaQzdk9NHyuAlh1nnAIFnXztrgVR2PlxMN6vxTz6
9QUkmOdUr/ylEtSrpRhzHO0Mw9qMEflT/nVuOnTS+hDap3aTIT8io3rFbNjCDReBKeT2dSXqv3PJ
UqTVRNq5MLg0fyJCqVN+Z7lywiNoH6pmUYhg1CMMEJFDGSP/PZW1yic1bnoJn7mZj86yuY0ABU87
TTlYNw7UXBUFQrkbCcUyULZ1eXFrjrQ2cmtdkM2hFiTuLUOfreGsrC5C7R1uuVZCAnEZ0BvAZIKT
0eCfaz6lJQU0T2c8MkCJTpQ35ltOslvwtxqsVAFHpNgEeiMiuD7EkMG11kfv3rIpcLs/4VcGdzHw
xVaD+0GO1tz2BfzHatpLz6glqg60gXHw54WjPNJVXKhmDa5sEOlyZyqZcvOBl7hWanychcMnt7j+
ATfUBJdaoPQ/QKwB/j0u+GGDEV5qHcKCSV1gCQWAoOBqCajuAh2lDGWMxuUphytVQ8R4UwCCM5Nl
Rkhv8V3ef/MkiCE3sgfxWyDBAaOKbHm8gRR0qPuZV2N0AIf3qArLryXrsAuAVmgZZ73sJLnZw+QX
DnL4Osto3u4CVbmJ8nedKgvkzypLmmFyMHuSRIZBlquzMxPsogK5IDy1gov5s8guP/Wp0v2zYVa8
AaC1eexyUxVWuXAkvkR1oPXKVSJBTzNyFt09Tzj5ufGm1gQMm+eiThqo1iFmjC8WXolMcrEyFJAI
ie0xF6cdQwmgsFGuKttD146Mj4L//i9sA8d7E0W6+mz3W5xcFdf1tBW9NKPkQD9aj8GLR1m1X42c
43NbT2kSEi3bRxstF5pD7NvSJlvKaxCfxJ8FJxIHyu2PR2k3WahKKwQiyV/GC/gXScSGMjO+1w7L
C5cBMPwpVJ1envHaHF2Poy68wUdTMko1HFSYcF6kiRcR3z76AAwIT/9RjNHpoAsT+9ttgaioTBA9
hKc5Q3gThuw6GUNZejFifQaaidKDlZtV7Vf2pCB+JlHDiWY1O4CtoQS+A+p8b4dPexoIbE9ooYTG
KIsy29x9HhtUhW8BX7VsoLMYYNkrAg5Jqd15W/kK6mZnwcKXTUuz8r5eHXzyZuURUkbG2pD4i7I2
3dJtWZkpFBjFksF6KrEkqpJwvlwJIdglLnHXkCNqVH8vYfJcwHa5YU0RVEttGpE6t3uxZKhymXZn
hqg0HesNerztwd3/KpmEDeMDvpBJ3vU/mSGC3CDZhBu2wzuHoZ9rZulJQ0i2QWof+qyg0DTVziIj
tId10soZUkafbKFL76lIMa79YkXPBXzlp3EAEWIRtyg2n6qDM0Qao/oS+lTIWy3mte90lJ3ksXWc
cZB8Bgpj0eQ8Jyg0kdKJbG0zkpAcvLd6NiQ4LDnO+KWr+LZUlOyiIUfthUJp+NoPzfs4OSxvjNDF
N5BbNBNikGdN8OXpfyDi20qt3eJ4cqcPJ16ZF0sUitVnCc5+VS744mX7tRN1SzsHaD6bNhDlyeBE
DJ6bg9+eucvvftqRIOrn6B2wjRehTlOJ+SLHoeDy7Xfk9LZDQCnLC/uBAIM0BxqfdFCYjWVoYcdo
YQoTePiqxJstWwXjia98qwh3yN8QF65344w2JtqGCRy79VcN1B5nFPwTpeZxam1HGJ2T2d5B4lcH
5QWS1h6pVvxlYjyl5qOIFDjIIx5MDbS7Jmwa9SI91pPs9wp1gYn6DOb/3dtJleohi5IHIJ9Ynm/v
01J67Z9k+4xp4hsPumIfuqHD2Lts9IPkZ7qJnk4ZRoso7EDYb/vwY8RkD8J3uKANriZswXxlAURs
rNvwA4//BxKZ96x0Uew2shD14PfVkDIhz9aYD5CnyaNGF2aOychryw0oPlx2XtJCQaA7jak+27XG
Nv1DA+F400V/gUS/JD8z95XfxIr3Gg6fXzfMPeg9u1oPVlnzC0WghAzqKxKjkDrLEdK4vTeKdmD9
xyCcW3xIIUGHIXrTZ1uh3T2eeE/w2SS/dneW8WB5CtMzZZul9NBucLoSNEFef70NGNF4+j+fHbkg
1RFzXujllxFBRjZ0032eSupyeydMV4efMgfgb5bm0BbHdvAzjCvDJUny3RQwtpXSEhRxVyx5RbwW
gjo3I+UlzrWjJR8+mhEwXJQq8pBZath6WMaTrR6kiN4XLpJk6Zcx4/qBjS6mbnJ6SPvS68XNNRlA
NWRbEMdqB35I3zeMU7CjGViInaYwPOIHfbAuqXOuq9oDhaRHLs70tnZh+dK5QNtjRxai2sret9Xx
NGszW27Te/9WQtqMSN5JgmWZyoW8WZRLtQHoRmTHTR6M9ZvmV2l+pyqTGa2bdWA9RltBPf+kQKQ0
/z6XcN9Uil6ybAZZeOQIMxpIJOoa6VZ3rv0XKGNQV3qkmRkQwVOgCfuFQny98ntzOkq7BJmrLEQy
EwF6HPqhHHzNL+ZLBWfcNdjHx9q717mZ8MS5QO+UL0OwNF5D9bgoq+FxAOirYeJM28sZsOWcgw6w
OKGDHWJrRD7ZLYcYM0TSOF82D8hhlhe2uepWDJtvTRvRDs8Q1nAnnFzyq71XxO7SuUGj4fNuLhbu
NpFvKyGTlrg9zgLYA47FMDreina9TcpqijNYIOn2iifCkLYrLjelBzP5UBdSN1PBmHAjhObScwCz
92oIFEPhCzV5e51taOupZiUOU2B7BMZIOsO2+WNqAVGjBUEmokakwzMMlUysluh87CYCpDbplPzh
uuYnlFAdXncGwkZz1HaHFaSkYLojR7IW9qZDNYEnA5bT2QM8j8dlDgrihfETMzrB7RXJbyHhoQoV
laA9UQih2yeLAxkcXQsZNmiRTwVBp0WlBMavm4rpmWTOZDP6Fy+M1qMpm35xxauy2XnPv21IEPop
vxnReIZFR3GSHOLsqKIxjmgsaei3HVGRuPlAxIi6wtOKVF70kheTu4lh23NlPyU4BGicH2zIRoVh
zTBa2pfx6i9xdoCDegjYZ9zo9tNomjZ7sWRmYgrLABkTWReQeloCSqgXzYHViHQHt+sxhhAaO3x1
tiIr6iIt/qZjVlbEGxAFGXjt8XqfBvlxps6V89SbOldmSy4v7YEI6hRYuBIlDUfdimBsL05UlmWN
BEgEbez9Tjgkk6nqtLDnZX7GW/3K25N8Noslyfw4j+8AYLC5f+g+BTfM6H+vw6sSo5dmEBRPeX2E
DF7doR4MOZMqQxmOO6/42cqxB+b+uZimk/PaLQjKBkuV6/7yhvn/V8n3Mfpt/dJt9ipqQahoMN+S
fkGX4sslAvRgkb+WGbkHyCcSq5obmffdmWSsHbFBldXmcxBs0hppXTlBx4RoUG9whqBAtDGBCWJS
L43PLKrrWPLaNEowcW4TmNN6tD2xyxv5CL7JN8sX/9S67vAoPmqVYdNRnU7kPjKbNM/Gq99xCHTo
RMPFuexGf3lQTYyOEP74ehUSPynTk3mMP9dPU7K5w3XBsl8sPSWKe6X1A6w8sv62DBbNgyb7WCG6
aGLMZgA2X5jQnPBgWRlPz+2vKRtfilRk2w1OsCro7mMiUqUOtGwo9ZcglmiRJEncmyZo4I40V3vo
EU02cDsVpL2XGECCOGd+gwaypm5e5butvr+MdMZxhBAEKmhF9Vzcgco+HksN6Y2C4k0N6sG0IUQx
PbY5anrE2mKiMxmWzQChOzCurpD974JOEKU9GD/VxgmAqb4TdVWLxxuWLbVnqzVurXVQFL/cST0U
pzHPyeuEQi0dtxnbDPgF0/XWz27x0Vn73ekbCIchiZh4G9cnL8SVEJD61tag4k0A9lfZ5k2yjEvL
al21ZcqgxMgRAtPrt9TCGC+6EWGGe1rwHWWhuc449sp8q5XYtDIpcMSxzfLAYOKTf+S9uqwuMEP7
4lLcFluLmfkjf/Q6IzB/WUusJ87rxKCmN8LFjicADljBMyn8M/AsyGYjIVfyPezOUKkAr6cgZgkd
RAxZdpse0SVogvrKEGVasLoUVQcyU+4JnGgBtU0CAsGo+WepXQ4Uw+7ZyV5r7Gv5HIz4u2+aXO4v
EEiKhKtbPPkDxXhJENJ1RXlCrvG1iZT4yLnqMvqc6RFPxT6vpiZK1rxl10+ilE4rohLyZjda/Fcw
fpQjitMq2QAZquFl6mV3z60ZchicbRdGwEaPIzgizhQgMIPIzn0YbwqSslg6PlgxPO/Ii93O/PFo
t/M9zVTZJT1V0fjs4vPJj9TxgIEpUC0S7Zgs3dZtZvs0LNddPVB46NkwgcBDTRT3pvETmP8j5OPC
JneFoWVrkabyghuBoLcKOPPRPapArQp6TsBRldBG9121mNq8bmxxgueu/xE2FAUUNOGbM8tgkZAO
87f58+oyL80otmsiWrN2ujkuc6Q0wm1/pIfHgNEKiTx+dQKXHpjGkiB0dpvWk/5cWaBerAUJBH7S
kITzf08AXgYg6MioLZ31JE5tyZd+5qUfWh3aJ4dNsumqFQTCeLKfG86uULJlJzAirr+cYXJKSrnR
whomEuywOW+BZ2ZZgBMej9pvx14oMDRczbzPxia6RIss0HObMHEuTtJ9YCDLJrlEtiEsq75MryTq
vURDwoKpjBdQEnBnEGvuZtonijUlBNlUM4KYh3Pj1+zuqHcIH9lcTbHPCOqghu4FVifCd0diiKO0
UZCrFl62lXgg2fcZxqDrpVevTSkU929C66wwBt04Fym4Tt/1ZwOQeImYn3MAdFYTDZTc3/VNxLQm
kH65QVWn8MRx1lKIU22VK7y1ua421bgJsnv3lgcapbQ+WWyMASyGUHoAFoC155+B+XaD1DDOzEcV
G2aL1rspYaaWuZmkdD35opSDO9a+78yzMAU2NFPVvZbepQazWvLQgmWVhGC1bcSJmIRXOSslXE9V
F/DBaeux4nlUd2bV4ac8oXtF9k9Ag6sqw3GQWHZDmQEEIoyL5d+qa1wEZryyhe7j409p/ABGbF80
AzF0UnwjwcHIAtdEjcAVad3e+k6mPIYhr32RI/Mqa8RAMPuAx2yLHUYTfKltSPzdj9MpgYt4RZjD
PZmImbkXK3tHP0+Uq4jHH45M0WC1yFKKlksdBH6gdHrdmTlotrg+YhZaYAxJOQRURqHnfZ6yhM9I
D7W82ab8vnoQSe3zNhMCwFdXv6BFabShU1NrMmJkqYZZIbK08WJVgsyfQakrQUztVwSfnmmRkPf3
1BFpRBCF4IfERWuh40CZzFE9FVlkfwqlCm43xu4QPdtnAdMdETc1cs5uiO/y1RtD1yEE9+7KpIpw
SwO4ZnohnhNs1KYsgtLd0VJRadiE/JeBKG1LxOGEu+FnahjdfCLFkMpIwcqmj8vlXzDN4HE7WLhO
B7hP/IACPqDrniC/vvR0rBIzjj30JbKaA1C2JeZJjIx74r6Jj14jx+4yIRKKmRYY4QbhLioTjELA
yxjjATe5XuFHXThe0Piytr7FPLOH95VTnoFzYHqd8OAQa5mjW38RJIC2JbHq2LKCJKMwJ7zMrMr3
XoPhLOkLuDFhLofS+NM8+XlZBKANxw2nEwg+mvhHS1bdBkcrKDk6ee4ZJIevG0RDEcp+5kqqxopF
MWheysWw6xsIP0BgS9WEIxD2gVK1DAc9Sn81y9eou3xoOQ5RgnHCXoCtJFwv2CMgtU9XxKR3q7Qd
LVoqC0JIlb1gvRPvsYN6rgjpqao6FShKPm15ibMKh8wNyes7Mqu/5/R+vpsEmwHbZ2mROk6aeWU1
njBK/gMA+1LwsE+KcoBHzrOGQhQ41IZR4idlDwzKQvE6M33CpH7eScxgqT3qGdi8LK9EadspBRqJ
7jLjtwQaYLjHybMf6z1HsIx2pFc+vUvkdf6v2XGYIssHQeCMVMHoa1aCYHGDnjpX6GussTC7hvHS
TBnIpFbZslBHFa0iMpGINWEM5Y4d0hb6TVUBNNeHPTH5sREac8kRo1XSCOewQxlZU5V2nmJ62Jy2
SJlFYXWYy/dtMHP89H8hdFf6JffxrvsTzxm0uI3JoNqrBJRQlfDW5AjK7GlLALmiR8bCpASmWZuc
XnSRdMQ5Njak46EMTyfLe+m+JxdU6RZ/1Rat7NjM9JL009OJ7GTZFwA2QazOr6B9tM+HZFjAQB+x
6e2X28ZGEDhh4SxOiKiVAfxzpRfRuydCmj8ILDf87TWDU/OGn3JOgb1lL71O9an+BbDBFVWd4ZQE
weVV9EZAaUiVeAaeWx4e0/1hWUs2VrJsrLx1NJSeabUVJa4Pxnp48S+TnROjMeh5C8A4T7adycAN
Op07ZJpO2ciBKdf+gohtItT8eB+te7bJk/I7pFeGJUHt3+3X9yaPpyUnyduW4C/DNWgxkFuH3woP
Jbh7PsZ0wGRGGnnf8FI+/cE/i6FB6FCDN0shf7ZLmOrAGOQsk4dmCpGyj8lJMljxU2cNkyM5djZo
xOS0Tn3iDBg8u3MBoGj5SciCL+VgNVh4MRlHxxtmFtBTV9UEqdTQev+wlnunmycF+7mtk1EBrkV2
U+g05lsVBIy5aiSYxgB/ys9krEAjqAKvxsu366fmVXRpfaZa/J8JPW3OVc/S9wtwnlAd7ovomiSB
rBFlapu2PhSkawh4revqo3lNGvlXswZC8yxK0I+r2k48w17DjuUy45XWUpsQ/mo8vyD4ZztNGZ+t
1ijyRFtZY2m9L2g9F+tqj5uYn+Q1NVdZbYhILk6cg2TKBIiJeDG6bVSXNau/5PB+lhe1ygMpsD14
LQfsnk/WgwqYHF2Cf54JdAz0YXGgd14QANjRIUdmMtlWi/UNMEzWUtyOASynBSo85Yw//9Bn5Gy3
c44t0TZXO7EjnmAmB1Gx94ivuciCxHIpdihPniRFDtDBOZD0DmUR6J72R86GB1zlNmC7G7S+8NaU
p6ZZuaefUqWbKsPuNef8AIIQEJevrj96bcwkXOhT4ilQY6eAztRtMtLsek8FtEv9BkIzGvBijIQV
NSTaEloDVtQKV2zuPoj9wADp1mL8Zs+4KRu1T1K/ZRxe5iEXbUT6HO8qd9iobCUXQ5SqIWnn+LPi
gg1xbN1Ju9vH+Mr7+4V2VGKsh3AbZ60h66NhE3na6bOfDqqEMIBxs//VDxXwPLXT+DGFn+VB5Zgf
7o4N6eP1ThJ7jJNkFKfF1l773yLsirBlJAUU9sqzTj0wuGX9sNsCTAVc3EM51+ZjbbxyojCKldjG
AGaRfAmv+FbJbfvLiwunes912gWlVv4EkEEutbQ4WYwcD+THIA3ltKWwEwVzylkl049UQpswf1KD
elEiR6xOZvW+AcHkVKi7it/sGMRvOsl+/GMcx/vDigfpNzMybqeiosFgchEpCeDoR7nBpAmbHE8x
ZJj8Y+BH//YJ32noc5yoy5Wggf2SypdqT0Ny1gwjtKrd/izo3dRxMCW+M6GYiSc/bCujAnIFFPta
sDCQhpoJf2L5h1CYWqCOoIC24BlwWhmhuvI1hZnb1D8MksA0hJ88KSAEzfcvioUQw3T+5znWPg7a
81aY2dPyfsINOQNhpHsedyw9azrrlNrNOdkfuSAQKcfgqG2+xbU8tJVYtMi2oxDIFo0UyDw1guXN
2xL197yWuxY+CVUETfXenQpRvepZTCMD3F6F+McoNejSzgQGD67R4CVZU0tSf1Uxhay0TSzswfhI
yxdRMlIRRB1BsjWVwNbA7mWnKPi5o/eEK73MInBHhDmm6/YZT4/2d5DEXbRWTs2kiak9SxCI7OJv
bTqtKXn9tDJg9K71ibs2Kg39mWg0iCbowrlLa9FyxYw7uEnIl9mTbrNfpnUQioxdPUSp8wYLaoxk
aejrMp43l83rlKKDML0rbwjbuHp1RuN/uigjRE9hEniPsDVHiTip9cHHPJV6QUDkxhJg0eZNdXVr
axRDKJCwSAh+gUUQFuaFgfcH/8tFBAk5iZutybDu99dBBfHscisFojUW6c+3e75marMh3en6hVvo
seacq6HE1UJQT6C9/nIanSRJLyglmclpwBIlcw19/U4aaiVhh8mLU/zSrGxbepofel5rDeXMDthD
ZBeMD4ExKMrbfTCdPVvbTJPo5UoO3WIQbzztjTJf4sqJyL2rfpmevVP4gXBk0P19Kv7uTzwm72r3
3ySZLLo0GULjU94fq+PgTGzfMDedg8qgS9f+CVJF5E13mQRDZnDQ602Yfy0cR6D+5J3Gy+uZ3krF
1rjN6DCnmWWsPWzJwRRWBCeryhKfncFcytsSH5Ets+9FCEa0gyhv4X/XbqtPQzHdZUNcyc7Ofn4d
tDCqWyuIeFOu4vxKWsmCnF9z9Wd8llz9ESO3lva+ZE+Wegu5t55BQFEw4JLGClEXL5SNFL0OR2SM
UOAieYSQJJ+BQWmBynlk3mQDhke8c+avpJ9ZpJvLRe9kSfavv2e9XG361NMO/OLV/E72o+sjmzG3
0MiUagJ9nuryFlVQviCaQYh5me3sq8YmIeas3572XTQenLhiZpaSZ9uMTgsZP4rid5XMHO4ytWUt
A2fcothGC+2bnkZzsozVSOWSz/pKk1MINw/9LPhSWk2L2BkMyDNlaZvfPpnn29DYNPBQ7h/uYYS0
N6eDdNauX2b67C9g+ImiJdMt97fDTXVlErYHsY2DvzLcZMYJMVQcGx1z4/oup1wGg1OyQETiWygQ
c6etgSvOFXOzApwxZ9T0vkMaRDOL19qWlXgBE0YK2WAlvK/78qH1b7gguLnS0nnXDWqWGLZceoDo
L2Ce+gWjrsaay2TbpgQiMEx8MWqy8QSe8pmMqzx8st+g4r5iDfjRicSywN5CzWKh2POU0ekL7rBL
CXWlRVBM2yqzuplEdrxg8fLORbMI2oZ3c6cav4Y5ASj1le4KtrCjgY0NzU+LmFQhIm9GsliJNV5t
0xdXzRUxbc/MiAlepHvOkkDQJw6J8BRUD/wjYfItaWfhKQRU2VuI2dlO7qLGAY5qborPG047Stiq
va3ei8CyrykZqPlOK/bzNSsEObMRaNp/FqWICuGayMKPB1pYocHXD/yg8Lkqi3XzUIG8J08NlkIl
rOkLY0BvuZZnxuASMRnskyI3N3oQJUm2hCqIp9uK8T8GPz6Zhn11H9oZedZ9qb1OYi68pP5nZCxp
k5JsUHWyyKXqGiZLo+pXsHHXwX2UF8emWTdU/8k1f+xxJmNSlQOq22IvDRYqEWPZ7F8XGNekOyZ/
a8Ow8OcFqG6NkjU47DurnFrq+GTlt9T3Pjhi/sLT4wZGAllk7OuMyeXYRHNPgaPLoKtZjXa4PIr+
dHzwcP5g2MdU+wgOX/V61U8IxuwKDvI3HkCD2h5dwVUkkhNYVAmEOo6yGZDpHfjzQ9lclIeN4dlr
30BQaP+WGeIk78Roj49iKflnpVytUAZiVFM8oeJNckecUYr6TME7tN4KuZeSRzL42Nb5wBf9Wb/A
SmQw6wujmjz0TMo2MHt38GWSoIMq1kSCePh5TNQkFmcMzXfhSgxs+ENydcgqL5vKXXMQ+1fsUv0B
bEdsU6HzQu3iGG4C6F+JD4tsMyY41266Ah1QqCQi2YTrL4mLcAeiWgKxcdFcHdM5ZVr0oyrWlSZ7
Rgzm9c7D6+cHjZPF2Y+FrI9RurEQe/0CXPv8RgBAGWjFi8WOmdLvrdmFpq5SsEPAkuqZ94i1h4P+
URkNRXE4oXqVRvwor3tUTg3zJXzTlBjkoNQ1rpw0MXItdMd7tThTDpErApUDMG+lhf3UWwN7J2YW
AIdGqGw3yyQ+NyXefbxq/Jbe2IQP5T2bYnVpxmeOfep4tKBuXWQMA/VM4zYgLtlDd4BB8yBG4rwF
NnC47biEw3bPR4N1spzpyW8H72k5+fcU3ElG4s7c2OOHrQtmRRQjGP8qfSqbT9eNx++n0mLrGxG7
b/JrrvZbr2Xse9HXBBPBYUsE5IqAx7x1GlFEPHMynVXN74jirDUa+DSIwVP11Yctd16qFuMKHixL
V/OCDwzIVT1CzzBU+EXCmdGOHcLS4qENmA+9nmwknjaT1h6XvnVfw4bFHvPOVCsFgXVFEj1u1AjV
kCytMMHsp5XQRkhMzkkioMjD89MFtl08XR4lL2KBo+Sm4tc0iWyYr5lI3rcax9yDqqdndwL4yUwp
xTtgX1emJaFdIGXfyUBSGbK92j7wTmvUKg3cvmrUU0u9GgzAlArS6eHMlq9ZW5AL30XPdKcoBfZz
UyH612yHFV2r8n1KogO4w0VsZERJZDtl9NlA03xKccmKqfms78r0DMrWPDts+ib+qNqSWY/ojRNV
SxjkT/Yo8y/F+m5D9yxG1OneQOoyHM8H3nLg7CerptbyD7sJjBH1bteagxRozCxWS4Q3SOP/lovR
NVjiCSq2NJYxfstz0NlQOB9LhxvhkyWNZtkwyFm+8mX3b/8vVjtUukW1IIDPWXXLzARs68BCxohC
zEipeWUTYiNoJrPYW5YGEoBJGFmCDah1zL5X/ebZMWWweCC7LDQD58eqP2x0XQPJP6OZ3prz84XH
6g6t+LCxFkWXRd6JoRIWl8R5zSD/NMm93XT4XB+WlH18voWXVVMq1Vt8ZQJE+/SUdDXTDKNk1lZX
vE0sKfsG/FldEzNubl2sFWTj9eL4yTpsfunIrWZ1HYrsNHM7/Ak3Kl2E5Q7whKKJiod19w0gCypC
2EP32nFOakAdpolNc+l+kKWLeQLRoERdPYyCuq3JAZnmcXWYXD/mOwe7e2XmxXxwBDm9unnF2++u
viPyksDe/Cb4+mdJ0Fg3UanEonhPej/w3gQGLi9d6udogbAy8wYx3JaVOedjQDX0e7WArrTmBxg9
nkn6X9aLdHond7zqpJ2UyfdgEk/y4xqrLx6bAgKCZHMHpNV6kcGrYq732g+wH8DXVu+EgXXsgLHH
90YA/Vi4yPPJBje50AYfWOgEy9NAIQ+vjpPEro2Xh09N63B2UZQtfKtNf6houyn/11JlVQ0GajZ1
TUDF0cVIT56aOUVyBC8zWwr8POB4n2Q+UUjjMzX6vI4FZcgIC7/KqmgAkB7ywJxRaxUzHS4pNjMV
whdXA7+kpfl9eIv82EwykGByG8hwvIjvHZQ2LNaVJnXX9env+Jjcs9J5In9Umm4ttlkMovUTg+g4
OppX3rBep6PtGyoWo20323S+kDecsex9Gx1+lU6bZDgiyJHjJqSN3hifBHj9hMdjqg1tYnPeZ953
V83eu5q53S0IyHig3H/qGaRCsfrstbSaEckRUL7W4nUHBrlHmxTe/lnwWTjgGtD9qzlH/oZpc9MR
UPl2PmCH+ApJDayZcOel61hkt9Dk17dJDB/mlZDejLHE4vhlFNQ2TPRiPZUW+nacD7nkCr5diR3i
c9+zVbF9rqa/WN40Ujrr1jP0z1cVlYZsw/Ql7YwFmpMNc2yBp0dFGzJneG9ivkKiaPPQcFO7B2At
cAQmNsipXixI/R7jGoqLSm4Zoyxo4WC14dCxHC6SyJf91ojP4e9U3rmF5n19C2nFL5adLVGqAWK7
EGC9lM2kxklPcaO8knMSqPxfCwYCapH4Hl+r0E4unAGAJKX/L2/SvCt1AG7vDEgoY7r9DdtGHaC7
ttSESDD08laT0VJFMkG9xYBV2Tet1O7nd4kddchYz1udDstbgzPN0Mc1vh0fr7/E6+Eos8t79zul
4TNcsQqs+OgImUGrySeyFUvaCUM03PINaUukp0XFYTq3HFyPoY2+MeGhsxwe2904T62hZMgQALtY
QZORCLlvKBjZKDnFYYIl8dB1jHDFins1LGuVLCyt96OH9TqkK/adBUUtWz+ESNJd4WgOzT4TNove
8EwhXATSvMzfIEwC6taz1KxYc3Lnw5oGMM0o9BxSvqdnWt0PYd2o7gJQeaHDe8qzeg4xadNvHGDo
SmKG2Wwe5buNCQayUioAgzgbN1YVFUtOyxnGc35cw/cJ20ONuruGnuUVWKIYsPxa8m7alcMiDG/3
e5UtM6LJyHptjq4PTvW8NNPeHwRr1RuF8IuvuzkMWAGSs9EfAi5B9iG7vmffophaP3UrTG/YFa8z
IG4JG8S6B4jzMkyMHZbWXRIn8qLf8vOYdF73GLTaLiFlIiaaiW9VhIkwH1uu2HQQaWsOYXlWksWM
gMPEV8kmMxH2hqUjMMQ9wCxXQDa58Ej5U5745m3mxfFajIAcU3DKnIoGV6Mv14OmjdHO316/593B
/jhjC9Eiwfx9uAhLerm+MejjKKg5WxLJoq1qFjH3hRCkk4T4uKjKXcsyykw2/pu5mFhRh0MwqzoZ
IZiM3Nr+LmotwBAv+Nu+/rrW7rUtgyOQV6XTXbB88S+EOXKoPoEjy19raJRBziG0XLTddL/udmGf
qfXcjZ6f/LuklXzb1hd9f58N7p+hDAMfW+Vaa/GGe7RBxwi9d3V61sPoVz5q5AFVYaXRs0W/at5Y
ZtMFEgtH5wTmhj6Mkgb/a0MEDjCdYx5CrJBmCNnJnhS7CetxugANXenvLfuitgz+HK2ARuD6pvey
Mgmvg5ldBDVacAm+pVPmgV6R99DiWbiUpvhED2UOaYFdEx9MYGY6JfzYkNh18APY9Tsu14whLvwN
YOQSutz2ETGtuHmLBhSN2Nxg3KBicgftaK7jJrgoIxPDDGHy3nk2v+YbVNPcFu/P5cc7VHHNuiR7
2DUtpp4xAdrFsT8Hp2pcva9TdLw+2/aSlg+bMlzBo18P/Hmj37tIKlbk8HegQ50wOq4pwuzGUXc7
6z/+sAqAqbwH9Lq/3EvWa/7UxsrIjGnVx2g5gjqJehGILdhi+rKR5/X5MlL65Ksy9usGE4R74BD4
82ViCA8z2KO/I78T2DPj0NeoinlBS76ULJw9RsiJJAo+emhZ4huEuNKr03qiI87ylfsz4ZfN0ES4
z2pusPsnTvekQuTIQkBPkTtJISXsaRxa8eZuJv/NTSwhKyQoDGCJ+F009W+WQzERVXU18m5QdDHr
BXKAlEawW4js8l+A4z2gvg28RawzX1F3cGEpzWIFekzAqAV1d3K2kAL1tCmbclXkMYPcXi4ZQ+98
mnC+VEMy78LYhx13EvRnnG0PY+/t71M1vAJsPJxJ407PcJmpYzRI4b+hhGDVrGMPONTkZesm+5ot
Ki4rdVKQ499k9ymRour88fED/5kEki5l+amP6tWOqACZ0Rrc/B55Yb2qyUlG0G3JjP/eZPPOLrXY
qmywA+Z3w3uj7yRGkPXCOyUs5NFBoSvTrKZ4uuK7NC99mCVcwjPXoCYpBZnzx54qUquAY0Kwjrak
NUlQ4o1/IyXJ3BhAHdxaP1uMVfQbEfEIRK7Ikw4X1Nnpf/K30VmUcOWigK1WHK9+qa8mRlmdT/Bq
A8Sap3CgaoGDUMs2ZbHFgRFKHGTwBFcGnJLF6VcuXH7pefNx40ubASZPrHirCAlhFpoVNtLrTe6x
WNYDjrieneix03+0Deq1VsXJ5JzQ5mt87KFYO0KzcaTRRO+S9vfada0PocaK1eGevoneH/mNerpn
vpejT08Atwge3/hiaP/MP+gmDhyQjCL+2KKQGRVk0BVjnrdOYEIBUdUs9+O8Z5rn8XQq7tdw61WL
SS6im2IL/8lXbWpEpou4Z7zMzyUhZZh8U1S78oZJRF0Z8DzO6tfGjwEgCCCuHiAGAoc4MSyxtsbO
XV0mcuPZKSGQUC5f2ETBk4P5U+6NzyH6yCNEYOLEF2Y4NMG13dnt8qhalGcW8gIM9KOyUmde42pR
GM+37MWvmvA2BsrfG0auhMXi5h/SR1L6QADvOFO0dUuFjKmDkPOr8b6OAmq30ZtfcQei/XJoXx8I
gOulQ6hxAo+GjhGMo7oERm5kkRZWuLWKJcEUp2rVaKR9m1MW4ZqnNYv6CFeaHunPtAuHCHVd1HGN
yxiMtGvgafg3UeKbX9weTIpHtkjwbRU2FfqVvdT8+X1bOxV1byCMs+qTFBbs9mTk9mtly1AHh3hm
UItqUBCbJnHqXbDec2Cj1Rso/vnVg/kXN5wehJuzo/skOkr+T/GWssrWEM9JxLIP/dbo8jYQigDo
Y7AiMCmJT63xyyLIpbUv4Xjwl074Fg+GIMnbdxYCmb7kvrhVrjTqDDyBNqBs6EosBDM3djiDsWwT
MnjsP4jkB6KJqumGyrhSE07ZBrWBkvqYiV2uiZVu0171/eemaAueyzyqFFmXyDUYPBz73vavKQ9o
2kNOGKCRaNm2224XiLqj2ROm6LVUDgOYiku28NsLv1ZoZYHTPkIjsYJay1cLtQr8F2GNYMNF6KzC
2xDLbeftYKgiDfzwsFoousfEVo+7LKgwGS5BuYjTGdjBgOuiNE5pBExX/I2OnE3d8ELefIVGjzRX
Pl9X9vKPQmEC+jVDotktc9o8vFV5rm++24CPiBaL8j+fSnZviJ/BVcOAruUGDL6vOj8MjsNw2seH
kn2GoUx6OzrNOGH7Xjek7V6dbZQQEhQNYehpAGql0B8/gI/gSZ1frb4ra2p2ku9HFMIoAnbfkLRa
C30AOkMKwkcafzECZKyNG7BYOwBYknr7oja4d+ys54/uRWSgjmq0ti69QAIIcJii80F+o8IE5uVf
XenhGF5gqLuvFwKvWKXew/NHAr+kJGNhsai/oD0cUVMfTEcl1Ii+C4m1nmc44rdhvt3l1H/Z5Tgo
/RaWAnnG/Qj741ya+yKsBkvkJ8o0rHe8dUA88wS2YtCXG3XF5Vk7fpZyKu40Vcrl89tb+QO+oKUE
LBHonRCPcETxErFmQNzLVFe4drqyyF4XKAuQdO5WD4AAvRlrgG1cD7W2ZpqAZwZ6m81Bm1GrZUXO
0yOgmwe6ZPFd/FBgZyI6Sgm2l4zeHiozhyzKAcfb79qQ0ZgqZubzDKkhYI0U8ZxQaknOYLrj50ui
iyslbhfbVAqMWOglPoJpGL7uxDOjLX3DLsGwCr8j9h9EJrVwFzAskjBmjsH8pCvlBOaCCDFp8e3K
GxRvORn810A4Z+q9g5i/T/1KXczXSOjN4S1/G03HrdHbomoRaJc7EfsAbOHMvwh8+B8pM+9Tx11P
+QxU2WnulbJeqLP4d85wCyJeDcpoxir3fL6K+6J0vBh5t+ejcb4BoUc040JJruvA1ww3urtDMCzz
ippuYJTEWft72HeYr0LzvEnNQDvwLeroPHlb1OHugBFsnSQpN9j1nC4szWCd7ssDSqEQPykc82cS
X9ZI/1x7y6qMRiXHUzWbeyc5PBjLf0GOLI8Akrl3vbECLZdLWGriKRcusVrXda/zsYB3udU/hW35
cNShrLSwbgTemOFPbTN0DoTtCoTI1j1ICsQ4scVcucSOpSbWodCll61Ugu5R+Ci4+Jt48Slk6fk1
FVlzSjqrEirtaBqp71gzo5OEkQ4URF+gr5lZftpe4H5lmSLLwhgzLL25dofqL3uzfek+NOVgdQNL
psYkwJCoBudm0R85bYY+GeJrNkFvnOhJfT0sXFYqeUt/cwEfVJDo0iQHdxSPph8QWN4dHY2stzJJ
jMOqqzJCzKmFLPEdu8WeqUUp3QP3nWgVxmgwWcrEu1Ef/XaR9T/WwINBZoMbCJJrp8UMHRccUDjr
o45/mUVeqw5k91dEOo2ettxinRUtUEVCDbwu7Tsg7RcagSyPtn92C7U8HzlgEoBZaT5EvSoSYN3P
yudFwok2ys8vfSYZl+0OiDqucE4+mM6ZuQPWU4GRUns157nDVJ+s8sEjB5dyv/IuzOlqak/TJs9b
bnhDux4hFgAAGH7mjWNjq5aD/ew6WyNDcuS+MJ0MZcMBA9vY8xNsCt5wIGufs7fyoTvVoEu5HtDW
7moFZk7BZU2o6MLAGfxQjFoKXB0tIqGJ264R2PJlgyxnEzFyhfHlxplj9iC5P0SiGcokdeqIIbOK
ObhbtLECLznNtdsdPbXTYhrtWK926njvg+UlNQ4m/oUBcEidynE/ksR7SpZ4I9DGe/ujuh6Fl/tQ
M5Bc9vK2dz1zPBeA2WnzpUj5CP2Tp+ltBTv5yrzKxNPZNuPjPITFEUw+2poRkfzWf1Roj8cBy6sS
e9o0mfHP191A9m9gYg9UONjAFrW2/qmLGxOEgmjQgqo+IVsXU3nDLGRVAKagvB1ClKvQYDDLIRlo
rgVYxI6xnuKs+yKbb2KAedJol5RMOFs42dZ6Gn/OIZyIz2QGnDtDUewQukWVS15eoWK0oWvmejV5
aWO/gXfCqzsiLfIXvLsvWu/pVUAIXmKEn4PutFI7iABALIJ7RsKJwGJuuJkLbI4UdvaUEAnjob3g
uQj8ytxOlbZnFJg4s7v9S7XqGyNprVZm9vZdFDqsRqCOHcuuCCSzwD8rCqnomE+SQ319m/6JdQT8
RMWbCZhcXbUTupLWPnKYB5X0Ky1v03QYMk4vprd/ps4tiUYqSJFSyghKVlX4qFYRQwyNkm/Wvjg0
3IfjY4kSvSj4BspoV8wDE5ARCBPtH6gVuP3k2P0+NGLtbA7UmCzFnsyqjfM5HCArc+W0mIzBDpG9
/Iz5gxKC3j4h67kIOpYGC7io++j9l7IpWN4l5NAFq8yxVXUzdROEGEuPAVm44df7kihK0jqyLfCi
Eb8qGaMOlBw0hOqJguEg9BO04iA7J+WeLnqm0HScmfi7FdOyywgnZh9TEO0TVWYsJkabh8dEPoVk
qn0rSG/d9SVc9zK/aAoCJm73qRtdk/lJT4vhJubCOcKycFcOfHBh6//E/iH9+MPe56+7osbF1vnM
z+GA1Qd8w3HM+x1/hIZQmC05QBbz/qlnx18wM/VHU9e5l9DHJoES1RyfD3b5VknIsPa1k4cQ0ynh
kx4sM8KgyL5GIZPzB3UPleL/WCMzkcm0B6SLkzdpBjbzxEGHbhNAsgmx0keBxbxIwAAWsodIf9Uz
x05BrI1jkjPsQZMEFa/ZD//neIE2mPGWXZc4P/gmj814Uuwh/IdW1z9bcM9IRdeWJVpkfw+qpT6w
ibiFSs471pdowxrwEtOIBlmTnRLYeBe7D97wKSyO+Y0EerBEz0JdvzDFVEiXLxUmg5HWCVWGLa/X
/UWr3Tf0EwNvKLR0JHuSkoQar+AoXrdnq0ah5gMJmUJGlrHqk3q6RvAPYwZVcJZ6oN3U7ZA2zX9Q
eGGT80TwgDdNuawvnLkpcIN8AtmsEDevuVCtkI1nYQWQ7mPRSJW+F+Ad+3RgZL00cDf5F3KMmS7J
ybPRMz/fOoQNnEJqVbgZzhwdgsr/VnrEoF+ikOvMbxmhjSiAP373vQVjhoyLT2+YDofyir8fF0pa
RFWtE6J3Yn+SUk34BtO5gX4/OXG3UVaGKqO2lrgdYMiaSRhTQNEMXKPZgpxQ0bpPYdR4sI0ai30U
uG+/NPLnBV15g7c9ou6KtBVT2oyrFVAAvvjsnHeytsPTY5RdbEctl8xcojF9rvyOea1P1Vcf8lWB
zfXJA5epcj2OSByi01qtGua7rE4OyxZEEuQu4DX5IQBDtuw3hlvHFC9LKyfGgteGB3rbZyqWPqBz
WhbixHS1GURvi9bB/XaevKKI5vlyI14nYJux4w+jpTTx/RTPeqJaV219aWObmn6uug1mSVkfhgDV
0i8Nt25z62hWFFLo4Az41S94hPTvS1ZQsKsThY67zuwqD1a9lCEdjgxYL1mwELnBF9BBgunW8i5g
qe+ElaJLsTsYREL/m1b2tlJAZOej6u59fXuZxh5GjT6LKxnwvOBVcImNP+6i7GLjRZQ9lazs/9Zt
mZV+Vv7KUuHoc6BNVh+ObRmP8rcVuGSJTcT1QFV9MCR9LvUGBOXB2/ZXCaY/P8ZCRBpwM5ZCqLFY
A+Dde8Gxd6ij4q+HuSEk8cp2tOGUU5tHBsi/06sxNfk5e61m+jqohEVYManXjrDEuiJpvwtGEmUk
5Jhg5Vy9+9nXctYKXivpSFBFR7D16X7je9vpmJt4IAP6LVF2saoFkXUAYQdWVT+9vO0Rvu0wRGf+
Va6yTQo3UFF/uVNavPDkNX4ZXV1RWczMGtF4cqJbqACl6I1Ja9tvDW3blUccAt+XHj6BBz2aEt9N
pYuSGCcGAj7bkEKGi2nACFrXt1nnZ6q1u2v9UQemZEIeOFxF+ick2VcKPChJ2g1HBW0JS9hQaEJw
VVA81P74Nj25UrTmEc56+emF4UR4SkHb6h+89aFPXrJ7epVse0pVRRlJCSfy+eMJpHn7yV2gCmS5
4YZONp79q1/OXknMVD93K43WfzJXLmKRIrrS9nOcyCS7BpV9YCHKmK5/gwIRD/0hNLeyReDMwnmr
ijlVX3oNBGbWiN1NaAUHlZRj6CsNfr6iFBp7hNBrafe2joaF15ZjBMZkjRUZpCcXRa5UXJzMvvdA
1+VfbkW6Q+9M7Ecgi7SxIWdjBJdc/v2avrVHcf7KAF94dlUywgGIECpHMeBd1HOJ9IY+JIrLCFAx
aIEW1dEEBofiXiOfuGLvY+gko61h9pmDSnFVVmlCBO+gSqpQdS0BwrJT4y6YjR8p7V/dOrOB1u2D
6leNXYBaokKI9YU26Q3VXYtsFc4CCycYWJFWXhngS7kdYFs0Z+2338I5evlr3pbbcTJXvkwUc0B7
SFIrkJXaZUT97Ambz8eawMWei8gWZwjVNqAGlkNYeANOqZ+uAQ4N4DvfOVHHtwJKdRfVSrwxiNdV
L1TkJR+4C9n1XgPDRR9iO0CKauKaR9U0f1MDQoEnzgWzwTHUiPyI50kd6T6OBrAAt4Z0UOtszXS8
4BYHxVY4Wyzhfy4iejXfhF8B64FUABTRwqw18gSPUBugk6o96af3yVd4HPszOfJsxeVIh9RgjL17
XWzL4t57sTjblwoTn7YnGByeK+qYEZ+yMAG6Rtvw2o3ml75zvMzgVkwcm3Vg8utU4KFQm4rlYaa8
+FHqf/pyzT6Om+bqIZv5hqW8NH3mptrx4b2qiBoQ8Z4nmvjnFUiisARZd88amisR/3CWsMTU8MUZ
zHCKIqe3SYXQkggVMjE4HH+gPdPlNnQI77jBKRh7vd9gZFl/+MYuy5aihZRjlkGZtDyG6s4D+ms3
QCgDzWuQFwvW4bQsJOlh55cTUzteAQf7+5ZoBiAkk5SPabUdyiA5vEcnrdhUv9CsyJDLhV25Qqao
4KMdsAYae2X/t7ZGUyKENhg+VZ/F6JNlNfpmGg2P3ATreqTBHZwc8LL7P2UrcvX3sGc3yE47yj5P
4f+eRCLBwjjvxmFDj6tHzGlMvx93guwgWKAWyioGFngvcuTi3fkNfHP07oFciKJ3tvx2QmHgrTvH
OjBRW9TaCRDoJVgrDq2+lEHdeZf+1hiQNn+XPB6l0qRq7Xl/BejkkpMXbZX3xUTb9XPXKr3S381Z
Gm3vPN7kqDYew9c3s8PPC6/G6NaY63YET5YpfYY682e3cLRLYLJlKCC5v0SLSlxte/37Kb+OxlhQ
TTe/DNVA9lDFbb56Vl1dx9eQzmvs4hxpmk2EVVTk2w4hEwi30IVsIVufZzTDHlMAJzkpYwmGqzVo
c0phIVVdsYqcGCd3l5PKSspuDpbA3h54s1icJ0FF0v/KRzSWRDB9EvVNjUitFYBedhpGK99tvHHT
AYs6shde0MNSiFQgpMiRaPchVIquFksiFNEbzGSCVHU9jxAsM+cLdqlm9Yyx7yinnwFEXTRSv1mM
7R/JXinxFoDpB0I4epuQ4wY4IDuw5qPbqJVQILVKCxLU4SwvenPqC/GP0GTbwxAZHxXVQLB1mP+C
v4MJ4V0Xjm7O4p+1LFl6E8hnLKiKLg/pegQ2tBDs9M9WkbSYNgIb5WbOvwI1bb3KGtjtMCQrZjHZ
hM558I1hv/J8ercGvCJg8bVPgQeIx4RwgqM21Cn423Qxx328EGQs3vZZs/muekptja8jwjZensaF
s/koNv/E3aJtzJHE8S8xhHVnTTAcnuPKQZ5e9M7u47y5oF+p89hpQ2rkiWIn1vQnyZLc3bvYZAWS
RO2suGYamXP0jVtmOo5UolnKUivfVP+lm0TfHCIE1wC1p7SzwE3/+P3ynDqGXyoPQQcBq0qyCD9F
8Mtc4KJ1xMoOt2ZY3Ale86TwaJyeNmP2Pk/u/wZwf0B9MzZYt/TuRNIW/pJ1l3liaD3SJAYwPVRn
g816hN2iVOw45EZaySUyyEd2cAIxvf0ryWfC6GVnEddqw/uBqWc0iu4mM+B6VRC+9JEwUN7kODJN
9tQxvqLEEHb5wix0iw12Etwrz9BxFPfcrbWf/EjnrpoSjQaRLr7WvXIQqsKQkn2iBKT1H/gpx+4X
skBEMxH2giqkKsWDqPvzcTkx2YnJES2MefOGR1yUGYcqqzpFKTCYWVvX7dELZoQrXephBjbfm5SS
K5L8celWRwMXWOsRMtgVVjhOMI17iQG8ZebZZc7gNqv5PNO2hVdl7ZGGQsaL3ANynnpS3PvwHl3M
0l3H1ktc92LpzEcfIIeDHQNjzF58vFYvFshoTC8qspITtYkJXQG8FKSqtMp2SVth3N9TydCHIDH4
KUUn4EENEJrtWZwAJoYvhBN376BlkP5rD0W08F6oROicN0r613gbU/uaB30swgkqqFDBOjt0UFF4
MzPZI9oihPEoJ/ETZd/QHI6D1KOl8cHseXynwWXsvTwMkuiE/2L4h65NfsXq3dAqUMVlqPeMO4gB
2DsAXoWgYNf8+/t6COPE8pfGu2sdH4fRyLntM1cIZM4RzmTy86NQa1BJ+7xcY6GdR+pXfpND1hjo
48Y5CrzpsiLdgR6mVoX1/DzkxW+tg6vjzJ+7Nh2QopWIadtMznRLoTSe9XAN4R4VYGiarFEVUiJg
ohgKvBIZoYx6+e8uuk24zU1T//BZU3eeMucTIs5gM/RCnNFBHyZB4ib0t1M7ZdYtFYJ+vUiyFcb/
Pa8Qu0UtdhNvh+6jFa0TqozYDB/DhDrdMEj3o0bYCbfvURqcThVKPykSGb3+rqVR7DTiBZtauQ1u
P5AKSOM/zCV+gtJXhDz/OT3W+suPbOJqpMxyIW2XAON6fKI2QXoB8ko7jJgxpO/6f9Mh1DoBtZfV
pX5/rHjcp7HpX0JaP0kZCK9A986M/VG/v7VhIVPVv1ynEcbZTQUFQBG0V8B294siPw0Ohx93500k
iQqU3+08Z7DiEiQH14Ni49lBXgjbOlo8RpwWV4WAvOUYBeuA2GVULaqxwDnCMUXpnMsDbUSjnjJi
GRvLTjIsLdwKTZrUkaE0IukQY17BxaLoPtGDqIKwOC2VjlbbakCibYVlWXut4RzU4UTgq4uv6X1w
zwNwVFx1GYR9Kmb2RFXQe/Q7THM6DY0cVLynH99bNt9cLJMwb1HJf7IHDylPIP9795k5JfmLGT7l
WQL+sLBxtJlofEJcak/5L3T5awHJQSQj4xpChQ6T7BAgg7DdWFL+vHncmXXMxNLAOEz8v69YHmYC
Zh9BQNATOOYVeNKlRwjtH+CO+o1nYUA6ZYHRAFjwkG6q2jPCUS6FmHcUVR0lsMlXvztwATDCnYud
CuuoB5kEwTL0P7CqRpZU3XxLd350XNwb9YkBLmfLmekUHgR+QFL9JCjmnp5E+3zve0x7ghMoWDOg
Cg242Wtg9S1xSkBYFxyXCwTJ9mTuM22UIn4p2zwyX2S54+NMhmX5HtmoNipYAerYjDngNit9gDZS
DZUaPGrHrsTdgL/J0SubCcFedLuW8h1j93XdYhHvBma8DRnHNRx6Jz8u+Zoxl5lQKC0Z0tFFjvTa
jtS7IE3gtSTZ4FosT20DBreqiwuLaR0sj/OuwTtVKkBxVi5qIYIO5vlDXS3c5Wm+RejUGecc3K3l
CtlMFlAbZP+ZHTGByz2+F4LKDrbbv9KItBClNZqMkknVmkIVgnL2MpxoJOyoYk85wQamYOEQ0p7M
4T3Lv2N6N1kTU3xXaYwNvULUIrC88xOwYrYc4EG7eTAUc+i1/i9Ti7kcPDNPfxJO/NUeRXKLCmN9
8HoFY/mrvYJmbES9BV1uhgNPRvcfq/Vbfnl+3YZnp1A/vnUeJkX7lap4AA1ObJiC0SvhMNsklCQn
HXA8pem6ggLJoTNcpRtnKPgFa8n2q9dcIDCt7GA/L2/oLz6mqaShixwaImGPxxEo4K/yEjPg8pxK
N/+y+6wbRsHpvTvP26SwJAqvmwLDgEd4PhnXviVmSYXaeQrduajHFSguvmdtA+ioWLlk+RLcNOYl
Tew63AXq0LqR8IIZJ7pcdZQS+zj7FWvi5cd7XN3RVZRpb2rpv8fdwfNy6R4fkbpaUjYFzn+dSllv
YAgf7THc2jS3kkHEwJZk2YaeLVYIsxilHKs4nFMz/0tGQDeaAPEff5zd3UmKvK5CLq47cGgntkLX
cFsRqRp1lJSmocsT4nJ0sYHEG9wr992qxY87xxWwdAbtjaVDvrTS/E0g+UNPAI++5z3dETYz7zpX
JOwrRMmVRay+kl7X8yjhxETK+mPuZKthOkjcWi5pJFnQkMkgiMfCM9Fvigdsu3BJeMOz+Irbvk7+
TWlPnTLOQrnaKVaAstx9QkcICKVFd6KXkrPsBIQw66iG8QE4HdqSvwKeeFNbEOwx0/u2ttbGdgsI
IitqJZKb/s5pLBKLpvgGKTb1oLBx6c8r6mJ4mUwcJfkGSrMtHqXy+k3hvT79kBSRMESrDKEUrZkm
wfG9SpFmzlcDzsYNaV4N9wTuvXwLhbYjSwG1OD5a8K0MZgg+uyBKad8LZLDqa5uhbbtpROl+mpdR
fsbCA83SW/3smGNFC7nMXr1mj4XOlGgbDh8qJq5wqAdllgFMygMHWr5EXcEN30hjW/Vo+DXTUWHg
dmDiWM7Wt4gcKaAua3OeFlCkRZPGnSJ3320fPI9xLYwCOBbeFeF3E+g53HlR4j/trYIOvOzG/qgA
n6u3rt92CBR4+JEZlUkyumUGW91WyBQx5w7U4mLq9JkRkGBKFmGt20myyNRAI4ABRKJ+jboEYnBX
uCZ8FLZQ/Dmnk36Xs54mghzJ8iJ6uRj2U4DEeQlxVTRKbpBrwUOuBO1YvVqmQmpmiXjo74ouWt/G
ODEgVh727t4Gm2RL5YC+6Y7hjR8s10nn894lvyJxnDLC3l58i2a10YdmOsEQpmNfEUUKwlVBhGrp
0QUyfmLqDYMO3Jv/27MPUoV0v4bedG00qchBZV9rhKqaUxoxnLKs3B+iV/S4mXW3vtC+LqSIO5uV
je5UAT7sQOXeDFhwN/SFwWdL9jBlaDsyRAWOmC8AFVJ7ydqxYUseEvxA5kTGwgfmED0m2m7xKbsR
5e3cvdKaPrRxwJ+0M64cFVdiTaEVPO7AsgxuhoQCfS02v7xmOyYxudqRGwh+FnStgGqYcgiGZklV
wczfQfkcJCdJ4qCxIVmY9h8YH8dyuBQXueegq+9IHNS4/28Kemq+3Iu7a1i+Wyqh2MRg4t4y7XcF
TRZJGo4wWBppTFdd58r56Lq3DZaSBi5UWapA7pEKsPeLzgWtHVc/c/HRamfg/sR4YpeE2+5C3lGY
rAwqZZigqxH3Syiy7qLoVtMXBzQB79t0UvdAeX7BGCIf7u37Ad+XwthieU2dvePlK+YeUFrmzelz
0ZWLLnU7HpFdb1VVLknNQIppc79WMY2rqX8HNtgh/AQI+acIn8W5mJoM5HKMQ+4I0M+gjtfgyJax
BRl34VYMLRf5jxC9ZEcew8mvUukow9a/vYnFIl9qQZmMo0vqi5Ph+L4kO7DMfRWGSM1dT7cHkGKD
irm4BnmRJV2uEV3N4Shb285ynR3WABc61jCr9k9Ihh3lw2TnTCqbb1OCMxqC3aHWEY4EimIZDHjt
/zOZMYNdq0m0Ivv7j7hDZybxX5GGd60EMPv7TpffCjBCv5vCH7We4ARFrDOj9W0bCBOSw5YdQ0w+
2+ub2cAny/UGns37YakxbVhCHblGzGu4XI9RubCKvu74voa2mt/V5cUloeolG/L9lFE/SSyC0zIU
olAdgHmFDfuH9CXOmmaUa9ciSrtEgOmupErL1plFT34ZJsyctHWptotcITP8OJCK7QdfHKiolcGe
q0M4wQZheO7PVFE01yXUPX5IfIAQlwxcTpsu1g2rKdFpiIoqvxBCfZdlmFSzKD8jH7+JoyRlC/ZF
evaBlCw4bikXQF7JAsKs21zht+o1qFUsgYGeXJtS8lf60NFhZidDyqL44xdjkm/BkAjYjn1sYx+I
gmtzdCbhZhaZJeMGdRvVC0vP1jSOdAWhpG3ycXg69NB9tH2XStpTBc4P+zMN6pwh4WLNoafhHX1H
O0Rhra/GXIH2J4dKl8vLBifWAZ16kaXEuYLWo/gvRweEyhZOjHmEUPDzydgz+LKYebkOWeqIFTnq
Iv64Sor2EnnSao2YYwbeUSaGFLTkQlAq/2ynQq9YFGtbvlbTiDWS8SacsmOEjkpI0af5VojDgWII
oPwx4K4G8GrwjeirYkrbNw/j9I0+RG8qVtN4mcgL0PZhtLF+8inr11wxx/ju3DDCbQ8D+XEV/i21
NfJHmCuI101V20oKuVvndVuifpGPICQqd4ZUM3zVxUo5X0sIafAanTSabkiLBoew+4k6th9xIBTZ
ANEogiefk3QgK0kKc5PMoRL8X2NrQjXB3R0GV5K2gGkuxl1974LRBX4DIdP5+mEVNPJPiMaKsAUo
E8oZNwjw1NqxzRiANzNqmlR3FfWEGXL2s8H/6Eiij2YXO1iyCLZtVS/yWLTnEyiYyacAPNtjDaA7
YolLjWNYi7t7LgL+iwL5bsFXlPJIQMF4BvqXbYtHydbIeqk8JakxZyU2gTEp8DXLMIcIjUIJ//j4
y06tyROZBlaAw5BtJEfrMEd6zbOByAmd2olkLJiICV+nYcGlSUTkE9RHZbEPoQEY3XqMiNa3Q7Oy
cN5jPcVmJOyCY9bJi4c/P5vqdCyu0WyTla+XbESb4D4Vq54YMcz6JwhJtYZf/rQcl9LGK5rXXzhF
q8gMv0BA6K/D/0ZRXKdjyxIUb+xokitnAjY9eTq+lZhwfhWoO4egYGX/bb1gFcbWUE2DwUdGn2a+
bTVd/Mk83lt0q93inS1MdArd+hItjlWeW6MR2NrERB7rT/w3VY8TmHjmLPgHYf2CyiTEDH2y3Tj5
SVSthYhNyhFa5YnJKzKT6CXrhpDk+mtuF43dL3CkJy4q8duq2h0G5T66nV74pzJOOI1dNYEGcwER
8NBxJSiL6sSsMRnWroNpT7EcXwKJL6hAQTN+rdrpjRN23/XShtr9R++bHVRvjMcxgB8RvOmu8EGH
CfJ330OenNApBvH+Dsikn2LlplScebhpJusR6ALrL/EWzd4EC8vtrNvtZYNUucgu/k2sdJypIaGB
Oa9wuZU7YNAyXfYGPCwyTuSyIG9NLCJSXQM4ajnj7CPnsrsVzxDYp0bDdBopiaaIZxguSHE/PH64
QGUoyp1pGYhex0vg1lYbbqZ/2WiBbuTBSbpZXco1bdLXVPI4lJbf7A6IaTPOfe06I2i7esdbunX6
vViYEurdlAEqnl0Y23rsvy1DXlff6yjmX60xvex5fwAb1OhrsbXPPTw6mNf74oDmTJ3vVuie5mil
4CQtIDSDqbpMcvQ/Qo90I36MH6MFwopj6blusSmm/nZUvgzVRUSvFs2QUSj5e6iAi8zfsu+6eC4O
pAOmCVxc77RH1fuAT5MPaMGpLgRT6BVQhn/tigjphkyFn6mDHZR+xTfXrrxrVr3oGvdA1+b9uwxs
2Xum4+D+H0S0xGfOlou0lz9NRtYUdvccSc6BH6EH7KpW+z91K1FqEMw2NgiNj3heEsUcDJTFmYuM
KMy1oBq3KnOscJraw1RXyxjYUVsFAEYchBICCYF0WZilkTBMFS0guKiR0kUdMYZ2v2cZkKpfSMLV
qTcqw6vx3ZDPM3lAfn8ZNYFJeMtDozmgOVBkE5Wo/IqEsGMw8hxgUDUAOOOIm/MHdOx8V9Wwse5V
wFLp8AveaSqn9Pf1iYdZAR9OgPhTl7t7F0aCKA8E7o/vECaRUgzyGucVRSDq9QSXBYeteVlT+Dc/
sxvE3d2q8K1Di8EIqLQ43goCX681+dqkZWombURVcgXubzeyaijFZbgDV3qxXKX1PCHHY5WXJO3A
RrwbzaLfR6fKjBFygAKbElnZQRYvbl2usvpOU2fKSdDdPn53OvEtcCk+Z1AVYuLyv96Il2gVFab5
2wFOFE+mTb/t2WKPazJ6jFOExUv/6iA8t/00wLMRpnGq8/ii7AWGRkA45/LZ3axCIS35KyKGsYBi
PwfvzC2McLLO4ydMnz6V/zDqx5gCE1N1Uaq0m1zQCcYxZErlKR0hj/W4K2979hOrn48Klm6smo7v
jTwELlm1o0yVThUPkE5/nKl9lp5CDaYJs79o+6bm6Knf3Bsh/gvlDku71//hHsz6brZKNPEDOWdD
7qQ1s2pEEv1jYz1RKSlpgX+ZRw4WQBLLDsKITARSkRa1AAGze/yR8nDHKy1ZRaDEwfJJrPAkwjsU
/ESYQnpJhCDCFHAkaEMMGCvd01xGKoYvwsiPMnB5B7CAihpPbFEZ+izC5AhZGT23cSw1rr2/oh9n
jMl0gmnS4v/sB68CDWcveN5F7iS6U8mUGkQedVqNvoMvKd3wXAQTVTDgVlCfc8OrVtI5rb356D9Q
L96eKZPN4CJRC5jbc0Ec4V6RXIaL50RAy7OHgpM4LhZuJ7i7unRtutkgnAvckFLId5bGIbWSvAcR
iGTkRggcxUTe9cnw2YWxgxpmCY4AwyOztx9tJB8C+ODymFqeBbUo949/j9K9ykyhsRn4QbpWoi7T
6Oj95Ipk17l0Plxjo8TtO5IIKV1ZYc8LHFtPmYYMB4Nu5HYwD3Yd8xsjMrCghSN0EVqJ9zKHLKRG
g5gVopbhsT2p8b5MUpyas3PiZO4rbq2mSoQzG0blDuyihH5oqV0d/qIrNFCWRAoJIdGl3P5qY/K4
2ZGpsXwu6COXjptwnww2eYvGGFxK8AYlBmc6BSJ3MEUafN/ZHVfKpRvuAybEpVnmd+K4cwRkPWDh
6WxB0qPOj2BYCpETHaVzdngOY8OXkuENT9XawRb0l/PbJTDPh82pIY2/1RbZxVSI/cH1QInjQ9Xe
/DzLZEKOspFC67CFOdmxo/Q6/jf4xNPI+pVeKecWmC69Ew2g4IQHVm4T5MIK/cOPGyphbioQ96H1
MpCgiYOhct1EepPAKVeD3kQpCX0pVzqc40vUKegiPyaz0qM7Ks9GRYvVEt11MbsVPzguqrc8yyxh
iSfgIHjgB2Eyy1tiuGanCCRJcUHycoAP0z1lFppouNvoL34Fx3LiKJ+8z7RsuPhE+qMsisuICeG0
pvtJ3fCpCVGW7eAPUc2qO2ny3+kn5p7u0MeZmHMmwbNyEWgednroFg9/yQ6IKR7FFzRff1zUnFxD
pbQq0NOff4lmO8CfgO+RxTqrfSp4qpcPN6HGANpNTCW4gfk7Rq1GCkI9Tdn/Z5d/p7M8R8/ZTWUx
mHhMQ25tB+VEjZJ3VIXVjNuCIX7Rnkg9xCvw4+djSZEygFzkeS3oalAvKffbKRZYXlM9Gor6UUxE
GRwgJSfS1jD+b4LHLr9kuIQ4mjj228rLnwQ9RI4cyNU6GhJd3Rvutu+zOPisqnirokqd3rZwJEjF
ROALOVc0RuJkaa3pqE5RY2LQ/1ZZZyfA0FGBysUM/DxJY5110MEMNjsNlDZvvLLEKht5U9xvYwma
SKi3LwqGCJ+E/+aoFFSoaXaUM0uhP9zGyW7gU+oEeWRBsCtUn7ZuveE2yEbehyAuNAauonH23+em
C+8wmQ/2GJGeGWFlSANK3u54dimZNQW/jtjqT/6VtoLVMQVwpVj2lxUf4qNmazmty0/+rz838kCb
PBbNktZka4YVe7ZGhsXE32ajlnZWIkRSAFntdqIWC2lKGYZQNWCNiH1QOPad/ByeyvK2JcixhG38
PzQPs2lN/uNjpYmFYY9WRgoRm1+N2XF9thYGhGXiguvLb/cBwjIXmjsFdygh1O48V8lBODIqkIg6
lVnX0W4j7HxHi06k4oXHk1kvDi3kY6nODMRvUISODxqYeFCpQA/mfg8NYg6/8jhmZ5rUbcSycZSY
eF8QAtOeLCXvatRJWe1TVURaNJT7HKjM1Ru6gKXIbWV67gQbEDRRy70nAWJ2ViDtQfxkuKRBJlNE
spxxs5Mnk4grzlo1fOcRzzaM+jZ/Q+5Pxph5mIiYFU4EumNeGBuqs51Lfr9QlTHlzc0bUlfcliAu
Z8GZp3LBcbTtewVB6HY1E5Xs9Yh5WMr6Y1ecIkWh/COcFNZf5D3p3pL2bMKbb4jHr56mrFIYHKBy
K5Itzkzzuhc+MMJWhGryGtnwKK1aCZ1IXPFOj/q2EL/DQmT0McR0fxHhDHg15Kis6y6KmiD3UTJk
BzheLJxmiLEik/L3rtkJMCmWrhD1DxhITDzzsgKYD4rDmhVu2ttvw63RWcBkjZQ9wZjAVWEiecRL
dTFHs8fqT7n2f9jQACbx78hEHmlvyR5AhBRcM49xHxA+ADjgZMF0ZClozdTX0wCyZb3l4mqRUK3t
ac5XOcr30iIZrXKAI9SkhHUccJclT5pjNDtIWjpX1DQN1HISpoQmackNfd9V3eXEPH5AFv/r46uL
PYFsTB7tEeDvrar2zaaEw/zvcT38JRQmA2sVWnBXUicq9dIuUlCCqF84Y1MmG3VyYa1WHq8O9a5i
4ROFpHrU6Y524jJk2S8mXZUGa7BzLhTf17TGC7xngJt3TPsQsIQNe1C6waurkfylUxY2m9KY7eId
k6YQlqEU9w0hHGiqTSDcgknMm80jnC2CnI6VMjt+lozYm6Airn7+YdTIrV6sovO44NUrIEsLV0SL
mPuiRFBns7EnBxoLARHwhnUrN5BAaBUaofOLVobq6ExUmhE/zhclZothaVMdadpWljiK6jPRVAKq
xS4LMMLMAFn/0Tme8yCt/Lv0h2IlrJ+nLCRBMn8+h+dLhWZ8q5+9cpK5BKcWgqUrWrQBzGKTHm12
rnBX4lJrM4h6vy5yyDbEhnbC0kGxZCti+SGqqY2iaELNOLBaARtdbwqoMDix7gFv2F5zwLrCBBQc
djtDWzPlUZjz9PRctLilb261aRWN+Pvo+li1z7CgeA0XYNVdlRlP7Rwrf/iOHLxSTs6MD+Lpnv+K
G1aMwS4cJOmDffH13x9lnK+FJqqnQXGpL4xxSKQOXWoB6ySViwSvI7YmIPkJRaQoGa+jDRcWHfLd
SHOM2sYBQcyyJAPHawuCmoYpbG3MOFyU1MvZen8A3pTbHSlEtPbBXnBe7ICaIUkuZTeFx/ZbfytL
+t0Etq+LamGqF4EuIL4e1y9GhIVH7BbwynJJSnfjyLSK5W5w67uz8GiniMBlYJPjx8EDtW/19d3D
7MCbvMVxooToFrqrRBJT0JAmApnNRaOn81hWHzYb0uzluO2MLy3QYLCihnPgA/HbyaylVnd4ZVFF
XPhbqe77LAO2LPpbUMGw/10fNfq6aNFk9oGSWMLHShLWC/edPGoPVA1t/5nhha77xQM357HBcpB0
jY7zYCAK9z0EF/WlubR/pYA+ineGscJHaEUlepm2A+jvDiBm4GzvE+Aqgs+n3JPhFRyFC2zGtT04
0Lb9qL1zp9FwgCrkL6fhc6yWDD5+rUAbT5vPSNVeseeBPFejt8W5tkJEp3H8WAdIKUjP069jBWoc
sy+Gwx8c/ZQ2G1UMngLPtQWYkez6QRPoCHgwxRdqWPBROHQbVnyiqW8QbD7a/nEsQb1qmpvbvgPV
zqT+84w//OtVf0iMoYGyr8s3R01U6f2s3V7TeJq5LmEQeQV2zX8C3tXgPnRZMfVYcJsBjXsuC3yx
EPZllt4gwNzc2zA8JYtxDRkb4FzxEQaOz5Ks+SS0g1utyRx9peL4b57Yi9QRGjrgYI1VrKV5e+tI
4PKK0U7EWSPFH38+s29YRKAb3K2wp61pZSfDZGkBsd1JFzmZNJ8v0zvtwuKUDGCXMLaf0iIyi2mt
s4vUNvwoXBCn9BCc4ej2YnyEuuZJiRtEQ90T+KpXz3jq4hZ7PSne9JEXU9gMzUXt3u3eI47VV7PN
NeIf16GPF5ijCmyPev5UfFEh79akvIttqGXJTmYEkzx4esbtnDJGtGDHXh6FTBx9dQtfvdcKtn3l
jY/FZe2Up11sz7WZUhraHSz+KvjPivm/qKWCpK8Mi5if3/kdr0J3LL96qkXjylWErcY3Y2Lgl1sj
O7b9KiBPJ3Dg0xk47KeaE+dNF9aPHqzv1F6Qs1YTfrkO1djJM6/u81c/a8z9NRezK51yYLqMWqiQ
xy6V39nd5PXJfykFBokKPoiKVH736d+aw3ekfBFjPEvwfXOEleVaNzgZUOAcyoD/W4LRX3ZbltI+
0fEo07DahQwYDR9NSyKgI/0TFSG2rKZFR92NOf2AgO/CbXR4wdyAUuguObSNaPTdl8x/3TPXIqy9
e4AwB30mtDUbR27uuFjVpgBLvB5F+val6xMn8K9YWEIgYtdQlKOYIurZxKd6tm7ygcR8cBSijMTn
DvaMGzBvqKufFTM9IAByi59i/7+Tt26SzFXvCpcOcWLwwsx8yhp+W1yjDzpSYDHkROfZCsqMWnwF
b7VOQ1GsmHEUcsyVofL6XuSi9E3gopjwjLGkzOgF6shnvPKrq7SwJzLaxE0WjQkkoAmE8Ic5CndN
PtftfYt+3pmfielTDLQwuE3YCKI6CUHBH2OnOsgJt4RPI2RF0PlSm3S8OLNH+6/oybJvGVchLsES
dOD9bYFzsgyTk0Ddpdbobhe0bfF3ENsV91m8y0cb1vMk/F75CUyQgowntT0mqC6nKyLgBT8pZymg
XJ6fB0zyHbwVnfe6HPsQkk6OO+gz/MGqiuHsAwCIfnAMQuUTLwIuzShg7ov2O77wz6DlETkeZ65n
TwJdiHSAw3RYiVpqDKhsPQ/6P+BucMnfrC1Ce2fyT8oX5e/Kgjb8ZiLbwtS363b2y8EBX32W8L+R
whlnQFO5QW/F8UhCjrmSFfWOckecxAa0ENQ7qGiZh4ZXSX8TUcuoqI3c5klKzTuYaUJfmSkjJreD
vOFYWal6nbGbgGnkkYpPfi0Z26P6t4xHvdy31O11kLiLJHiwkBHKftYy1qtlKHAn47AP4G+NMH4L
My0+FFrBOvNAar/9706xSwytGRn4XWizHoEMt4t1ma2eGuKOU+B3ZZIyg8vRKZvUM84ioqiNScpM
JlpvPMEJ6RPJx/7bVm4ooPgBXi8/FrvYGJQ4KrFqQNAQ+D93lH2VObK4RGh6JU2Uvk+078hf2PC9
mMT7uzR3uGRNRf+gWcn1DKOultlZsmZMs643ajaNy5RYebLRSsDAGCFUKsJHVVoLmG0Aw0+H6Ec+
DUuoF3rCqdQcfZVeDixd0lN22Bj6Nr1/oi/Eytni/hC1FuVOsKabfI8B9NOWc+nOhAH3hCQ4gZ07
yAYKJ1xijbSTRt1YTqti/VL+C6JbFMW1x4eLKKqBnXQx+Mf687sn4m7fnhXujBvqWfYrgFs7nUuW
pkUSlTis122i9Lc9z0mjvWOskPoLPCcnZD0+PZOEmbzWus1h78jEObMlvzmIkk/7SxatGIwsPJx+
jdYiHGPEtPc9/xonQdLw43djV86Jl4G9p2DLu6TlFJzVIivAZicUej6FJmhfh1eOgqBbBl4pPhTz
ns1qQ7XVKQ1Lhj2Sg3Nyj9Bopqe3GwcBOe37CkFQpS0yHQ22pvV8d00UYh7LN3ouMRanBIu1SNcO
sg0b0j9qHRElqZ1Cfi9FZPY0KzmJU4ccfyHTQn2ZUCqgz/wKoM7EczdTtpVdfngCe5qbRqRS15fm
FDbBtSJ+Kh6s/61QRbh0HnNbPtTHwt/XysXqqWmXxFt6+klcpe9ImXoyRnHiLeIcMtBuV16lcUDZ
1GMCd8iHGQj6a9Apz3qb/1yt5xkZTietWscJtN1GOv7S/CMDK2CfPA2jJhW9CZcEv8K4ddgmP1FO
/li9C6sv0oNxgQolnA9Scg2PgVU//R0op6RQAMyXT+k+TjuRla/SlnM+2ZtQAzosVsDwOebY+A6O
BELezMF+ee+5f7Hr1pMTC1oFUOnQCj4g8/y2+4Mbl0OOlAuma5itfMRX3YXaikDP7JzKn7AXlQsj
oUsvYUVyTJayO4NM6hD4y7nMB93TzFniXuvDXcVkRGihIdxaTqrRFVVb88JW5p3z7krFHNRPMQyV
TN5aHXgO+xD/Zg9oqpVhbeoQhUveyAp4F0GeGe4Pod6Y7CYlze0yLg3WBRkVmz0Zp8EXVDjRHQyo
eZ0x1/OzqHI92n6NbEDEinwvBtbJ9dKQC56XaoANkUeO+GyReyd48ppIFMuCyYCgi7IR+on6/9Ki
R492YMr5yt6JXMstLlouhhw/f4RuKIlHtt2GxXV08sLU76LfV2zt13ANN6VtKRO+mjfsXCJNnXtd
kBce+d1NIiFRtT9kYR1IS238QRtJBmjk/hI2c1rHKu5hKg2bGLNL7C8gkjvVtrcxMnHpDSjES+GZ
/j710zTFDEOYpAu1/crZZ6B29VJLbYyy5G213HOKtDHBW8r0VzznH/TTznMcLW/KvPDEXqloEwjg
qhBF5eYmqVfdShsiRkurt7sGCmICyuXxEZdEWOGx8dyzNNqv2CM6VMQ+vn9U4oufjex3cNmGjOhc
BHnM80x/lUejQstVT8fYEPEk5QpmJD9JyX4XfdFDz56WozTkZV8nmtsjGix486Yl351NVC+Qaez6
3JCKe1YzRP+pkdYzYsCmtr7VqiLVbCTpRNmTvHYHU5TnZ849lWKrxfRp4rcgWJIeG/7E7Qe5fGNF
RMBjH9S8mpqRWiM4VPwYURr2Ypq07/oZ7a8KqiT4ltb7UupCVJXUitkXzIHRRPeUfmB1nKifgD2v
gABsHMZEPzPqkMbT2JHbRSIDICrDGw0/dWEuWh0cA84KIkjSSbCS4Slo88CXcpXt7hMR2QwHK9L0
1qInKz/4A3HO7nVcU9xlG4U1XVMvf+/mTxwOvH92oyTpBgIsf8wKQHRUDhoRo728IR+I+dBZVdto
4hMH4f7QfK5kJtK6ysoncC9XR0F89LjyiiuviUZPI32+GqkXK41xbk0/u/I+s7+5mm28qh6SKiXN
RmyTfgZt+rWmCMonMQzjMPDcRH2Y1P08Vkcj5XS+TekqM05BgvQfKc8lTLB9LlVzraC1CStgKlfw
5JVd+hEqJBuZrYvdL9UIdtPUuYZpI6whWD6GNmVnNJppxv1KURRpjjVS6asq/KD+dAmFIh4CDlPV
hZo3gIFz41cCDm9P5utCgvkN9PbTu3S30AFyUTwNMoOa0t6Oh1GfIWvXQ5x2yFF7OlZ3j5G9ZMRD
BomBSANNMEav2BKyXBICEkBFGaOChixCYZ1rzidJ3XZG/5DRoho3iMhvRaT1wZDAsSx1RR+WOFfh
yoRYsasPlLMx1bzMYebJK9r3rIXJ3ogMsDG3fuX/hH8xE3k66eqGVTNCBASNrje7SIRGM/QDFlpE
78vUkQLI9B1EkSI+xIO50OM44792OiJm77WRup5PxHAkzUnm4U6Pw3ITmki2KLQbCTi30/9BCHUN
Q6MTVPVlYVGYSWB7sry+l1PYglIRDS7wZ9XctMBickoAU8du8qrgddoLNkSVwOsoW45G74Ex6wjU
Df8CmAI1WRXxAuD56scUXlNY7PJ2lKRLQvsPz/lUj6845TSic8+E57k7ArYQ1JZY7nitnF0u6KQm
0SttYiwH62aKgfSzQXwsCo24P/BkBvUG0tqEwY8zQWW3Y7cBnwrM3+KwUovC33Fbi1BOwphNUuKn
VU/FKKvGaC2tHGiOhTbYkH1/gssuFDkNwQd+XltPyEWu38V5GIk1M0f2OzDO48VafRQ+RCDyHs9R
A7nG9TQhLASKy76xC4TZPSXYAt/RzF2oAobuUOMEct8Uggt7bqMyDB61yYs7pNY13K38kv6eFOQd
83F6OwzAfCUiIckWlyHae9KVvoZNHHlZFgRzdHmAHwg8se8nMolb2L1HyVcedFH30EEdqOxCk+5Y
jWq9n5SjL4It35UritYCXq1ECGAy3rtHoV5gstvoiDYF9D2l/QvKjndHjvfp/LmMS6dsoP+ae0IX
GVp4UrAMhKTo4rGf9DBftDw6KFQVyy09NiFxXSiklfdr5e3zJjgDBlPF4eglXpdtnQ6Qq1JkUScH
JFijyzWq8ehTo3+GP9QaRunVE4OtYkC1fWH9dH0S2QvjORIHbkCoDqIufYpTPfvxg9iMD3gmv522
j+L0LFkBQvx9lSJCI/GPvYHpEN356FhBwgUUs/24/hQ8FICFHBGl0xdxLIZ37H43GLcfmzJ56pRU
NfE/QwQIQHygJrcaMWtyspYm61ZvnaCmjTp7Nl/D+0RSJLllEgmlPN/fb8yq6uH23HdvycC/8fuZ
dNGB3u0DGxOzcjaObCGxy4kmXBaJeROxEquJw/69VcQzeH++MgTSeqHCjn2CO5XarBpYiavJWcaH
qH8RlZDBd1n6bVUU0c/uc6F12aWGyUjIeQpfyx/lilgywBiild4yW4dTxQfjI4eD0Y/koPv+J5ld
Ok8aNq2G7UDfMVxkKqum8f/ZLTNjTTNi1ru+oQplxE8PZQUURN5yeWzdGHNFSl55KjfD2UJZY6zP
VF9+5MPPmjsPX9fj1jhTTrOvkt9APW5865qwJSdDdQdOIiHCMoik9IzjxJj3tm8Mx2pFI/E+2snf
RndwOYbwT89F61gojz3F+TOZ1u3ksOoZ0UT91Ev3VpDfgVm6ljT3Q2Gjng8BNMJ5HKungq0NyXuB
7SZGIjPR5R0ul73nbqc4sfbMKV4xtDVdx57KVE/DQzoCoNvk5sBodQyREU3j7Cu8yDaj3yxBc/0E
TZUZ1ft+A5YlX19b5NqodrC+deCaehU6AdyCRYYdJqCt+6uyOPJHBbW+E4eusI7jgimRawIG+qDb
gg9c7JMAmhTwczpZ1Bz24pS5WmjBhT+wr0OByvIxlWOK7uAKTVT3AiZWqb/qvmTPUTI9Q504b/7P
kIEkNuLImQqYWdDfTq8DJYadq/EaCx5IcNTbswNyc/V81Rngd0wIgqZTXIkfwsacej1MMAHdYVZ6
Hf2/MrRj4IRRf1/EXZ/XdAopO4ZZ7QxLv9hJbto6nS9H50ZYMwo6IztPfVX2Hli5HuTw3JF6oOQ6
YNJGykdKKLIizPeyneUtAU/U3qrsMFv1ZFsYsNOv+Vp1PzIgCNpM8yDPqLyduayaDlFgiaZdHjzx
GsynkbG1BzLpxW4dfgTBNt8Km9gCiEAFnTZyj2J5/YfGGppQw7i/YcaMaMbTJsoj/Z/zIpZPIJ67
F//r4aIbF7F7CLBsRGOiCOLcVtJ5OldoSPhvCNzlHYe8RahsdiuvN+mPJUfkg8YWiqgu5ypM6eK2
LQirYDHUcXgFzEnBZqCnQP056js2C+J5ZrvljAWfv8qo8rqiVJmrDtKtKv5ti2Gks6PJJhQ+qmfk
ymh3pei9wircnV/tQAUa9coKXYuz7X6rbtRkSGxcqWmtaBdkSs97Td+cJe9SP3z5I1ou2neRK+8p
daYybH78ulgK0K3HQhn2znUYjSmGM/olXNht1VfGFrEEAKSEBHmPvl1j5HDBKWYMRBwpHz5dAW3F
G78A22gvR/eN8XB+TShu3YCaxrh5Rtd46red+mHmfPEDpmjYVi8JY6cNrBdfwdLoNiTOrMUlW/pI
HoiZbDsMUC99C+uv90Zs/9sGuugexiOkzrq0BIh0pLwAihMHnvUwRsQxxjHwxYoIeeicCZ3zDs+f
PGY1HxShip7Aw0s/oxjgxJr+J7wcL03r2dlPYhk2Yr1Jw0WkLkOv8GRqeQeLy99r9xaiux+wOriH
vxtR500i+adgskzIj1JN8NLd9QYgAseC8qHjcPHi6FYmGynXtMtvozWrCGSCzpGGaYdROcaJCWi8
TmRarqpzR4yqvI2DXSf1lZkPawtgWN5KWavGWIRxoVn40uZ2t6G6QOYnejkw30xXaz+Xn7ReZdeD
VWpe5Qjo8Q7vzkGHwAoqMXCpTav5oytI0Lqp5yxwlyQ++J40Twrj0wsn904f+77nymuYgtYdzfJL
4QbGiTTwF0afxZEBD6mOBL5R+k0PTUByM7mody5J1UD2bfXnszB4Y6uAUQ30KF6KpMiMi2iUQ9aN
dMYMZT0Oaz5FoQk4pU9CgTg3oU26h9l2qpLIewD7HHL0/fIYaAnwRhJz6/CVanyLEWidOWyvKjAd
t+ITKl1MCHDsM5LtqjptQjyLVvplk07ZoiGQ9M4THFhxG1yi9eBNirKqwmliIWqwLm+5bW63P7rW
DvCtvwJDot2TY+YVxEneZsUTcmKUrIj4fJUpMz3LrYTETnZn/lrCVgFDNO+Q/1x3qTLs+snGDakJ
2bfG61JKvo/PnD+ob6YFotsgoDJWkVp0svPQJQ7At6HcFlDCeKIkJrE3c5ffAOZqjLlVZoSY1tEM
OzxoTN1E6oFx8mh+NZMiZFxb9WGlf2WPH8yP6NCxOTpPNyJI+niyOJOlq0N3N3VIO5F59GDs26be
effYh46+um0PR31pMFTaqhWmJr/f5bYM4fwhrGJywX3mz6fQEHY4SSF+LwqcGOSG9YrY6O6of3y8
Fe5GIdSI/Ey2ciVnpdRCj3rDa0MMdSSMEh5RenIDP8xBRw2AOev3Xz06MTYkNYeoBDBEt7M9FRQ4
bzvfcU949yxZNaa/yLY/I6EM1UWrPQ97c2XGBDhV9ys0z+IRwa0daH3pjosKfOifdZJeRuggjgiz
DrVFKcdskY4rB0ZhO1ww+pGGn6XHhtrZ0ubh2CQWNkvvxtVFpRdR5StRORVqSYdUhiYc86rehy2D
HNurQA7UKa5ETwYJstGXqadcFKVl84NuZBHeUv1CnEMejkrzZclrge5BmNTKeUz/R5+42+k4yFuU
6aphj0rWInIdvq72/VNzHGqHjsDSjA3bt2kQn/xnCitiBWkx8I5fvoW/6ovXsn/vsMM5PU6tz9RU
xHgumtsKaRO5KWaeeCpYwGyz5d1vxw4E7WcMkbropCh8VRB9G8knH5UfXYIEgiBSC0Jg6tlq1OMx
AYft0Xux4iuLgnCdMnyfB2DjSuz/xnUdTBYdS/O8C423S8+fJ5U/GCoti1npdkjlPl0KsGuE1306
a+WKJ/yDCr7sgZWJwBDjcVNljKUP+tNTVqViBfCtEyawfzzbJMzzPo/7GmuPP2hBZ0ehIK4d1+mf
1XFSQc5yfl9yuo1efLmz3R+cQ4wefkvUwOcE05Dn9k0JwJAAV2ZTX1dq+Xc6SFhc2LYrogMkhFtJ
kVT2gYAIcEelglFJD5AvcmrIil45wli8/EW6mKKbRMFL5q9rxD4fh6gfilG8Pm5MTyC7f6EpGZS2
5n6dsUekP9TMP0GfdD44/ZMw52EQzFVoz7LLsmxViBSEQ6GGMBOsSBMMn08L0ZuD8Ph8RLT2xpXx
9czhM5wi91g1gUe3c5zZeehcf8rQI9FaKCGGCYjwx4qk962L01lj0bVi1Y6YW0V4/+oDWRc72sp5
LHm+DSRoSeG624nqalGZMixOx0xHHdNQo9/Lyj4PMsvwrGUPGFCcaUvvFjht1jlY9B5ghbji58n4
c2ljTRAzqPV17LsvP8DTanhLlkesHHPHOAiAD/RkiObYll8y6p+NNXWi/prT6WvfK7F7I223ZxeO
va36bapxxPCGc046h72sw1pVw76UNpWUnATE4Oy6wv5EhBff3RJ05nr4schp2z4s/7w9lWTZ+tLr
tdhE7UJtdJgA68ZZpjmSsK3/m7xZsZrrYKtGg4TXLKGBW3ax7ti8f+Yzn0HkQl/XWGod0pHHd4YL
OHBEf0UPVGEFH7ShVcjC+54t5UubUC2eTeVh7sAiiNpdV99BQ0TOZPWa5jVRf+Vj7gEwL+stq+2f
IUkclvcOEwok7SgBBDNGB7UgnU7OpP77lTE+97rTzkMxhL3n3K/XbSf8At7hVmv05egjroc/BwS6
YWRWQ1v/TE8/0C1WykvmzH+vWorvItxwytgdfIlnXA0qx8oalnFK+EY9FYPddMjqJbh2H3L5fHge
FlNs2Fb+I/kWKZ3nKqsMGKRUT7kIFPhpC2BneFyetygQV+cvd8GWKHH231b7CMwRpChme5APls/s
EdjIooEUUiwtyNj1onTQkaOELj8oFOPRheUXWBnEJw9EbLiqVCcGChScPOlDH1FNyYDZK7ieIsQ2
bpGqBJ5s+JgXBdawwo96g1fikrluZFKKg3MKQYsWP9bSn6GGSnm35NJYrFnUmvew5ZbAG0ObKV8p
6wdzuuLfP5hKkp5gzpY0/jr5NeooktcjZyJf1aFusR9PwkU+Mxa7J86f41l/A+6qkOyHVIrOzptU
tinaKFwfKu+RHGLFTOLsYdJc/bDV/aEfiKe2kc4/CdNAPMYIMPMRn/0HBa8qkLdleSi7eocvm8XP
jEUsBVw1ao7YC85qsW/Et7pyby2/EPNF6KusMXOTfClOJDwmkgMISaolCfIh7nsIFxJ9DfbnqcrE
1w2PTWn7t11IqrzVO/mzWjSFON51iJdgQ6KigkPwDXkZzXKrnLfEQQxg4xFsLM7HMVT7wmjzxc68
RKhuIg66RvdI4gu+A+cBGHzxZp2wTA4ZW5NEBz8QBwmp6t9ExEPPT4nreSvpVSI13W7zMNHek5PL
TurbDpMPAo9sxcFV4Uf+LZghW6emTVRFJ5H1/X3d03JBjqW6blPPBZX66U0OEBEaJCt7JnC+ceZZ
0cIlaSRr62XNc2WsB01CqDVi9YY+nyxbZ/ucjXDKtYur91JxNt4P9AY6G/m4BBvK5hW+5QWdlTC8
RRMIiesdPKzzRAn9vmRvFCKrKCteN27LCZqKRqRJVoVu6/rqOShd9gMRa+DTyTFrbUo4f0Gje1ka
vFfhlizoBNMGtyZNp5Gij3F8GDrsjuQ+GlI2BKWCcpJINBuqjVz/aXa635TeEpQCHWHd0i1ZY3Kh
Neh4rMObCSZgSnFwsVYGhM9XBd7+F6RgB6VxDaJiH/2k3ZyQ//9MUX6byvHhI47vMzEUsIF1fdtv
MoBkC6OKzODhh3skbrOlCiSwQ3U28kG4CNViqm3qLuXiv/KMZja6+kZWXu5JnTXEfcS5a16t2Orw
+QLsj3nUcgxJ3riRFLe7fFIQkcIWDsO0l6oPgvxEI6Odk9LBElOuHxmD88bjsTMqXDLwvmVR6hMK
AvsE+1iA+ChZ+niJD12xWaBUTFT+uqSmsaP/dirlps+6zh67SS1YH1+dUpuXmebiSYbnswK3J5Bb
ElRBB6rD+CF0vo/z/iHAs2iuIQKHdSu47vp+1Bw8zFGFJvT5xTPpl9COSLITG9/amj53UWS8wCtS
ITEvyYM4KoVpLdpDGP3ymG6Kn/TJ3nEWtZuNlHEq776ZNKZ6AhS8zmit5aVID5BSEx59vBGamoxX
R8L9bs/sKuwptV51SSGjvgDO4VZBxFFMav1Vcur7RMmn6oPEint0UlczdCgmLLBfb7Y3hJHpdWoT
somCs4ZZi4gVl1q3Zl+gGX0DDRqYFQ5NIlLgBfa+Rh1Vl2TndK5tB4cTjVY5Y4gngzQBTzhD+enn
DjuoUhHTd/vv1fw6WRk3niEBGVGIBPHn0CokYtS6O5s+5J95d/fK8yTt2M6qBG2caknh3SZneneF
VRM2ZJAFSdE5VX+Lz+JIB3AJsrUEmAMKHWuahhBeIo0lP5GW9f2/7xOcs9y8eO9B9CQa+pq5K0m/
CyhJwjEEv2onEncgn0pVCUzLFEecqlXCXR0xNsJ+u3+p5LypXXQaWNrvb2UbsNXIzJBZka/BkBxO
O6Eo20/4TP6wu4sCdy2p0ybY2KJV9RM/EZ9wk37G8rjcqmY4Ce/PDPpnoM04sddyGeCU8qBHF1ol
UozK1lKjx4YQaeTk11xTKtsSRmhAE0Na/nmLTRkuODe7kj76I3JqtmFK8Ps1BMUkwcXPKo/jbKU1
g0xcHGoIj9NDYXp64fFH2Vs6YS6jxIngJKctQ6MvYNP8/mpRnbKfRHQQTK+LGy7en7jBLr0WJywP
ktYPxcbFhQTNaiHoBlX9jNCWgziYDvx2Kwehr0a6sOI9Zrk97Tvue+T5VDJmqilOc/wJBRKnZ+NH
VXOAMGVfvRFKYNay8oyKKK5sqnnw2aDpJJsvT9kCH+yr1XRGfF1y3xpIWm5RBZQRWLds0XXOJ11T
36amo7lXnUYaCCas3sguS0Szthbn7I4RJbXqK24t8JIiS67j9muIGZRhqsBlI8Cjw/hL8RScbqsI
wE5MrsKUBQ8LgFVNRYmrXddfxosztUGy8uq2oPQOqAcR4fBK20/N8OrMKLR1OC0Xj0oe++6NU/Cy
hydb8MJAgfiYDExNXLAC+lH1EIsf4nJxbFhkzu4knamHcXTfIkkV9wIWFewRYUxSGAzb0a1LYcAL
djqvM1J3W9egmmlB+kUPUGS6ZUBGvSBPLA7N9M8spXFxmzBvzYpOQvCAH7MiuHCR2EY2fwLKGCvb
VCY+PKIfGuSSyjX0Cywq3I+ht44RoIveRdTRVXobFkIOj1qVEyAJhc6vxlksLCIdWsFgKw5hSM4v
V3yS5IeVjBWokIl6X309KTpgELvLRJx7L3pXuP5q6dbJtAEr42Jr/eFPOB2M6vtUxS4xTJBLF1rj
ofvegLhLa81SzoWlmwAXUsLHd8MJt4ZZO7ehFVRKGGShFC13Rrojl4CAEb1LzUayEebDnwJG+kvG
Ghs/vyzpQ00nvvxWYAZd5idebLYMRhFF33OynR4zR62Mp6CGm8YGU58Ho3fXYl0pc2J0OfrwwHai
dM+aH06rQ/7mcqXZ5TUlfORdHaVfnZ1L1i61WLwc8hjIcyf9QSj+rAGhbbPOx17k2FP4XqO1uuVd
fD70MSF4782F9+TvEEs7sNp4heVIL8aXmmVxO5qRuyisjGZaZkVyBOjZuMDFv2JNTJPgDQc9NVYq
SNBtifCWxjtDwS8JCXk85njvUHwr19BXpPMGLuUpnBQ9s4ygLC1yL8AdED4uPtP4s3QICtDWiPjJ
4EmsJDwQyzWeQ12OeXEP8+CAGTmy/TIcv0/mk+dUHzsv8ruPiB+tkSwpLi9rGWTPFb9t/zcC51B8
5Y7vaMN4mRVYMz1syg1kKYR884JD1Bu2GKd786v5xM+YewAU5J4rJaacI9a4KI8nmD+DQtD8C08h
IjKq5whmngrDhYptSK+3T3XaIwVmC3eXKYemGTvePdpchypg1cY2iq8ekSOe5nWwSbauI/iV9ByM
Znwb6fd/hakJxfwHPVpVmtZ7Rnx7h/5mY3iTfFjhPAAkLr6mMPEyN+YYJTfq9SQmvNOGoFNn6tPk
r/kzMriM3+T/O5kYbrGAsBrvOYWYI9NvB7eZrmFN2g5yDkMA1nHHfQSh/SAVCTGN4DuKMuANTaGp
9IoI2Q91/K4yRidPzWTVolmYmGOancuKzjVPZxIxar95rk2aVdrQYKZM5NykzNkqTdmxDLQivLuT
UhoBjg+1KkRIzoe70b6rAmZ+U51bXo7njqzbJ35ediRL0tQRLiOdQ/wtPKz+a/igdizG4x3WAleQ
Vwc+92q1gLLrgA6PJ0RRwt69RFpiOVJ8cW/2LVXbu/+t+0/FIk/5GWdZR9YYkHc3Q21+ByAxOh+v
vkcz9/Ih+fNgSu8GaYaiBYAkJjMKetkWiBW2n9qMve52H1zAa4GI+oCcP1E09QQ+x9mGiWdD1Vdp
bHD3AksJZdZhtCY8DwCCuJkoWU13X6NLItQbaE6Z+euJwVT05LrFeEgy5DaQN2ZmD5SfoAwlMXe/
o/MIQWNGM7TEimgMRxP4oTK1yVdxE2aPx9U8AUaAM6c8VjQeBpE8wnbdTuBigqci8tFEOoMvZr/g
bPa4VBnn0C5wM3qUMrLy9GVdfvbKwtQDB+dOm2AftiCEujTNHz/TQNMjYWxQ1Ux/O714SC+IZalM
BIGqtu43jfTEiHufy5GrT2ki1lRp6rcHiP/4sRMI+fmq+7gxl34Oaj8ZLOdBfVy7AbvqK688Kyc3
hsOX9CqV8Hr4OPqRkIyFy3MpydAbBOxieuPqyNcTEuuB3rUjBa+pQXoV0iNO+LHxXAU0UT0OmDL9
gYlFN4iilEvodlzWEmajq6/9vwWhgZ9srFGzdT2CzcfcqWdqCEi0Njw5BN0ZFFAExuJ5Wk/7hrhb
Ta4kzNdWepbnsZtxkTHAVgYxFIn0HaHtPddPOdhkXU0u7PzI4TCzeVXJlUkNChpWyBfm23RCbXnC
N/kLYJLPlLJHA5VMEiZmULckqn1iSD6f8EQNGKXprTC5kkEZ7wg6HFiOuMQVnNxiFwOKbHbNC2o7
nLycic6rcujWEO+GKihvQO0OTBY22DNbv1MQmmuB8efe/usiWRElt7A2CAW3KIia/ac8NxIEQqRu
mdISPxRw3l1OubrRIrL5sxbcNTZsDU2s5JR1+2VOLKnpx9qIq8UHaRr4ojRVJ+Hhk+YtJwy4ctgF
HUOEMprwBn+O0xFHpBCCikeX3hTW8VIaH4/D1puaFB/f1VCeUlul6kxxQQZiSW57z18JX+RV44IS
oO5cyYDxm2DEwA1dQt2iX09txAQeEz6MCC5goHOpcUZUGe66Ffm8G+XRJzNV4tV4fz/oUaZaiP4i
vObQjpow7Ype6CjQfEc9u+OyoS+XdhPiwkSfnSVvLzpL6h0AAvFTmWFEIZ0bIxbhQZOmhPw5KNuo
WLQo/o7teDrBfoJwTgXvcD6XNNbZDJm3shGzmqmaMpvdtNE1a15Q/Ymqm2IbhlojHt4acrx4LqX+
IULWjQW6LSHZshKXHKO7W+mvJxwb8hy23beikgWTgfRGslfcLhDFQi+MU+2rVltf4MzO1Uea72lx
nIq6a16Py/DI/aL1HW+eZkO3nWCBmfCZQZUqRZqelkktKnk+6CVY2eD0GC2PvELk1JtT5kBjavRw
oxVaK5NXYPIoY91bsoBmw3+ld+RfZG/mVESl4LYV3z4/EJAi/+l2VDjSBKbZk+9N7yH0ojN4G5D+
iyiqe3ptFmz/R64syRVx59qNZhOR2NmC4oEj910fhiAyU6f4eobvo0H8+hHszPfV04ZpdvTYfXb7
i4Ay6v2hoA1Z+2yVfXe807fvtAuSbCuVGaGWVJlgJsWpJzaILB2/P4KIr9ej+s5ZCv8FgMijkg4X
hUV+kGtOFWKQoDY3x7cDT3qRBGpn+QPIyWARXl71TXWXNmzUDWjAPwqJzZigKtE3PQlOcJaONfEC
Vs93ibQoVTjNPWplrt9PDirzwBZn1vLDFr1W2n4dEXBoSmnGtQQDLBKhRMbmvGS4R/umhK1RPkqg
IiJM7cUS6Tf6oKX8mLgDwpmr3Y8XC5RsSvkWUp/P7j7VrHs7IJ58MbPH29+73tAEpfNE/RdU+WPc
OiVtyk/5uBmqYM0thFVUXu0cCDyiJNfSaiipNDYg4l+MMj9JA1hFBskMWc2v4TPIn7LGBiSAVpSW
LTiflTrPqkKKpeEg8lzo2I6Rd+LlRMC8iZD3sAATdb25pgElfuNux7x156bBEiHjsfVAcfqVEEAe
IozSuYidXV6aiuvbExjWzqT/wIJn0wUQzHtNoDIG8BsQu5xcS1STy8mIS6d0JUoCCZxI30DfqsJG
TdNZKxKI6TvKsJE94yS7VEPRw8GHuv6YdfmoToJavaOSOvJsepLrUYJ43XFbwt6dURKPcOIqXRv7
gL237GaIf/lcrd+yW179ABrDvskTLIjtnHBzvZt8RgDJTxYNxDcAMgqWi1XyB8O3LNqLafYFLH9m
qGFc+72F2bIQjUaLMrXlWtcWGyUMESvW/V3rilrqqmYFzZyZe03aGa/WgmtArzHI3+fpqjZWNd9c
1SF49OGOuK9XX1DHaoBAeAGLRZuNqRe5H2f3mEmIxk6MUaZeXtzyTyU6lI0YUg1ehVBU2oNlrqkN
KU9BO7KEyMWAYYvyx10pBaMoaI5LUTovbK0epVWk78SNesR67m9ftdroPZyIsZRrzyAGKLEcfZbs
ft0q14X+x2ErDJ/ZyuxnHK70KwGmz+evvNOfbkoQxgkUuWVUrPM+yeOBHD92SqVyFnFG3r20T3t1
AMpSxw5/2r1tGVvHBqn5aJi9BGjlmUsaTYlKDdAW6GVPzt+/+sJ2YS7B9+A1PQjJsocVUHXqj52i
RxDFzkCLDlQz6TNnr9wJCblSvxV5EwCE4AnygVm3Hx1XMup4qn2VBB+dVaoRe52RpKxfXAYB/ldy
nycT5oKcAU5lW1SZ5Vr/RTY+MI+MSMQnRmT3mxC0SZQrNe/Xoonea2rcnLCdpItm/bzMFMArktz5
F+l1m/O8oegjNF0PHhFXFfT2aHZd0lWD+U0x3eqcscZrHwgpsRlmCNDYOzjVtK8nIt76hM0jI8ne
mSQrpqwexGPbN0TQB0mA1n/Z/XBM/ZWzqubW6rA3UlZ8zEEzM8VfMW0asRr4Vq87Ixv4sxphFccf
+iX52pHWftgrgjyigUu9f5uAlf186VhvrNCLgKN54nMBR/vpzw+XIAH7Icz4FDVL9QIqXdzyr6Bs
x+UaeC8Y0tpY2249PzPk/iIvkjq4DiRhsYgiSZ4FOl3EoldRgdUnaipIhyvDa0Vf/cNzzReucNhS
9zzlgR20Vd1agDKl0UUsrrdXjDzsiRfYrsPDiYworIbbf3rqRmyGpS08HNKjETUWE9c3RRQe2LJW
KYbmlXrTMm3CRvL77r3sF7ICA3dDI3O44Kcb410MGr+bSVrLBFnq0MtzE9wj6FRUBr3Z8FLMoiu2
VJXyf98omsBSwQDdbDkrEpn/tAIP6vIAppXDrX2byHgCBnwWrU8v03NAMf/UJNNGKFDfoyPxVqLW
T33+lJUfWmAm5+BbjRZXtExxAwV3qM51gBBAisGSsOr+f6+tTKZde8B2Ya1pfMSy0RrtBuryWlu0
5iYZIam7eCy12gNmEqa9s/yUIU2MD78fTHCL4cNqAY5BLwvslMe11J5SPVKAyss3XbXF3rHtxKxU
o2lGNu9CixqYoosrWibjGnlgcPIucKuoMIpz4Y3/mLKkguOyHRbs9sP0LcZzhO9SR216EQP6lxYc
ai223gupw/VVTE7exyOYKGRS9FXR6buZuzmVGvsJaEc4p1+n8635HMHUttP6KiPyuor43F6Bdl4L
20GUgaDqOI5I2cgXe8sMv7lTz45eK+V9JJrkuDutWHaPKRCW0GTy3u/4XWUPsv7uNa96/71A8p9x
ejKWaA5MqTlB8qVKD0ypSlewRkLxL/ZpE9sxXv8xylq4Dh0ex6PDgJM1ZM+VMGgB5J49EcU1jt0k
jJUc1uKmoUoN0fvqkAHyJHIv4z5afGsagb/faTnNyHwIs3F8mrcFaHwSywYf4bFCYvqohtfQINg4
APyeTti+5SRpYlzOnALA9KKg4thYeHQH1auJhzZ8SvMI167chtqzIkYPUVgceU3e5/RWeBWheml8
I9QKdvafqdu4sP8SUoVHBYNXDWJ7BElrRIn2F3/RIueshG/duV+GZ6lWwvAUk8Wr/lqZAUtyw4wu
HJT219TBkodvvyDeCpyeFXmFnAdGyxwRoIshl+1REGiSOXw6pRxgjBb6buOARImFwoMdRtSQfNwH
shfTbIuoCk1F2S/d14lsTlXl4OZn0KLIeXjLJNUkKd2v3KAP6gO1d/pjiyQF5BQxL85g57wp6FQF
Lmfw7KBY+P3iSe2SXOhQsky6LN6FkbbIxRNTG32WFZOJZ1lEqsRAUCIfqmC0nxTRqZihX8YISLlE
pHEpqaZC9KZZiKIcTMGPV6XMeDYrNpARH6m4tdNBKBYObgOTME6rXGZ0WUJnONHpyOD/pBdeAg9i
kyoXgU1sJgGgt523aN3xXIZDibm7aIpQGrdlZ5o+PayGzjrm6P2lapb89O0Q80NgrwN/0oqJCz/H
WPl/iGAa/UPYg7JyrdKQ56J9V26LWZtIH1+bpz98LD+KesWOws9tCnLnXGcp5QCgdVw43Oi7q6N0
2KYtfojeF6mvMasbdk+EJJ+p4ZPI51UlgG/JAI+qpihvD5MwbD/iJV3nXfYLSM8yYRdLbiopuBa2
IL1ABA4BSHLk88daE4JU44wYpotuNcKhKG2uVRptt03rGj8jm6PSwOX3vB7mGQFEzBZAcrltjVYV
t1n/HvV0X5I4w66wXHEEQskvwtgN/fUl2IOOTtAPOERBWEoJMkGl+Dv4Vyqz7VVQZy5UBOqI19AX
Edg7nCz7ib0bn4ZzwwbckP91op3vQLRSr5pbe8rzHMJTaUrCKcVosVhBPvTB2RTJmRgZZb/d9qKi
soXaLxTmoVE4+gJIt6Gd3Byaw6qz4UfOofKebZho/KfUssfGD64Wkk+62WWjkQIDxLxEm0SxOKjF
I2vdz/Te9H/PwWZYVz2nTONqqFk4noeMpRMTmBdQ5FpVNJSxO/F9+h8OPLCIELpH01XeEB+3U9Ki
bxalfO5N+DPt4Nm/MNbj2a/PnRoNf74/vntA0wF4L6kKTcbE+F7HdirxURvSpMAzMwXWsJ82uaXt
oCBENCqWM6IFrsgbc8hyqgmvLGJ54NeE0x+KmJTlo736I0sfEs4+QdHxO4mYk6JFu2EOxIATLwXy
7M7cTTBhWHt66M5e3KhY20sAAHT4DZagbj/XCdyNAAiYJcJ5umxCO3fsrBifJ5BQM4sgVdl1Ap0c
8lGUISFpeLmjRjl57Cwb0WFSLaS2WjIY6bMS9LiGhWCMUEDAje2xay9Z0yzeD9Oz/6DFSjFx1bAd
o7azg/CF7qMNmY61xJl5j0mYeUA6W2H2zL1Ajs3SXo6JMXDsq5i/TiHLE6Lq2OqQ6TmQakbOWIyI
rT+Nbpty9PoHx9+QjZZgyI6zbzejDQ/0osd4s43L54XqOH1viHE9K2EP/2z+CWj/6jDwQzuK0j9W
kb242BTPXTR3ItLy1lsR6d4if3T+ybAPBDJtio7NL8MBm5Dbnv1AJbT/fL4XAeGu1ByE7pRNGZm2
Pr9WHTdlr8JTw8RM+xBE8DDRCQQB0vgo2943JNcuYR6xbNN3yV+/w8ZiLe4+566DISE7soTCS8Ac
AMyGI3qxiz7iSoto1IN6z1RhT66/rYAoIH9pAgGKxJnxs69WTGcLolVH9ojgBfJtey0sGGBa4wV/
NxAw2U2vJY9yOywD+IF3J4+QnlpzfhZoVLakvcjS6r9LCa54CHxVGBnHB2MVaJgAmMk1pe8kuYQb
3Cl2GhX5AZvyCGE3ANLFM8fMHRdH/f3gkOzd25CtkpgvYZt4/+NPqcNQ8CKJ3L5NXhqKVjjifyya
GY52ZyoyvyYDDhE5XjiZF+33b92PPm2h8TpICJr6qRWBU1q0FgnBVluRyXjLgVavA5FbmB8AxKAe
pMCqbRCbbxH2MtoFvmOuA/hPnDXKCANx3UAmHMm0JrqZlvn43UsjvfesxB0yknKvH7Ps3dKHbWBt
t9OdQ320M6/ZtlGS+bWDnQ0u1R2xvA/RnBeIk5+D1oS9/uWACyw6OXcjwzrkASZtXTo+Su1N7vzq
5faEUWDACWO2MB4G/U55mS06EyluZE30JCT361mmXFgaIDh6t78GAZwEaqKghHK2rABZLu3pgKLd
+WG7ELFwycic+c/poqMYwEMF9dUxvexISlZYLDs3w2h5rjAqymDndf5wAUV4HAXsP5PQqYGdnegL
fLNHx+8zGHp51RqIohL5IUB5Zy3KBjekqGGLuy6CJMng3HZzzVp2tJuQLtGdd6SsiShH0qupgGLe
MDcpD1XPS3FtNQHS7jrXFkuEkQ/HcS3O1k/BG36BHQGomRcdJ3oPf1aeJEcWN9MF2V7ZOefuwkTJ
Rv5B6LvSLjubI8TlkzGFQL5UPBsS8KAlnAMamRLshexrMJeU75CxkeyVb5fclRWzV7+/Fm2Wc6H4
ybYgvqSTx8qFaDW7IXBl8Ye9aM8/dzKopV/AIDJr+2MXcwPKGnXYe0rqB9KL0IZJJvZ3eZ9PR++h
BFlAOY+QrdhW4Mu55wjqHfKV+Bsd6MzGy8e3DvsY/HlWICLnHJIGgujVF2kJbBEsdodw6tl8bUpR
3KqTi1cEY24GRZKyV5Y9hELF2noYt3PG9aC2bukpRM/Yz3VWjlZThxF/AQhRfQNIhbwKNRjFGRbU
eczj0DpPwqohjyeGlaiTQfyVvIBIZKUlGLdiUGg8/F24JetMVfzZ/lp0KrNXuTX4tahEC7IZ+Rl4
I2VyLsxtEQ94tFO2eK6IAGM4+G6a+jNXB7/bFvPX/Ynlc0TWY791ktcf0hNWJhIB37A6yF5BRCQM
WSLozRcxwMQKhwb0RaTK+wlcMWYEET7kIJiDb76mzxoVkPPxlWDFNCPNGdqmQ8o2CrpcIzkN3wK4
bBIxk5gmeWfN8rfz5NWc+9/iI1UhAIvSGTmD2z+/G+ns+Yn3NYH8zcjQRb+/79iMmvaq3L6osXXB
esIgul0v2f0QksHNv5HM01DkaumifpXYnEByVrqmINVbrETzC3Prr/+FPOoyW4bweaV/bPxISKqS
Wbd8OpNFIDXGNlbeT/iYHxs9NSOXRMEDGUPu5r1m7cRhAPEFZX/AMcklcTL9GA78LmNeWZYXJ1W8
a7zAD5jjLd4JXuon4XoD3eCoykJwbesAt+rBbZ0KYa8DyDg0xzKA4dJdXSfjkHwP57nSHsovzSub
W7+aJe69Xr19VOK++jLYm05ugcJH0PvBsgVs/n3YeydqJmlurZrBG04wnhHviJkVj0KfsJHIK1KC
K+p/Nw1/E0OhLv/yev8gZw7nwszDoiYcTwagq3GT67D5wf72jxYbKgqtn1QaWW+aba3GD4ETFWDb
zfjPUzpbfziULwIpZtZeJMoINAYKL/qzBPibfYbw+XgjjL9wsySEC4jiIHcjod1Lbvrkj/4p28Zu
1zGj3+QhwanRhnxUPsAyIa4j4aER3dq4972VHI9r6LdB4KWV9Gh8IKESC7F0yLi1hWXDvNEZTWOq
0v2WJFdJnyisH+tSy1GsngkNaKnWKDCzyhPGrTzuU4YFXIE4NcHGgV0zM03u/v8mYHulmxmshuk3
rxXgRYcjClEjliBPVfXmUCM5wwc4T8DxPpJ6LZToacNDux8VcWmk8S9V26IhtyTVI+2iHzAmbLUz
NcQ1mEbVe4nGgIglA3QtfwuRdtDvo49Qr0gTB4O/Vmknb/tou6VJ5hsgPU6WatH2LvHFBzjDgBnC
4WM9WVXaUdNTU78mESbzgXr9NmQWfoom/qSvphLmoLrIwE73AOrALg0LnfbvaGzSHAfRvZE3TZ7w
dwvUmEb00B8AYTXbx2Y1AqyqCDZUKsODZvN5tSw/KALfjpaoAgpl8UL/+SLQWRtaH+xFQdXBzHC+
WaCvXGi6xaNnlrcRZBErTuCOey2XtlDzTUagWTMx4m5fct2G4QQU911i7Jcu7BVpao0DJZKJlaJf
+G6gp9Bwj0xVgNAeWwp0hF0K5gmLWoF4ZQDLfBvSp19HNmisaT7DLarQUqxouxexVam7sCFba8ax
8T7tHSc8P68/jGsqqFeUybcG4MptxjEI4nW/giaws9jjjlGkbM7+cMdZIchi9dJUugnv2yX8PcnR
JCz+MTmIlmZJt0r/O1nedEoQ4v5hJTmVG2imBqBuTHW5DwreqZosMXA3RhNGlGhV5AieWNqVmUBd
0b0cOGy8H8C5OCCQCT/S5ZOEHYBDKwgo+HCMzmhony5ZLnX8nRDBYPZVGD4bX8OrWvkDdZ+vGLlU
9iyPvldJMRMTWP2a4Gh5CC8ryodTDI+ru+T1Y46lPbqxPr6+GSFE8mKk9CzOHRpVCAaKZzSDcRG8
NbRRpUT+k8gInbx9xYj9j48AqPOiAKytAWzhin7oMCHjvTQgm+Sx5w2CLkeEXfr6YTJGfWBEriUd
Du7iOXg/UBrF27CxDnHOLRSp1k0y9u19v2KKi0Gqjd9SNE16i4ZWel7sUwWEx15vI90CQXGGwdxH
9YWmu7rlAMyyoWKaW6z8DDUuWqPYR6u4lHUXiqgSG66TtYk/RZX6lXu48Hy9aQSPp2KFJ4+EQmtk
uUOxvjmeZ9/u3gaj6HKOz6xIGP5U5hWd7YUJmPwpUyb9Z/aYCvWsNmAXSiSKkARJp93/fu7Vb70q
pp+LqoqVQ0D9pASDPgLKhfqgHxDEdzjkwbxp5aBI6A2vpQpUMBqy7sVTiU9oKB+5jMl0HOEhkgUB
b07eg+R/D2lgh0WlV6qoWlq56AJO8354vazzvwNf9CWeTXPKAhTAMFJaJ3VEgmz3cdOokZAG0BdL
GYDIdSu3Iw0bnjvM4QiIjApxYJwFEy2JfDaydHOd6Hqvu3D+vjHIHoPS1fhUdsi2GALlsxEpf0l2
Vr07XFiOIhLRXFHcKXdxqzuPuDP2GLSvf0JcwZBrdHP/OUPR0zQGVEioaJ0O97+51cetL78WHEkH
ZiroGZnzlhXJuJNyHIkzG+uRiFGNE5Y+IqWjWsVZfNnrcY2HQXKSXxVzJ9/xZt0LWyohZQ6soL0Y
TVfpKO/pgcFM9dVi/eytpTjE5Caoi3xTpRrsYFE2zGi5aVTAB76wushLVlVyAH31/XB85aZ/ldVm
Ye2gAS23T88/Ugra8aJLryU4qzrblddXqLadbH7tKUrNV63XlKCGWHhKfi6TD9lW5e7DS2Si+uMX
SYyNrQiyGgGuXitkoikOWq5Va1suc4mGVO4aTYYUlwclOaAy0aSSP1jgDs24HXtTbjakVGuTr3FR
/e4kUAyTO3MbFrXASrsemkooMUhF9Hm1h9mSXiLfuDAnutOxghE0beIIGuwrabu8R5tkByxNYaRJ
G9y6ulaOBjqaCkndfz0y0yWhXxHJoMBS6ezgDsa+HqGn55zseoaEbijRUrO0wuQffE6PdqYuAX/P
2eiYRRL6NE2/t4hFtrZ7C/sJ1/5gHaLs8LgcYh0fPO6ysRUvKXf9+Iq/6pLgOeqTsvoXpiUeRen1
/u3W4ZvkcssLQgOxtE8qWY8Hqvgptd1Syzk6ms6Vxa/6jHZy+80UnRCGjqO22ZTWSPdkU/mzpEM9
B6Igg3q8RxGqDqKaiac984pb70Adyg9zZa30849Hr8Zun3KvTkHpFUagKr+I4FYijmC3QqT0C4Mf
QFM1cTHfRSFNGOFO4rukeqA+d5JeMcmcGMf0/8oGIBMGVnOBBS8KgYOp6b5OjHDuivE/3xS2UhaG
AetEk1U5IVDaOtmz+iN3gQaqhXsGZADAm04RZPie0LJp2gYhGcp+QOljAESyab/09prTMnYteoX3
AAdeiqV/VWRQWSbfaNqicmWx0/SLd4GynPmtNOnCmO8lDf6l7SwqYLCA3KPN1SwoZjuiLqejM4hx
9Whh+x6KN6Glz5dv+EJJ7dXbgXxXBXpSfSjF2UeCg2HrfOgJM6C16oIznVT+dHsG3EA7MQ4Cklxb
9iYSoeW61FbM2ZZCRCJKm6QD1L5jMz1TeLXNHm3+kTP9BJWOQ+0Qb2x3sU0oAU1yFQi+jd+0Chg6
X5WB9cDptljKzu66t1ldKmKjKpjgP3EnfFKBgL77/AME8BZPI3w5IVYkzPaw4n3KQAzafTEfZUm0
bAkebIttH5Kox8JjRJh01mRLUPOLessf0/Ln3pJh1STR5QMNjgwvNzXAeoSio5Xwgv7BS734azas
UpkvdjUZC8HGbSR+1GNidro5e+STWwrz3hnp6lu+alBuDgN9syySUqJPiIZ43J0Yw9UITKn+0t0n
F5TAkmYmDpQIDUAP8k6eQnnR2iJERQPvb7+rvFcfbm8HNbg4E6VjXg43o8mpH+tEPCmhzVaItm7J
pZFaZePjHySDLEJ0oYgcY9OIA7JkEAPndBjgn5c/Tv8YlF7Xe8MUE9ok5NgZLHHWWGD9Ik8rm9au
B3pA6ZjXFdDUNFlM0cnkpTT4t0wlxewmhOj0taoyhDIuD/NgYiPoElW850V91sIZahbkPVPtGdNG
qwSviUzjhfkVNEIlkCS26/EIV0KKtTRPuZxK03AahWmexYqPkf72faozJqYmdUosRjv6HWVZfMPU
mWtJoDlY6sXZ1CBNbdex92GNf6FbBT+OHPay0qviG1oVQ3b5s9AnUKUv+r2LIH9nLz93xhUfZ0Y8
1bxstPwL593JNSJgFYyC6zTFmkktGUq/XQsJoGKPgbvxGPZzUtOvJfK8HL8kob1EFuWY1qn1Aq/j
GTaeUKZ574LCMykbSHg3hnSWEHWsL44K42Qp+ntEhxtB/WHsARl6PcEecSrj3a/8R3kmBTlUTT3X
pieZP3dBwsYBtFmQHPx9GOu4jzxQBsYpJQlAC27ziqAcxGNLJeB7xMAXuuEvwhGr2uvuEFhZkYaB
UIatPmJTOIIvtduqjaXUWdbmUIRbAOU6zLLNrk/I7h0z5xTCXORBI/BrX46eSimGGYro5wql65Ij
2aAzUS/x7TTeH1tLEyyYY1oL3wKTr8lcIWQ5pDM10YSesy9NdM8LM+QML9/bVGJxQhdZkoh1VE/j
hN3NyBK0/cSnMABSCpyKqgdQ3pWSP4GWGOTI7KzM3Iapa6OfqKUK7uiQFU1si5gbB478yNpYKr/C
HjABqHhVOs/Vss88V/nX5PS4An2WBM07EeVizir2xZRjWBBQshdgbaE7UyFXjl5QWynI6fLzD5T6
J4YXjJUP3g9pBMwln8IRuf2LG0qwv/pMNj76MacUGBtV3Em22z5wcVM8PYYiSfilZT+Bfn+vQTs9
O4reSY9fEevTolOMiSkikSRI8RRct7gQSWruBNWnsa+Op34vP9IiY0pKInCbdzCRiOHsrkMo33e3
I6fXqmUOVNNPt3PcN/NER8UPKK+DPhK4/Q0CoCD7jKoLX3tup2dzywmsijuLBvVNRNX/xi4wbLZ8
RulmYy2q15OqUBs/42nJrlcbc5Za5QEr9esaruvL9OKY6RETsXdcLiS8a8AxgAo4imSPg5vgUK+v
p+/kqBBUBQ8JEYrp7ah6eNFhvTlKIJRD0TaYFkZRFyRjXlJd2fFhbiHm3cyTbgewTApM8Ac5+NHl
Ez7pqaaoQ/+9o/F/3buglvS+uSNYzCkvR0DMVhyYoD329arFXYAWyF5dYqr5aeWE5xnJR5UHPoC1
r4r5aDFV0CnwXn48k8UWvaCe0C6TTgXWsnIlzkLkNjVJyFYEbaJRbdrzMeD9XTxMwUIM0MAu15gF
u1AyuzDy1ZuVWEGcR5tICGgeCisZSqv2HSJwnTWb87WhcZk09+cUg1opLu6KhkjEWSuliE36yHXn
Ae59+xDvKVZF3V7iUXigcBWJ4OGbkhcLchGrwPmQf/qihTZB0yHBgJ6EJ/10X5ONxrxs5yIdfh8w
01iH435Epw0j27wEzGmVNPPsJ/y0XmFb60DiCWE+jGM5nMbRaU2+XX4hIcHKQtugl3u+IvWgi8iu
ZnnB3xUPuYGGnFmIwmkCWA84BVSM4OUC2YZjHaiYb5g2MrM4hXFC1NY9FxhbHsBopuA3Kf9b8N9+
hfo05xqeAjVBilNpiJZ4RgBqgJN5iIujziFW3ci8Xgu62EWQZknS95V1zUzWb1mYLn61NT0wXVsm
JUoJ44vKNVUY9bYYoxq1rbdq9g2sxDkGwBjD5NEY+O4ZH+kohO9xxBrfOSgy3swPPk8Vu6mZT4tW
vcTyrE3As/vrYaXUfDNbfBOzGkB+Kzq+ZdTtb9kjTYFJiKfxUdrmu95Z9yEH892ddmXr/PuGfohw
DR6C9BbpqH1Tnr7iqz2y9IDDyYukLDVcRSsodYzaJezEZuljmrb9EXWKfEq5OyE3b4FywczuBWhV
wYqc2xNgjuLOvgWQ2ZL1ax6A5WusKq2YUF2Wf+7RJ/kui9aRu+JxZ5NKAlgpoltOu+mInsN3RCkL
TJ5fcoOOjWxQ5TmBQbzTkHp41G/Yn18x2xc2qhX++aPbpoBkxsLkd2AratQc7bxfWiA47UUgd2ly
51QgqtrIhjolq1boDB0tp2nZwWLkG3tMUXXeASD82xk3apJSGWb/YPmRQ9Ec5rL5B5YYZQBCIRH6
VCdpR3VVl2eOsJkQCdUT9SLreY9XgTdU5wVh1rTpBCeelI/S9UOhi+gfYZpImuIqaA5KCbvKaCvG
GZQYU3ZeYe8tfZhGAT3FGn9cAJWY+wDXCxbtmCW7soXgdqSI2VVmLvU0tAgyFHf5CEs827ZCkZE1
5owLehm+4uvF2LlCoNJkqA8Wv7EPlBINfvgPoCfep49Ogzj7fbLX5m1ugc/ASWkllbKFObGAqiK1
lMQ6+SvsOe0aE991X3J5fnMaBbpoJREsbZHIuClob3vPTDogl5f4Nm75YRWxIRWwdukpoU7GFDkn
z6+K6bBtjuZDHttvR1mC5HJe0xC5NkNw7EU6HTNJxAqJOYRxxszYrVliYn9FEq6L4PomRryJFkO1
DmLobzYbPiYov3X5M05bOiBfZyRHzOuefWAYyB610PeH92uxG82n4236XHp/LDosz2Vid7aGbYBf
Dti4NVKCKnMdprNx2FbRrIghcRKsEbkullDxso1C4no4r4IQWViy0IMmxV6dZMwEYncBomBg36o0
NSDvYspQGwLY01K94UJUAZq7ZMIWp2O64r0pBDpf0ApPoZInpGoK/RED6CX8JuRtaXtosIfxGERJ
SZXyU4HZMMSSyzspnx1RMoDcts/0wHS9oUekxW2hHE3DmtJYTe7Z1oQjzorCH4c3Hu+SKPIKzQ0E
ib1hnsA8wJ8PTEqEOzdgcvQ1avPTvaOr4lECsySnI3qkFRiXLE/poC+Q1haHPRgb/KtP+7sSyMLt
HWG3sPJJuAb/vA1uyz7ejJSDqlp+s/T15b6gaVjCC573fX8J3yRXUgp4K5kcwu08axW+UYcstxnj
3F9sb9zT2x5KzH1tw00ZN8nO+g7eg/ICrPvac8tpRiPC9g86PK/VBSK6ZNoUe3PwlRnX5zLzQvh8
U4prrBIEouL8xrxgY33L6YfXrUdAkySXwfIwyGf1N2walTn9M8nvwl1M0SCWQrB+ElC49bOEoBfF
/Afu+JMbNFyTG4jMhGqz2kMA4DiwndQsovi3ntcDYcxKgIDdvA0q9eAYKdrsnlNEyX6UEDpnIUDX
viabroPv1mb5w5krY85s/PLSz8vZXj6Y/IwwJYKqlaCJknbTPmeBR2U96T4Th2dmXzSvoNNOgsY3
Bmhp23SWt++Y2sZ39/WqjFRvJEpj76OWIRiaAil/bPQKFEgz3V5xcnkAjixJtZwTXEvQdNl16jew
dDSq1coRbNu8U+FCyiG+/6HWSccakgRUZnxRD1XxFgjfbhKHp+SwDfzsdodGcKHCrrfsLFzZeLiU
mdRJhn9kUpIaeHzspdRE3yqnJXtYtZ3PM0Ef2wFARNxTJjjJFJ3ZZXlDyF+FK1w41HnnqEAl9boa
fxj4WhLk8NzlD2hsrrc71iov8YvSEFd1jitePNJWLYT2fk6//LZQWFVHftaXn1teICdhsOLiK3Up
OlUn1qRvIRZEZYxWp4FpWYj6/zKYYK+mfrE5u4+w5FxgPTRq0aoQNEfz+y9JSMDIIInpLxzXJKHG
c1kmAtYNdowpp5zqMDSflS0Q557e4u8fFKvX73E4vF/Tpt5UBL8pTqKYSoQtv7TdTpOd+dOkj+Hn
2WvHCaqMz3HnyprQulbCXUEcSrFZV0qMtyb9T7nP4Ju5nETXGpOhoR8I5i6Fkj8eYYi3h1M1NBc9
9xmtD3aLjwCBvSRf3v9fSbaiNo0Er/FEfcXvcVNmhpuTMa1A2baduFE9+Mbjw6vYX2uuh+e6IqR+
JX9Mxk7WTBrSBkOj+7ItoIMkGvqC3J9C66Si80ZEwe/NJ70DTMEJHCd7P3MOCl9a41JpgHlZVonC
QCGWMFlGOCxMupFcIX0yoYx+78568diiq2DjS3JwGo2u5+hXPZtcmcJRKc9JL/3AzSV5CFYTAZpm
lZRgcaWfkE7UlL+x1KpFRH47y+cIaSWGBzc43MG19MtXx9jFwPDhIwpldxRXCw5AwVIpvV/pvAph
xD/AEfBfsqvgYPke/oWwsaQPweOjd5GHvUbhH0NevLD+mqFHdRof2kGdnVUJp0SNlFBCcnkTaMr2
WO+r+ZgNIx0DQASjgwwBPZSmzk1jMNr9zWPKl5CveX/T4yy2Q0zVzJFjXp+PNRnxKzVUv51Jsm3H
urXZKmgFuMmTnMqGcxxSYO6yvT4ASIUcVIq5f85TkpuppEjbOrEebb80dXxEOpVLiSjC+MjivD5z
f6IIQKeaYUcZOkZqduItFH805GR/zYwzVIPabKXQEgvzM7/lFbBQYu2czM+5Qkbld5PNd/FSDejQ
hd2G8MS7LnpKAeTGAFaxcebMvY7mGLfGiIk78046Obsv5ulJApFFkdy1Es1mVPctpLOyOfaGHIH4
14hngv2qM7w/06rGDviHCKrreRu2Fq7E/kb1tliZ37rx45Y2CGXffZIMxy31UwALHDHVR9JOC16h
9Qv8bfefmKzp3TRWOsk37np0SYM3Ui6fpY8CJzFssE9CNRUiOlnRpE47bfD+X7fDKc75ZsFoy/b/
FeCJ9810co/VDAgEQe2uYAJ485+cG2urbAmBUlxaDQiOAzhgfAhGx7iHiPjdbXiuaYn2JVmPbKmV
I41SaIA4HdDcxOOstXYlPb5F50JacsW+nWbW7zbhYFF1fF0Y4Ibtt068XxCWzIs6bV0ZU/DWrS8t
NrQnoXAtGLo36QD0hNZ2Hmi8jFJlE1t45hJPHVv4Qa1kB+/vLgLDIML62wYEAYCZaoxHhof/jW63
0Eslkqo2j/Sfxp6KWt0IkNQHqcF4N3BxTrARUqbG3/X5oP7OTHQxYnzOiwb265Xw3qTklhbDDL/S
EG1YWnD+XjKRUCySd84k+5SEdSmCak27k8434hM1YaUpwPywM+X9cJccK2BeWDoG3/+1VtUnJfXL
g23uqD67jRhX5WxKCsRBk9A38LLaLM0XvFZaPnghzp7W0CmN2Wp+tTytsPaOir8lJqA1f97/wv+3
7WhKRPORKRmofb81dOqP8ZFMmR6kaJrOeFR7T8mDg1di1yjd2KeCKa5HN8Zfm3D3Brp5sktX47eF
p6YlAvQ78uu+zMdbMvwlNtH19xhw5YZBA7ucZNzatPVfZGer8vHvAJnt6wDZ1XRXCB4ZtDJme556
aygnERvwGjwzI/aiGoHM7wD46qExG5Up03zubY0zrNxJcjooi4bW99TjXpggR82YXcrTrVOy0vW8
9Gz8Qzna5J2DPiUwiHBFXICpFf5CQuIm4nKI9xdShfTYFJXHHXi4n9nMrvXBTnD9MUYa7oySYcsZ
LLZeisQMu90JURh4E9mEjSEkAaceC7f59/TvImgiiw9RRLWBREvoHC5uCLilLUyDLFNOutZvwf4S
YDv5K9Bhm0hFOknEakuNqnQcIXkjR6tl94olomJ4W6L+P015nPzp5NKORTzn4v5umX3jBYQuHr0a
dWX0fuIrk4GTTcRHUNQzoVt49o/jkTQZbyXRvF3EVn0gSdgOSyxbCYymBBN/BNpRWu9wfw9nwkvm
oum4JsxhGBQEYvAx3p1dZQ/DpzuVZnsTauy/mJQPKpVqEJomm03KpZOm3HSSxI6FUfWuL3omoNoK
SgsQMDVfw095gvVt4QH5tmk99qTychP6LS1K/z6hTFXkiJJNmLyskXTptReIBGY++gfxMArBE9YQ
k086Wh5LMmdILfAehUhSmfjsn5Ze778fVfbFDWU9W7sKryeubX7D4XVRxYOPbXJPL6yww9T47x4y
mu1OhaXmjOWhtjFvokN5rrzWLlLjNdE8b7PVabwA5gEP00MKHmmg2Ukes/RWcpjd6sh0FY5QosRe
MDiK/P1ohRJ6dMp/NxVyDb7n9I7CGbpczBHSNEMlJkuxcA+9vplhvva+3dVuKUaAJGIw+HxgXYJ8
k0M441lwyua0Jr+qLsFUNBZLHOKmrjjwE3dnK7d+VUiOHwVRFmaNQgP3LSzoF07ez5JsIBMFZfIG
/Mv+Gl3mo9bX1kGmt1kqyUQYjhQaqCwh27R+tM3Y06O8yRpA1WE737iQtJ1pfHeDg9x62ht6Rvpk
blepe1+o0GATgYi3axHfZm4tze0b/IB5uNVra17YvKfrSy6Tsj9X3FIA0cCkCIqZH5sE8dHrE2pE
iLJIIsMfsMCAOGrMw5wvMRMmkJptuijcAl/9eg25y7VdTQj1bC9MVlVOwjCiDXD4IaGcSqWAnA4i
uwoWeWSffbQqe+8JW80yqcC8c6WkCKpLNiTr1VtxcCozWmWuWIGxEw894oOWFaPtL43h8Zcdh80J
nHYWTr09OpvN21fsVlb4WL6ur/c909kq2xlv5u4Nn8ER1/xzPM/tzghRCE5HO2d/kHVlRLElCVNh
3ZdeSVwzER8Q9cp0kRzLfsarVVymMsyWcRJMoz0mYWdU9z8/Trkl+e/sDkBtdwVM/nha6FD5wk5N
816+VswfRXh6FINjuzlCucoWqTvCH9LNZxtymiDqFPT8snB+9mpWYUKEFC4q9NWJ7aeyk19TezhS
4pHGy9/K0o0AEpqvJCHE6661fwsML3AhYo/AZ8LC3k+xS+L/7HnouhzdRAGSxYotb1XF2dBTuDue
ubn8CpomkSUcwMnAj7MGBQfVJ1IqtADhXk0yCxo/xX6gOYNBdyDPplqNNrHsGndw0J8fMduwcOLC
x5e9bJihXSdAyZ0e8/mMEEphWVZvA3u7DKgqw0UcCO9oqJwIXLm+aJ1+xrZkjXdyzLyMrWZgk04C
5E578DuQ9QEDji8aDFG2MM9xgMCG8ZSFJYBVGic3hrMRfRW80+FDSrpOy7eReWZV/HetQD4/RKhh
aWF02f2NQDU929dW51NGMkdfQs9sWtlnpoGEtoOEPsUBUImdr9UvAEqpcB5/RlO5+sY2Oo3f2gLq
2A3lDV3kOskeKg5pH86lKuxyRs6TE69MIPiOwyLhhgqPETONnhrGncEeDDT9YBsG7tZlByIfUXSn
VFQFHZnMe3CzmR/i3qeSFajAl9WRYfb9+t7rwTr//jRTnBTRFE3O8hMPdpmToKNS9VlJT9+pMAub
VYYNH8vTp3Y8jyxdPE3T/WsfWxOdjtbLSu5XGgOYp0cNarRpYWxUf4OE+2pqGbWGn2G34C/krzkr
FXE7gbT05z/xGgkDCyO98+LKJDOrmQWlfSaaweZsVTLx14p17dqdWbU38LvrZa/ubEbVJYBtpXce
dgmkvUkFs8zwcy3lC3eKvyQ15DRTsG3rT55oL2WFszMAB36aNh2CAmsVeqOmlPt7mhz9XJRXIb5f
cUcd8VRA6zllxM8anvyvLb2iR548loysqDZ3cg+TcpbFJ5iP5wtr92ZO2Cfs+WVP1K5yTu4jEsnw
sZJlBaUOpat8qTkbUghPqeFvPGk0aEu5UI1jvRNuBoyP//k5a8vglIBh01fSuPYkyjraAJzdnj4n
ZBXbcAK1jQ+Y/VQIkNl9+YhzInRXGNmIoCe/B86epGCr7aCqrn3ArkdmsGowZglY7OZativgd+d+
qeaXInW5VlIIG39GTq5mkxizMkqf4a3jKhpQb456pACGNfqfB6pvmDsXrzQrB3FP51t/vPNnOAXq
XhVFOCrWgA/uufWvX0bOOh6lZIO9SO8bxTpReZB6IHKyjGqQm+N8YSQbNbpev/doUYL34PXzdvoN
aynCETRNnDgeHA0z05bPUj/OepuCNXQHY4ciQMoz7ut3pUYbAWr27i0Fp2QJO0DkTkjjvnH8eWJC
knuCQTuaTUQ0CgzRg6GuiCS8HHGnKB62jF6AqhCf1EqDxOcsh4K6fA8RmMqNJCYCPFbPlp/zpKwS
lGvyZ3nJpUN+SyimhHK+Rq5Usg4eD6RGQHOco1dG+J7uVObId86xWQ38b/bBCFshy5nVQZ11bJWR
MzbYxeSgtk3lfe+RRIPDbOvaG5RfWHWmxZeVElqFi8LdvlQVOMoPbKXKiGnUoBaqMSrU0B7YujE4
S3OukGnKtv7H1gNRNVQG4s3MO02yng3cKWStEvPxshilj28RW/MfddcGX5Hcy/Hgd36BW2VEae1j
qrKjbqGRXSr5QVT1+dH3mMGL1vEyZml+sONQautAMH0aWGJUUy4rvh9KhJWlE3E8o9MJErYSNccM
mNSNofxBBeSUJoVNe/Ky26qdMLzr8S0Ps/2k3mpSx7glMYCI1+9c7VTmycj1+zs/YzJn4C5AKVsQ
xWo+QMRt0HLieQl5RCClndSOMeoqh9fB04mZGJbdI52HPGTwTGi/u+xLXbbPoXVrbQGazfw1DbuE
IxVDfl9u6u+oywZJ0RJ5yiy0b5Y8wQreLYfVw9BmMYe+6NAEdgWGFwTEzo+eZ6fr5q/+6s0EldWl
w4wFYd534nHtSPYVIR6s1gthNvw/kbczuIPwlQIXvnojegVM9VW6I12LK2mRtHvUwBM0JhwzzPrK
IivQUjC3Gt8OQ+U1hwcs1zFO76bkxuvL0bN1kH94oMC5AzUmV2DfKVx/S7c+9cVgeuF9VZdYlFeF
4yhUrYNJavPR+4aFstffTX529C8Pe3KoBclHbun4NAkPUafUJv1ys8o1smQ9c+6q4KZXuSOfOLLy
F5q//tEkLB4HGtGsTWxBiG76AtpFsmNaPsBXwh1M09oP6667OLYTYZ0xNMh/3ht1fflLw3dlfd4/
aqSgznQwOAtY4KeYHfSY7ih+U+W79NBKLtN+9fQtmDT2UY4UCfOEA1uAIRgFNZ+/C06Cy0isQThv
EZ6rE4DbL2/i/EnbNT+nCXlgIeYxdOlmF66Cyl2a6pmjj2B5iFeX+HT6gvLwbYTADq2ugHIQVgdC
b8LoQ2zLEZUWXaePEBynqlgFN+sbmp3g+LOpCn3IgFW04FCW22B+Jtid3uRoMEK9CGZ/2LTsIG26
DGrXTu6qL3D8B9xX4vlSnXs1JE6XingC9JRPOdm4Cp6lOJvMTslAXF/Zd8T+3QCmYp9YVK0mXrg9
8PNzxjGCv8pD7q4rk4HXaXVKr2jbJaBSIPkzn3KbFelEZZq2QeT1t4fPIYE8mY97n6sFAJeuU5xk
LgN/8u06GLDj0zr+wfjaUlX6648sssix31zsT5OnfE7RnVSwZcFpNnRfhvYh43zCBgCM906ZpcD9
OsyrdQPwRcRuKsiFezBVQmFqARiXG9xFaHwlTkfNrEZQGRor2E7Ixa4u+XmEtIdYIIrtwOviX8e2
PNvlPkzq+vd5SGTYBiRcJY5B/WbH5m/KlCSz1dDN8VPGUNgU0Gu1kmaIwWa1rMHMrh8la2MZ5NUc
8f5pqY02iJ12bGh4LYQ+rjDQL7qCHWyTfXEcTqCcsUTEqaToe1iNbbGt9X24fvrC6oP4dpIkB3uM
hG8fZSKlxSNrgLEkZY3cX/f4mpqWjbWRxp/4u6mN+mu3tipKjXkuIL2TEyWaNPVffQ4r3FkNXfoa
ZQPY/3pKx+1ryRKy+H/oU4z5AInQTouanJmnmnJKiEyrAQKXcq1/UsDAOCJCmtlioxcFmaPt4kAW
WFRkKidd66Xreh1wJc9e0p90xdU/F7Bpo2EuDrIUBaxbm3Hk1aoBYW9d3Jf5Su1r2MMPOAn6zpZm
ZwgMWB4ZyTtHeP0ajCye2zZ7xQ12jmKPDi9HouTy18OnL59lx1Z25nCzQkWD/jk3D6aZeI+IEKTX
rQBce0I01RaNbCfAMWVTEXPIhQBN5VZ9WtDzZLkmZYX2tJSzqfgWcmT+P5+ttex2SUsCmvb8v8Tu
tR6THbIjUh5ulvMXkrxq8Py6he78IkzH+qnb0tTpCW/pptgmYselnQuiZDHrvsrxvwm/ROx7fvTA
DSXWaB7N7BI+PRxcpTMA/v2Y2pzG2uti4boUkqqNxQE4e54BPEg/tq/4fecJ3Lg+qWfBHxz8W1Cp
WtwbkLev0amd+Z2nY91PqHJNckzruZaTLT8LdQyN58X14fFTFUsabc7MHQfy0QyFCuXg76MFs5gY
lV707qzbGbjuikxS9VRqiE0agdpZMCWBl0q3afacy3/IRTxaZSXexX9FedW1x8xfKnBtLvjDdfdi
jkMeatCTDqm/l+aeRQYQUeEkVS/6B/yuq+55GoHeAFwU0q/axAArkk0quzcY75L7BzeeBGuSYkSk
uXfof03t1Z4KPvxnJqO/nDPD12JZ18d9WCRnwCsgu7nNL/wYJUz6S+qSyIm3qt+gVsnMFqNL+k86
5LeFrm4oOz3lhhVydaMUfBBFOg3jmxFk0FJOsaa5Qw/NX8ijMfa9ofhuduJJA2x7XYMDW1gHy47N
fVjJMzv4N9Gmn3A1Es5oGQXY6NjF5cVEaCcFN/lElIAmAUjZuCGf1wA7zU2nDpST34qQQiuJVEk4
msqQh+Ua8bX71Oon9L8D/YAsoeu4zCOhJHeno6PG8bR9QieYT+zkq/t7ZBqgt5W96pFcvsoVamit
/nuKVS8RE+ARUqfPmM9tZOyoUh64s0JYJdgKnD+8o3QvHI9B7dheYZmdjEfAjmp1WuJbujlR64WA
L/oxBXf8qh+3LlBI1fSlSUwingtkxDfJeVbWrycKgvZTvoc14DEWqT4QS/oytTHRJ3Vr3Qhh7ega
CVzoiPjvx3dBgf3Q95y2I+Vv7UESBwK1hpbh5qSKM8VoWuK5PQCz5CSKQKwl7jpxesZJ0UP0cBPz
n7TIBjUp3UhyWKkOauFzldGZGt1H/Tup+BDIfDSvdPzuFTLQ7KKfpMTg1eeXrQK9UHCva9eJ38z9
HBSomYYL/NO1r/0kw0Ka4bKOml3YJrRjgLCUQTuprtAfnkV3iHOZRoBG5b3abg5Bl2QS4jasDEuq
sHqpuEzAJaG+YKGkkRa2d/4eUccoH7jc91bTM3FntEdouugOx8svL2Aytkf4USVmMNohXQwRY8SN
tfAIFVbins3XG/napwcBNqNmg8Q0yBLzgngqW1dKGsl+eUsBblSnj2Vm+e4JInHt1h+3tytu3Syu
mHfkY1GKHpHDbTZAJRFQk0cqKIUE0sWierpTiXLyYb6NUhEd432+NGtCLW8J/CLUqK/cO4M+67Na
e/s2Jq3x6pja8t6izJt0WQwNIOp6NJUvYL044gvvT0gq1TKNzpgNqDpBctW3ONUia6JNTNCfNgwd
SKoVpVVjPL0ovkDMmOmR6L6EU4ByonQQakgfiqUkEkK/Bg6SWHbXavuQBpwVqkjRJ+FuGq8f1jG2
yx8MuSpMhkLjF+ZsZaAsg39JJ6EHgfp3aQnViWKxeelVQL9V02A4vBC0KQKDnLO7B3h8l2u5OcB5
FsGD9GO6mppmWUqhrrfs1d8fb1ps0sz+iex6f9AjZ6krZo+jmh4DFHnwYw1JwsrJOpgl1hQVyTz1
aasentDdk4buUl9MdupsapEMpr98nTzFKozndVBXkc3xBzefcxcZ+hH0Kwqb3yiGvbRvpXQyPLT+
8Xf0NUs/tGQbDk2BN20Xr7LE53UAARWIq60Chnhs0qsZ7W8bMl5LF/c+uZ9F3aJod4wdCUjIsfUz
wd+9yb+Ke3a39N/e5ZgLRjdGL8mofwfjbabTbWOfzmB0Dtt2Rxf2nq59ADrjz91BHV7FvEO2m/q8
xvz6ktDEp+9eHt0c5Sv6AfD57dYSONqhhVguw8L/Z+nI5HcZ12tWIUmzPZM0E5doo0lUMfeU1lsy
Ubabrzi+VrGUut74BzvxPJNlRzZQX9TnWdRyCQxqh7ZGPNUYYCldCQHh0WSmE2UMoSFLB5ThFUIV
Xos22xoqdYd243M884nnc9grn8rL5AezXzJqOu4iRywfHSG62FeqQD3ulNcRyLYCjBzmkPRLpbgd
CRBJ8pElVRT+Z0SL1T6qinadr51LNzk7m4K0xdb5/rbq59+xYTfhKSH3l28Cag6JWuVh9Pvyteo5
4unKdbEcpxt0hkw+dnNZYfMbWgH4NnpeK1crtEcw3Ffhy0NnEJRzKCOA+m/rOfE2AZHQywfRRCwV
l6EN7wD/HV4sRM8MPW3BbQNQ/R00yEhCFCZqeGUxDIACWh6ajQJ7lBkjpKVoJ175YKb/kUwiC81D
B9YsWUCGKU9RjX/I5f44w8VOCT8EQFxc2WU6IYKe9YryLzKiqYmBxfsvVrrEaRgX64PXCwXAKhDN
XoGlZcll2gmhoa5HFpVt3WAWn01dKXBu2EhARjHner53iidm03FKrB9r3ISFuBxfXT2lqkM6QvR1
kZ9MMlPY+xJTUDdSewlgnP1zRW74XW7eSh6kqlITuWjXQncOMvf7o2cUL+M92F3I+rIFmh3I+xT5
LOqps2cTLygGNyc8Hy120YXMf1lUUhMAqbvvwcqCyoycV8dbGKPVOcrrwbDdwKKtGQUKowZIYEi5
5DaTAixs1oBL7Z6qFUnLrRLZFfKBu/JmAgvAPC8tlErWLjNZGXDFh8vQ3Z+MrE2G1WiCp4SIzuPY
mjOe73m/cHNmr9VV/RdIrmqT5fp/k+K7ugzcGprViXUbPzQNSy3ckzrzyUx3FQV7K9BxzRhTIguB
WCWUKjTvHn15/lfJrwlyew9XcNsRfGQfHUcNEjF1lrcJ6arEpQluOV7AY8v9PXQ5qE1lJT9HuQJa
K7/02NHGhKsgDklRBWbkZhqRV9ezjTkK5cf18EcN5jq6NTcy1TZ6SX5CCgY5jHBPhgMHBzxkJPgJ
1LZiIsUOYYNmQ0UfwuGrdR9mnnwiOI5XW7QkIHlfw4/Onr5HiBzODZA5/rn7qOba9z2Ho7VTdp9n
ySbvZafJ05yZvKA/7qbqYrfqXHHqjURwEAesdJvUz5j6npWGAwNMcSuRtvTvKUZj/MIb3yec08L/
uRnnS0i+0Vqz9BJQkgaTnnnyu/6s47pJrz9uvdbZF9Rf0/Pcvqx1DcBHnK9vJ4OAc526w9qYZL1/
qkl+tkT0vVai/6eWD667N+UpyNTWOGlw2XW/NNQvEtp2MFc+RRv9LtSldst9fwFhoDbM1iD0JxSu
1XW7t2Vvhrjzx6QvQJhd/Sm5Nq2aaaOJkXn722umoYh1MlC9GjGHT/jVpqjGn6DNUqbLlUZ4Hn7a
HnjK6WFek8RYauQ1+92WbrDkK47TgYOHVStQoyJrS31lXmi6khYNZtAjVMtVFbKCVSsytj+Wf6NT
ws/NsAj6tmOQqZHF+5QMZ4/08+krFaDwwz/J9VRRRbV7WidZMG81MF8tN2Z8FAsZgQ0geiCkIzZD
teajfZHFaEhteswA6faxZklSxtG91l/Snbrz0boMUyw72SbBebPg1fn1w7/cAAjTmbiFUfHub/tO
zICDoCGFBAfGaT4XubL14P0PSvbsvphbZRjzp9OP/Ih0PlmdvlBbaTyVGruhtybxxQZaviANlIK5
oi58vidsmsaBYQNp1l/WVSLh1DPMKbvZfYwSANbFJeSt7y0gSdLXlyGp5G621ZkU6zsU3sVWhx3N
C2VrAEIpDeMVdcL2Z3rVRDVgWfdIoOFN0OwrLOP+DRmcUlvoqSbLBy7Q462+pBAfHPp0ubLGuuaM
4MAA6boIqS/E93Z1EhNIJtUbxFvHvQ4IBfUJHoWCDfolL50+wrA6MBOQ6UmCCreK4I68LSrc83y7
XRemuL3AThe9yRoJqKgtWVJQXaQMGHVgD2wKtT98wlTFfTwsq+cwGnTeD0teqBb4HRsLI3Nsgqjd
IO/hO45aJQJK7dRSmcPiZKZTbbsBYz54RWp1QF6gDJF7P6J1SWMpreCLkVp6t+vN+MVj8E85Vf/Z
Ejg/qpKIuMl7/MfVqhPCMP8Np+fYpCFNixePSOZr3xt1yq9quYzPog+Ad3YcBrV7Aj22LKaWFqS6
/ZZG+aEswSDS0xrs6IHwivtMTyt8p0jERsVfGSpNY/B42V829RMMdx9tpkhJMrud6b5KzT9vhgY4
9uCPZCS5vd4NXJUuVEGLWcdWoDj5lKW6NhBSQl6B9JE0xZPP0jw9yfSrXzI+Nh9X1SL2oj/sjgC3
3yS95p84YJpu5LDvL6zBrnmtGoocMp+RxCF6oYyGR8WZUGgPQhIyhC52FtcizFsENRv8VNc3UP9G
m5Sou9HOoD4LMZ/r8nJ7GoLoUC0cbI56cwkkzetxgDmhwgW49wmGYbA3qGK1uUWrjNwfNDiqThva
yX3L9PHBsZWlYZyRpniO8uGCymOlLJ5hBOAQgPHSxoUxVgz5hbRk5ujDYlBLnGInBurKe4XC6jdG
2ZvcftTyqHOS63ESVn2Hec2H+AfL1mD/0/D5ss02YkmIMCpK6jt3hTB+BSdM5YHFoBCJCDuGaSGY
UmtPT2q2YgsWrkOCD5Fhilmq/CRwpM7FD8xLCQ48mPfiuCF7+9Dm1SQpPryvuyvfKlnNh5TnGIDk
UxQdqfpm8QtVoEavLso5alE6N8BPQzuzyoBLvpXEvx7cGa5Bx6FDxUbzCusVX+GstdpfaR2hmVs8
fW9MgOXCj9TlYupb29JrolWpk7R8PnYZPLLI9DmFdFwImKsQweWVzheSRqHEuX44+gnDATi7YLNa
cwFRU908ArfG9RbL+xMf5C6+wghRqYjfWpWDNCuqoihb12BxEZjgVhCi9+yKKwvQLp3PtFDAsarV
qG286inIdMyz1fu47JLemtZZsVyZU0kWJLvQ/fVyWWNWqZNvJYkOAMXivay8LjCCATLYe3yWZPDY
z36q+TzBYJcTN/L2XDUVgl+tE8OVCh9dwX5TaXjNM/g5+/H8TBTsKuJImVj5fl+uN4jIesv2gvvu
P2asCtK+WMGw/DQE/cuSho2GjKGz3noLn2ypvBp23W6S5qNARcAlShrOz85AUumR68f90vhAoY8T
tshUMJlzEO82Zom7Pw6cmWctX9+ENYlpSzbz9kxeZRDK9dV4u1MKyjgVplSPNydy3/2BZWQL8LHo
dEyJz2KoRddwDdYkdeKagCRmThP/2mvPSpzCZmQ1DdqlZLM8oX6a8UpsOtOj1hiVd/KC8YgnSy3Y
YwxgOW9ebMOy6aTpwxkNj4P4IWjwLfgG2C/GEFU1X6fyoMSVIGPWjGgX4Rw3zvlOSoTjqDOe33ei
Gf8d7dsIm4pQaj9jJ3nOkWCN0JfwT+Wa1n448X4FwJfxHCjqqIIuZEuw0gn7vgrsIf3qunCd6VJP
2xkOK+spba1b3unCCi1a19K7VGeHOGegs5d2TuMLRj8LZCXDgq3Y8qTFiWyndnjtA7RaXDDfLSmp
ouA8auJaTt6z3llIfPtfsHFlhEa/aZeL9cEz6Ps/qzTbLNKw9JXlsUgcfHdsepTf/DnT70tVL3Ar
vk8lWCnamKVF4sP6KnFfNSk0FT7bysUxybFw6JwJOtk3z2ZsFdxTHlT6xPYpemE8ICVEd4B7ppQB
sA7N6QPxCV2BmmGaFyn9OssDcDi+w8AN2P6Ym09SK09P5MkKbJ5fe8M5uc0faZnytMMgpGvTIE1R
oQV5GFbfaczzkpYGSlygSiwFIJ7je+vcsdzaIvd0bAUVHVPz5Vx9iX+JRVyGbiukzHyuETuseThd
X3GhJJknK7D3QunWoUj9T2dObR4/opJgAZfsPe5HH7U6cEUg4KP6+YbzBtCfBSgYWtISsde3pbM3
IPyzohnO5uycu6+ddJJu+clCnUfsG+7kKFjbpqAKlYsLSU3OBW5MZzbM/YJP4nV3Dy91UhQZvSZP
bEGUg5/EAqrld4+uptbqCPGEAZK6organax31sWabDS2jxaLhrhy/G+C9bdwVm7pxiT3J5zB12D4
WKPBy0BmXYw9Nu/1IH926HeBAh7aX9NKM1oVEzvYUqhfIhPkv1KTpqbv6x5rXcU6Kx3RL7dSsCcD
z8lp49FWmC0/nkE5SiUbKialgIggE94hUFgyto85eX3nE64yHPy7AralQMF114NndfvNzVd2J2rY
I0Lnl6rO2FdsJVgF7q8z5bL5lmMTU5kgW/KrtCWrjjFMoLa0xsGjUqlfyxxLxLPu/z2Incb5LjHv
c2mBJ7GJIHzTGxybH++0k2O3Dme0JpmJUZdAdbEveH1A0zEEmZZJvrSjFL2btQr4EJXeK657GkTK
WZz24TkioYelE2VqzNwPTxZlTd0sWbS0K8dD9Ahod0dMu0cTw65ZEoc+6Bq37XM4AgrOt326mB18
0qbbccf1uG/bq/rt6ynodCgd9WV5/81VX19eqy1JaUiYyaiSf61lZqD7txfRGH7Ggq2SkF58eo6c
w3WWVhUS2SZNH4XP8MfMXK7OtRhPisS8YFs3leUmDCk6QuJnaBUn+Amo+EN7g5mpxEj/vx3uoA2U
1JlIGjQRWMHVaZjNiKmyRFMSTs5FXOUEP+pN5yuI7w+Plbf4y9DtaY6u8vAUqmTmRNAIvDR8wShK
PznnQLkbM0NsabUSQvpIjCU4pdfpdLHSeEaas+rS7C/I33KcMgF/BK+/y8U3MtYzT5NxIrx3Ok6r
tA/XXYsBik5JBZvrf8wcF+y5k32XxMDmTu/Rkj1EEE3y7PsOhkwqoa5dLEyZvCd/5qePZaZA3k+d
F3Ge/l0OGjxD13jLGhxkOITnft/eZyceNYKETnoH8SF+MAOHHIO9vUNHy+z/ViR964bcL7p4Ccy2
HMlIM9mpslfGv+6RtPq73O5JC8hntj08+K0w+kWTGfUNwZZe1cOoYG62/whUiJxIsdig7jbpyJJ0
7ATuNyKQEdTbKUZjrIL+JceZ8hBKVaVtO0C2/fKkwigbdce3PwSctGeya022u1BNnabdlp95riQk
Dmdrdsr091ZQzYMz5xoVyEAioBGRQyPxVQc2AVplEcIhr0L3NFOUxlirOPmD22BGfNmRPLK0C/F9
FiTxRTlN83V9BfFVq23V+WbFCR5tRIgUoRZfony2QlhBoDsUh8kk80MYMD6qSarKwn3ylhfPaF3E
EXMNUPzeXQO1iSZ6lwWe0wi+iSbwlyYi8UG89up/lHbANrgsNm48Gk8u4+WGzsvSl166UdSAhTBu
97HK6lcRQAu+tbZcCjNQAA9rStkQAvmOw4u983FTLdSqyUvKEv09DWJMaAzzrCSitIyqt8WZBms9
lB0SNAf5Mlls95/NHES7yZvBxFYPrC0/YcRNFuRzdxjXCWbNf1Wu37NYJZ7OemQZ1D0zz69SoEuM
e05k2gwsxuO2TO7UCf6BeV33VMPb6JuTxnyV4hJyj60VNAFKPOYrw+WoSqNHFGzACNdEx7svHf6m
g3WjefQW57oXq8+WGMQkfZ9r30AFr7Na/OB9twiFMLpvHPFWJHZ1rJmHCj4wgzt7qlkeAkMJNYY7
QeeDIBhMZ73u9nZjsTthii3N72MQUKTSlzjjqyY+D3OHjUue59bNhjBl2kCGa57yBPF7c1mIGFp1
cqVR0j+HuMUM+A1jyTdIPRBxR8oA34VMFPAnesoVdDhO+7ZrzkMrsWEC2wGorrLtTfekMPHss2jd
A9WnPGnBzZhm6F3cqlxagSbBGUrYJrsF78SetOXz/ATYxMIL+0X7xdKB5qrV74FVsy1Iwr653+VR
7+fc7vJ7Rvfv8yNo3S3c4UEaDeOXmfG0UTE9sVcTOLdu4nckCWnjpyNBdp5NHlXZ+ZJ1/B4oB7hv
A1GOw36PIuxdcA35PFqZCydWmKBids47sqKgvuH94bmEA6tixCrIcMMAiWAioLLh//1iVwasdPpF
kEExcF/hNxRbFjUo0npHl5eO2KbrSwR2q2RiUg2mtfmVS8CWAvS8zLOshohW5hDRQkPGDbfBLA/t
GDHVpgfZ3AHwCLWB1d1Cc8Sr0Ns4BK29MAiZYgiKWMT8BlWG/6spNJ8GateKVV4EJ5suQUSxJhSd
JMfd4UFfj0eLEeJVi9BLR8S+hEbeynWmBb7DbXnmP+YiUszTcmD8lmVkW2i/R6CUg9obtcnOvDHZ
sZozKb+3DoQexl18RTZJOKfGJgKc6fLZE7x/qXTGG9hRnR4mjDZB0wUiNLvJh1Iot3ek80bSYYc9
W8eIfV7BSN+fpGXy0dpQLNz8Ndmqwegk25Zi1zu2AkQZcSsojIwO5MFV+Kd8HLUmuDdILWqHDcES
YpIOaSZ0FrFevEOnU2ojzZj9LXWIKHbNdC5m4tqF8s+h5vN1WU3g4x+Fdr8HAVZdcJg7+HNfZJx9
T6G+36YhOtJfN+voMpF+3TK5eAK0ps/qvf++jAV3sQUnhK8TgrasB8vbnfo3MKSgQZGkVBW1T+3F
ZfMXONEA2sLwCCcrCZJEqZkDGgFsMBZvyd2PzO20LHSzvBpo/Hy/wbdZ47Kr2w4YbXiuCRxAcfdC
BcUNfBVZLpRH6xgQMvtTgdijStXnaaGHi82sYfNmpUon0OJHhDL1zonuwPaifPtJrj5WXHld80nH
2ne+TOwNtIkBDC8niVjg1KxSMNuqxuulFTumqyCDT2iDSflbGMC4CnXYR6NqjQZJnKQJWeZtoQob
8GYU6gi3LDH9s8xfWxv506QxiQ3cSbNeL9WucG46FEEZjo6dOPOv6gCuVPbj8m80mJk1nWAuzpkG
BnactaVgSrY/BGXcJSqRDTa8URdnhwE11RkizRAnqUZDBBAw0uTP1KahsZgpI4l75m2wHMuDKYB1
5f3mU3SPFsEM+kuRb4LmduKMUNaZeEpZZNP6bks1qG4KU0cNojY1xvIqbDtivjoahIVX4T42Qh4P
/300EHTHDl0Cu8GUqA9HO2thH5JwpZ6xsgDUTLrbwqdrtwPV8Z+rSn/0KwJd1c5lHPdtiyDl0XId
xdNDVmekHZYc6LsgYglCyntss+9+/dJfrAavGB3sbiiraiIXNRcPwes/l3JzgqP5w+CkNCZ+OLLp
UaZ0o2kEpk4671U/9HPGdub55zpV6TiWVf3zL3oGWaaBFKh/txY1c5AB9sau8t1rsoPwhja/lbmW
RznoBooZ5Mdq+RyfQD4LUl9CHDe7YmiJyKkfEU079TDFSxGVYEwj/nYbEpvqrlR/8hVSmMw4A75Y
3vO0upOczFa32LAYFPqUiBUwLvEgP70c9rUlaIH3aqG/jJ+3X5GGHgjryoWcT+rLee2ZPkdHYKij
Kc6sHTK9hQqDTOgonuaW3poUhji1mgLCyAYl9hyvjFBW8VfuvmQGCm3wS2qEmPEQJXAYIHHB7bO3
Y7s5D8SEqN0qSXqo30Zo9oEpmLE6rysnhDdMPahMdKyigIUxuSKxm4+JcEK9GwTphlSEJL0660kg
JHA7zRXms7eMYYEAwd6HEMFoyBxKImT3SSGGUstDxYELVbGXT+lP5OHsJ6BRB326Z5u/P8B7XU9E
66zqqIbH3QNi0jRrqJXE8fQiuZrtdIWQAk3tve+Ks0kSphKDYhC9tv3pW+wBF0LE+/2mY9Mm13GH
9763pDFfcNH4KgJaqGS/v+zyRUkQk62rCwVNvEvJfZ7doiQtcOiy+YIasAX77/+QXs8oNWVyCjej
qPmpTrbuuXG2Nn2kpqq18Y8VJ9X86JWXqWsEyJnpJamYVdN4IRQeQkLo2hxra9IV+54nNFPH7GNq
gxcL28uxbUAPo5S1uCmGu8mLLjw35jYyKC2Nc6U1ChvAVSM9sBVK7s3z0xB+I/ywrQQZ39s/ye8T
2pe/c+PC/509NZE2ik4vISz/czNgFy4KKCx/IBjbZuLQ4aZqSPEwWxdXoqcfCLig1WOVXL/nQIHw
XEARl7Hs3K2LjRzSNHLJNwEmslvndd7fsaUp/aBKMjfgju6IlNsrI1gX3QndQn9sOUTwoBkTSWdY
U/OoQgNNLUq5FpVI4LX8RII/jF0+670CEmQBpin4vXXkLndatx97w9YjkL1mqMuHnMOccyLgB2nk
9rzfBjqK2ThZDZ64zXVvvRRtBL/5ETQ1tc6fL1Ynac8s82tmUiM0kmQ31zhqcMzuisEX27uhNaw6
5o3BlySMFijFx9GEUAkEH9NeeuLsjFlmvxukzYjY1+HYB6/zxC9LkplwTxjTy2F7YiTbdKkRne1Z
+Xic/gfGutONm/AWOKauIl1cng95TzzGuYI9nfmMs47xEi7c7Hy5rutYqYngczMIr3QCVBO5pDok
6h+IBIr1SnzOWQVXVfPz0a3lJEbLlEkbcDWzI58pJkHwzDLp5WIJagGvJ9/W55ub4NgjKZHq9LTr
PFosDBXYogLAPVUeWLmGSG28XofVhjcWWz7gImzpDC4g93a/uRZe467VczgMFU1efCUt+NNO7Zk7
dk/o5V5KObDEBuMKYJs3u++WEi3BKBFBtM+VS9K+SqsIvkisMURa0VusHQmagJglttBy3AiTFxoT
9u//ejAhzyyWj9h+2JT9IYsS5I2nKiVAdBlDcrxTUXfTDisdy9pNgWMbvAkhZsIiXoZiiwrJXwvW
HJWcJawqwG/+Jn9CH20x7F+zpLUg0JNmDvIaCd13Ol8bO7nMh7zfFNdMW+hKV68y3iPzONk5F3Mn
nOBbY8c+w2iLwj1yJAiND05SaBidMcgdT7R6w1a2R3odzTntXkRzu73yJeQgSa5kC5plB+cBQPte
BWRvHLDi0mYyJNaIAwN76nq/bCTCbQGHALVJgoMpSTrZHpSsSeMX9FrDWE2XcZRzk3eMj7j6mXgA
jqgxM1dNhB1DcRE5tmw1AcYMY5tbfc6aH3AgL9V3jQBZNXjm7M1xRrjS2lNMUEi6lSD1p/6U0WW4
zfcy6s4Cyi0KsiYTONqYLM2Vge/DKsTI4HkIU7eZ1KPiLvMYxY1lZMd7LeEd1qMvDeb+kU1UvGqk
FCprfHyll6jxGhSlwdQVUr3yVjhM0UVa+K6OZQjKnWNR3QkTJTFcICUqRZECGDCRSdXH/4ZtVgx8
GUA62Hi6MBS6QucHpsBc0kO04jZLOVTwNTxMXy3gVp/T464HoIm5leKVqH7EVvbh9Z5BkgsTE2mG
47xmUwCU1m0QlGnMXff49XJJzkjQG2HfHcFNkmIozBR5rT5TBrLTyxuF3bdLkGjY+U9VMcLHYlgl
kbOf2v18UAa0bVrJQyHjjod5F/UlVRBMwaVnJ5CRmVMwxIyAr5C0Ayl3A3eK/aR4QJJwzFCMnfED
CqpEQAQ6M4XcnEs+wN3e45mjy5lZLg9njANtelmdtiL8A+jkqju7Icz6MrwePylRpWwESiVBlIni
ddPpykJ6AKbL+rSvfSzCB4GXV4lGxX0TtHZT0/HvrzQPGkmBXXAe4CL59yRt+VqCiKr6o05L1Oz0
bsetAN6IsykpA+N/QWPEFt/vNQRUU9+4iQlHMYe38yb1809Y70owH7RLYocsh+V/V3eCNj39WH0J
7VKvIOWC6WKzy6TW/YDhRVf9iKesjIxHJfSepzoA83gjLPbya8hWymxQNI9zt95C2FsYiSEaHIbi
YvdVstacLEuLefzNuCfgL20bxYpNLAFkJaHzzmf5GBDb7E9Vm6FzoQtgqmaJA2u5fky/EdSp85Xb
HZqB+GSMmv0zs5RH10eyiGyMk0nTYB0MqyAWA+aiL/83zNifeKwYJ4TEUJcudMALdLDaEWv+Ugno
1aJtfy9P/W+XLDocZrzCzbv0/uTFZhO8hS1GARe9Lx3qXeR1qMD156E55Z1LqLjfEsuVg645J63G
4YkaI2K/Ugh+0wAw5NvyhQ0Lj5eh005eYvNzN+KriRPvg053BkGIH/ZoL24gXY65QeAumTNNFkN2
3rMeIA9p+WMybyTIS7vTTqbS9U8mynYImCUZnIL37eBKv0Oyf16eKEe6e1qbQyJgNBp+tdTp1/pr
DI4eWSy9rAVybnGQScX98Q2GYFAxAOFPQxVdcvoZOVO/5SCtAJkS5AuJdFJxz813pLpSrvUyKnEV
BcNPKl9iJorO/DSlsTlU7z7+ik1N7FIIzAxipKIZXb7+jyedu2JYCh4mSyL9KRGS5BbGrlsz0smZ
2OiXslzDqWkNPbT89lNcBcxaW+LLiWQmbjGHPsBFkCbi1JfPaomh3NKQ0DivAHTbrXCWPFFYX0UX
D+mIJuMgwathjlA1oB9U9/d0eAb2hom9b01Ggb1NJPu9e3z6OBKQm1hVm131JmteU8cs0W3kWwfH
BGGA8VyYI8IQb8631JTo6XyhSJfXidMGNKFxfJN93VEjhTxp/9q87D58+lChw3YwI+TsUv5KuXrK
5/qcGaAUGTSdSPxa+Eb+/7YyEwH5P4aCROZOQYomIRs24NFlqQooeNvi3IjZ8L6fgylNirZ0bPSs
bKTfuo6eZHDBjCD2gmOqJ2qQYs5a+7gKYJOaU27yGLUmsuFFryOxUf3UtuZM6GRaOJgQM+xQT9i6
zAoP78OkacT/aijQjlt3D6K/WGXtDG07I+TQe1jfbZL0m78CG99MA8Tx7N52e/rjAPBO3FHqMKBG
9PlQ8mt0Xp6TDYkvwycfqhnwUN7pUm1XRdXyOn1S0NjWc2QibiwTQJWTG5dbaaILye3Bx2AMOUbf
hMrrtUfc6NI8jPViCrHLadkWet6KBEKyhT6+4+QPDmXs8Dq70ABmzKAotYjwdi7/PNWee3bwZM9e
JkfUJC3BwcKajWgKSR3055G4MWPt2FaVhIRX2lQZYFI2/YIeol7aX1vx5qPqAZNmi+skbwBDBpkZ
7O+rtCvfJnr/fwxP9pTBsYmN3btKKnsIwagV6c9DfA5Mr9JAab9OPFdZzWbDAUr9KKSeG+HfZJ+1
5iBWC7iQHkpQI60k878VZin2ZHXjnfs6JpN+K08cMHZpgTdEKSZbPjJwIOk0dwbrgU+ZJoz7MFla
RcXoiA4KHTK7J7JwQDuDpYNYRB1HXaf+KDm2m3sM9ZeN3sjlfQsO3HL7KkRhajTXDZboOOkk3Ux+
PgJdngSlFVIsHNCPat+OQwUMMBvCev/mtW7RU9caUu/76eoXKmQ1MF3QFTMwpIbc53o7oIu7e5p9
ZXk+npGvHalVPeaChCOpk8QnPIgzlmtdqqgiUDAkMKdoNzXtt2S2flcu8J8YcTj4fV9F9zLHv+kK
CbRsj6UsMls/Z7B9/Lhn8TGqay8nunyjH3JAPMi3ewH2BznLw3ccloTk+AQth2AdcIAJYRbER3wo
KR++7TnxsgRiGO0WCu3fW88+y8vLq5DldJVnvO5IlMKLrJU72b50yoR2uFfkMVm2poOdKCvQMwWC
KBxpzViicJof2FJYm3du8OQ1NMXq/wY03vbFBre6ym4NqoW+H0U1zGJ9THJL3DhquNSqfY2nVdsh
PhpjquVxr0ZX23gVFzv9E6TYSn45KTUOx+85V/TdjaHCjkw4ZQ0n/WFDKarplt9RN0j0/ZCsCBja
WnS+f6C+Qro/dXSrP1GkOKNZaDNiysBrIT5eRnB6jGUPdy8ReScBhOjX7u5DUNfWHijLsWKn4pyZ
D44ZNaAVlYJsqWlN+4Y0zhLYL6UMXMTjmsaS3aFgljeYSJPvFx/StOzbGUupdpRu6opIm5J/TEbK
Y5bi/u5ik66lCnmThGONZTIjzqFSY6bOmj+y+iKeN8Y7RaLptex6gd9rWaof2TdSxHcAlwGyQ2Bo
IFq+ZFn3tcEkujzkjgt1u5zAB9e6GCnvPabuF4RJSnfy6xrfqedMZK8p58ahy/uQCBHm5oIDETCV
MLmZZoqQgv2P+hOgQpzDGosotZ9iJIhOSJl3xfFur7gqfQ0o3ESIP2MPCrc5vDWHDdPbmWQhtmYq
TtF0q4RGBKWn4BT1g/mmu7nwjnXfg6268/ElEor0PfHLjQ3KdH5qMltsKCXq+KVjCNMNia+h1/RZ
/b7IObQCHT70YswfsAqsW0lk5bX0I5Ys4KND93JgX6vA94CjWAlQoed9u6QK/SgOwSASHoOem32i
8mRVhTrqetnPJNvwQ4KJuYSL0yF6xDKLxs50wwwGvpAkFNnzbtIJ5tyBFAH+DFyhoPVgYe8/jtE9
WiSYLUIT69MT0ejPiHmeMQMe0aoykvTyxn3Twaci3TessiwlosVNB0VI5+i+ZJYF1KQId0bEd0CP
lsWsqt10yETNT9hldbnHCsYzJPp1+LydQVCFNjEvngO60rqR7QTL0LTZJ2w8Vj9lTSxgKkqQGSUF
ay6lOKiDCNR4cAMtN3NFCkncDjao6pE4JnxNocK86Mddc57491OXhzOR18QLGdLs02B0ODlR/8iL
CRqZ8m7RDgTGXJ8+jbBtXJRFpKKscFihwaUlayviAHu65o64avYXgrxAxEsC6a/S5C+OAT+DmU1Q
nxlb4mCzIOoyUBRGu0AmefLJovzBn/StWV3np5E1liWhucrq/F1UX5As8bxb2N+CmN1TPxsFgTLQ
u6B9BjyhRf5u2NaBzfLTtq9mk8ucE8HcseG08ogX4mCQscZ4AjHxbBXSY1QjP3+TGWPHtT5+7NgN
bX0elzcOv0b2GmiKqpFYH22nRJAFt3KIGE2lvEgY2qf0UD+1+WvAE0KhKclwpMZCpDATl028+XOx
vekVI6DoPZNfTManVbIwcExnh9t6O2HOsNyI5WvmhQXN1vl++wMwn4T8NkVJSbSlYz0+ldm5uj7k
oeU6pCS5poZ8rYXt5/eoJ/u/Zw5FL3cuuxNj0H3m2/yoILy2H8EH1qPxMrnWG6owKRrUONz3shgH
18uIfUJ7OpYVit8VfQsEvYHCwrO7uCDxH1J+d6OikiN8FjcgCNP368JzWHFHQw8SdCycDpIIS8Li
4GbU/7DWCNFkWcdV691v4Lv2aTskP/UoI9cpXzSSXAa/bjeoywVIWc5cdDukXYXLaz1R+9iIPN9W
hVBw8gJ7nUtkNzqIbAOu2uvgeP0bOVNq/u2FI8fqJy9YMNd0yy4EGC+h5WiA3cZuUQY5Crmtq1LY
89KM4VPjqKpAQGSaE4eR24n7Ob+WKZza3ZaV5avgZOfLtQIUEL2DHOwoI5c5SAutxGK0JE65/aH9
DgENK68az2EkP0P9NBfUG1IhCix3ZIwnXzlsBd0AvwfgY0fpLl6vrmKeG/CoVwQkWHyOJUj+4w6w
Eyawp73lbElLJVP7b8B5e4z1V8EaDnaoeyXWujGm7ceaz8m5QmF3kUBGvP+31GcXAm1vRUnL7Mc0
lZgSGFDIL1Gi/WB71fGlO+MA3BBXTWA75OAkaytRitFLGuK+5kK9Aqbz/o6YDZg1gLrduunCzJFQ
yMQuYOcIjji0ty3tSyj7FR5pGSw8P3iIvqG9NtMYJ70IOLKI7QW31nQqwOF7rh545Pyl4zks14KM
PEBCY+MATpOSn/7tkv30yBaJROHwiz+blSsaIWOZVUlUinIvycYFgoeMp0rImrYWGEXlbhtY8e1H
8RGA07/hoXCdqGoeOPZ6NbLsl+BSv1Um2yaMQSLKnhzetB6HRwOMtRTPpXZ7BPvoQYnY5Wjd+2ZF
QzMNRKuzriTUWG7T5LWiKGEE0agjEA4bGePTXHbpxJU84OynLF/XuMwJuMHOivYdEw+LCSvR5hmk
RhkPi2jSgoltMidnaZndReki+hNx9EvSOsWZ/O6yFbuQEeGkiHj6ijB0+r3dKr55+FIX0E6zTfDN
S7sn7ToEXTT9Ra1mPe7iTgoxVvwszh3rPnuk3xXkkQnwUoj94j6ts4t64gqNjT6uKeGiy/xNk+VZ
DudVcYqY3iFgJEgjkSJswiB42ifiLfzvt4gtoahpZzrN+KzGBuoj0IACxPVBRipIm3hQzdy4yN4X
LQdEvBeOADwsd3BMpIgum4h86Sts4hfCC9XMkJftPllaIB8NkdrRGZtFa/PHtvumg7/VOzdcpQDv
Zkkg0kl0SmtsELf6jCcuZYYmsDXg/4bGDGj3pHGVlafUNj2l6Gb+Ta2O02WbjmXm+au1zOqX/wBb
h5+tfK6LhbdPbYHec3tlJusqMjbRz873FVB9ACejHy2xqVqjJ80IbJ6LYMS0/mMem1yP78IEEG+s
lblzYDRvqfk1tPa2xq4wQt3SDLgA5qKqWKTRVyD+WFytWNgf9GXVNGjjOr9bTyd2njMjLvkAiHhQ
PG8Nl2wkvdwXQjUDh1XmmFTy/e273hxa5jyR9gYZHIEOQSIyf5XfCpbzqWBinsYsgsSt7tUrPeyO
CKKjU5dOIVbe90HGfy5tWi/6WsAO041WNF7xL/k70gyEPkfg4OdXuWQFMRgSKsAuk2LvwYgZu7cj
J9Vc4dS7ngSocndFrxLduI2Cb1ISWxrinpbJffhCCs+4in0fWIgfrDN1YS8hghcOnZLxNxGvvDg6
OW9F3JNfIbcbeQIp1f5/ip7P13K8lGQ4Ei7hnPRWa3pkMa53Eb+veJ6d1lJY0+Y0ojXziFggb8km
i9Aw6nojHjhPBMdgNO4kw6NNrLk8Ghh7XVO3cZjGQ/PQbYzndZSGrCLzRyQoyPQLEtksjRbFQVfH
ItqEo/vcHsIdWv+SnoVRjBGNS6gX8Z+EuAOoEFkXxuoTDfcVAPgHEOK6SmWy4r9eERODboBXir9f
rQVMfV82KX98bWSth3D1KFiqRDPmmLFVXfyoXRUtLg++hRZzWtfCLNvwZlKgMhOuZ9+t76+9HPv3
RZ99XcLuACHKi8OvmuLkuJ6ycnlfzqDbdNJ36eOBh86Ei8EJNddD6Z+wRhbtTM5ghXl4S3VB0WO1
SqjIi/NHT2rj0DJl5hIwSNsau8lxUEMoKcf4PKFHK5IxWwcLH8sw70ggzVZSpTimmj2a6HSJmqQP
CxT7RZwnl34YNaPBBrVsqi/s9PIvlU8tqjTYkDBwDzK2H8r8KOkaKBHbZtMb4HEJKIHzT1H/mw7B
VAh0nk1nDB0baRAVeYBNKMVt6JC4zrI7rCOA9R6RiiXCZaiWwVTMkis34tp+T7oLG0HfiyMcbTG/
sZTDm1MBbODwk8oY193RQLZjmXFX7VcUxi1YTyJ3dK9wEpoP7fEMubSt/07PSHPrjKDG78Dcg9uJ
cm/yKo9C777tyKKBwHFjEQrYQgM+Lu+44fzNA7uEL0AJIdpLEu0aeqhURmWE2+34dMLGRc6b4BDP
YZILxlvxfTJjut+jNVmRlUXKa8zZnIuIAR55CyAhTYbsu5P4i1Iz7vV7yurabLHGtYhvx8utlFuA
86Oildp7vYxuHZ3uIMwdInEkiRsomFNIbvMPHhVivNG8gpmjyAKNrY7/QLB2V7ciy6+JT2geuDmx
TX17WKKyEqLHrb7oaIHSnwWKuDTVwAPcZA/SfrkTXLS12/CvdYqOgL832IKH/nLBDDTLXHmu2ykv
1rFxF7t+cagN6V/2O8FjFAC2XI4HOjIUx+Qs7OKpkuUSYVjcP/XcNf53s0FqNPLGBIth4XObJyDb
zNGC+u764WDriJJB4HLPVAgK50N/XM9zaQ06hQQ22w1UFX53kYavIRew4pnzGRQPVUrJy2dgw2y0
FytR0wTImQJ+KmYkLkFbmcBZPQEr3mX7juxzIH2uKwBU0WjnABFr0KTGla7osnVSzuKvNjk9gASC
2V7DzeIXA60WJhHrYxuH4c6GgfFLmIRzcNWlcVN3pRQLmqov9i7EYLGQTTd80r0VrEOKwMRhYZeK
z1QCIMuYVw9zri/hcEtdl35adfyrthjyDb2E05sFIqNM11xsmRVzfVEJrUXiXNHF+qjf2aHRiY/B
4AbEr9e9dV5O/71gQ8bzGsxKlLhkEcfup2iQak1/y2MtClHXuIDZkNtAC+mf+PYfpgc/S7NduOk5
n9ZQVutxxPiFep1OoptL6bA89XkVFbNfkpwgRFW09a7Q+mB4uoxg0CEXgE3Oodc0C8Vr73jGz5P/
hzKHVZoO0VYL1jRNqGqjMubYxiHdO2fDSmdpt6HHGeiZYnFZ5nPIYTodFydp7gNF6HsciP59v71W
sQsPsqfG5N0LKerraL6zlroU3KG0GWGEBjEHHUNH2MHyamjWYb//ZQV38XtHv4alGBT5JkNcNbow
vLAAoCe4PSJIbkYe4Mc+j6GN32ocg+mLW+2NvunMyxheOJZsoqykGJY9Q+lbwbwPkRepC/JBLJ0V
dZAQhhMih7EjMOYTATW1iDpSWOXQTA4sLpDsSP97/gBwUYW8d6dGlKfOAQ3MlBmgiPqsM4yIvp1y
zlhh+i5YZyDQ7+wWZFBMgyP4pjUIduO0/5G9qBGCP+Hkwo/Uwr+qtZcwproZ+u7lRAs7j1CEehxV
8uI/lWABse+uEr5k+Ra96ozPdCf8BmyNIKBzmd0AQ/PTdH4wtOipcBznepS+lnKc/VPuraELi924
/MI7wdPxCG/eVWJ+yxh1NWcVdTvnJUEFMmCFEp+dA5K49XjS03LM6u24zRLUfBuT/I1KGsnqgvHe
fNJ79hx+xHs5d6khVmeS+RDvzihA25YM7tuW+R+tt8WSrgcdgCXKnakQztWMqFUPN8EEVLuiRWE0
fV6eT/j7TYXZdWN2glrVYn6kyluYzZrPYfyspCWSiJfCGfJwDY99WabUIIrygIAMIjbw5SRb01rx
fgAtChmV5ZPMPZNebXfzM/8XdREhFLO9cR6XPPKLcSEL6VndCFlYYY+aM0XdHcZza8M6NRoUoOfE
yTbyHJoRkqZsq6G1vwY/M3Y9kpq46Cdle8T7H6plhG977wazJRXJ3IdCfiyB9XXCNgiwSTV3qxBl
n52Ab99zi7l6N54gZUOxmyss82qspwvmXMOMliQcf3WrduEKXuEznw40N3zakGO6rFl5JmWGOJ8n
QpYHqeqBpj3mAaf0LaHmxyEbqrJ0dUDXSCBOpeoKxNRR9KUFmawwIA4tOlry+V1v49Lc3NO4C0AH
Nhfo07O36uvF1mN+hnfaP0woEmUbgzFCncgRtOsoA2/YjUzJa366K1O0PwxdKdJ2XiP6WjwcPPZI
ahkWTOFA/L8ylQ00NZyHdiIZOQl068AitliKXCh4PNbBEBSspm1iVm/jMj/kbiSTAQsEEvzlW7sr
gGb2pR7BPi4mrZApRo/zYBRbwsMeMgenBgVzi8hK0wr4x65gcrd8TTBaiVIOwOPujw+6o2LstxQj
9oo82y5fMQ9CGhd3Syx394bscgaOgNAyUk8U8ACnt3rsTlw/Tcivb08v059sYNaiiRda7/BHUEZ6
DQAnCcNmKhQZfTxWmRWk7jgjNAJr//yx8mfgX+NnBUWLIw3qzAqP0zi08U1tprdITEFYdlXLg55c
5CFjJP6czFxs8XjA1SorECbovSygneBqcLW6Zf6DgE3Q7k0vMOj3fvzps1yp9mD7efYGphDs8XAX
BdC4ymboQdqWyRquNMuZ5zA0XxltWENOBehdpMhkBJv1jBBKjaWYVqKqe+cHdGZIluxN7ZT7dnOl
DGpq9D8yYTP+KTLeqRUX8FM7QfnZ963sFPXh3H5MNd4oKahQsMc8UcPcZLKa7ikL9XFAfnH5uScV
YoO8SsIXglBCeX+2LKZTHkxOZ5ksRZI0HNzdk0bkSPBMrUPfpN0UiwMdL0D5Cailzrd4quU3lKLM
mqJRrVYhiXThaYVBcIGAgUtIsrDpHydnVpRyzgQvaRwi4KuRFE4dPk5yfvyB9Z9U6y4UtHWCFuTL
5hT49b4YEpDfL0emdI8n3kaDdfBz1WypLi02gYAf0E0QN2LjIZaSm3ilJvjThYifzT2K52Gr/MM4
42TJ3FtyWWMeQLEsIDWHagUL2k96hNqts3CLN+HbHhv/iQ/2wDQllw82xIIkutRsPepdcgBDj4v/
mOt+gxX7E/3wQJHIzGpW0OU8jrfWC1kwFGj08JZi7TzHsG76Tuzxud19E4W9rRAUS1pgEuxbWkdO
h3QdKm8JuCR3+HufXBhwz/16zTTX2GUBhCx0N4lMJTa9ObjZN5NcyMpWBovBlkp+xaQ17Yd/39q/
Jr/TJ//1fzIrn8Jn5H/uo5zQeUMddWgj7n30xEQlRwnfhuQgw2vtX3b9e4OVXrB214L+dSGLqFVL
+m8FdtX0zhvOQmS6DxwoSYvWEL+vNOmeEnWaaAnF+150E1fRuWA6sU5OmXGNNmeMK+34OZaYj2Fl
6aQPIvFKASSlsZ9M1SvXY0LAzJfW9gIkuFiQ6uGZBGVtIncmtv0Qh+ZhSxePu71xLsDq1iIG2621
uaz09RJt4QJez5GUY2BZoWVy6L16x/neygesXRgKkYT4Vz4MBDsxYZtN2Iio340DPjFYYhh9G1XN
nMRl4jl9SB1dMIiQpXxHx8Gj7sJ/qNO3tmka1pv4v7AMH56ghVsLCkalwSRnJU6Ou+0sYGGOX6pz
oD/8EoD6NXl0tI+0n5sXIliMhG3Aafbd4AKyNxnU0PDiz3XaZns5m5my/jCgFTN1Xhy4xQ9jXnAx
s/yVKEnUoNtt6SS8CpbqrNkIuYoLH7vrgp4BH4HccRQAZx/T2m3b2B6YsndjvadTbZI1lFzCWHgR
7lJPSEnZQmfxGdVmSsdb5bkUjjI+DIT5YT11M//c2f0m1+DjyTR4MBfXW9PrZyUU3tBBNoHkL9lU
pHVN7xP6Iii6TnrRbk17QMve4sJug/SvMweLQXtIp3tty/QwbwHhOGQKvmzE5XWwIcDePNzvEclZ
Sn0I5uFbwf0I+bgbJdkMUAdTzZnCcm/fnsGU7CVDKOpZHwpXIdkZUUwOQZWyZ9hYG9Hmh8VRJknd
sdLK6cEHt4M9i7gDS6jb99U5oESeR1NesliM32O5vd4+w4D3RtoFdE+Pp7DaVipLa24zanq9Saf3
8GJoxr3kD5mImUYQrqMHs7N86R+bU6gX5DVScYUSc08VcWCLGEWYGqTv5OJNk9BwTBHzjE2zCUrr
PRPnJtedDxIwfOtpunAgqQGuF3mScMNL5F0BuzkEDxuBDOVLWc4qsoAekr+eHdIaJEWE6ZuzQEb5
Y8KxlhuxNSkq27BYwXBBzvyaZq6GyBvgLfiwSje5qkPrv1y94Vhqd2BSiG0tBSkI/AvYdSEkl1+p
q+MJwbWfLF1L7O60CXbSmgVF2fCat4sbUDXLOIBCadtCDS8lnME/ifChIPDggo7NnUHqXLAm2+my
Uc4r1GtEnSBMyTNKty4igf0VRaUFhDPFqXinzu1tS4gDsj+L3aTLZKvMHwuY06WJQCOhcqQRtV4d
sNNDDVuELXir0Rlyv2DLWZWpc39PDxqcGEsIKgjxzSUfHzmuUsNz5frGlq4Vsvunnra8NW7EwF94
OU2Ohg2pNDpiXlRisnAcOVaLayTSl/1Dl8P68byGGwZwbZBmmynG8es+F6MqL7EzylpBYFJ5YOhw
xV90fkoIfcJvTfQoh7UWcCMMjBRF46eRjPEXmgCaGlAvasX4AvvC8eIPllrbncFJhOKvMg/3UBmi
E2F6Wrsa1Xv9GNmtZYv7HP1HPCw8977uTxbojCJT7OXbVMph6O1Kl8BeJwSB1H9hP0uO1tyy5sAD
3LC0MSzncC21F+32QTLaBxbHkahpEWpV0UkFhHFF3PdfKfEi8Jj0IhbInEIvRyfA3MHS2soP5m/y
fEd8h97cTZz4E5sLDU2TlFJrRi0cJRvYw5Pmp2FB03CTozLC3kXA3kyf0XNBGix0N6EwkSicd3C/
5VhdTW9xowgziwcbkcdX/njDXyYyTSraGjo/gGQYiDAgWJNksTwRi3RE2xpd/N8f6Eul0jVvYFsl
bhxubo2CgH+CrDwonZmzHAcfKfE0D340Y5zIQedgKHNfODyWHP4xLXzbtoDHLthp+UiOPMYM6hfa
q5bFadf5qGA1QWrmAdp8XSRf8dqZt6YmE/MO3+ux9h8+85EHBnB4AlVhwExH3RSiRrIiooO4NnRP
osxvNrZq02DtegTuY/yL6aFXsAhbIlcxUg3i0LxG13tUegRkMu1DUSo5w8YnSQo0axkw1r+8C93e
0BZufb3YewatZFBmTptzfsSHkR7Zq79xE01hmQ9DSaqJsInGc6V89t/F4qelVdELbAXi/B4wzDya
i3MB38YzikHY7OJAjr37wzBm+nq5+G6G0Y3asBLQBVJafTI4ZI5i80Zpyz8FCJ+5FRB/m9ohtKfc
4TbzEZf7FlKDWbOA4A5BgbKG09LMVxPPYCPfmEtTC03ULa9Kaqz5gsDiM+SrEDPMFZ6LWxFZJ8ag
6ZLZdjUAYT26A8WeEqvRkiPU66huF+Pmwugje3WtjS697NKPh36E0Rgs0+kHnjOMOZpJJWdCiHnS
/8TTOsNTEgKjBCOzeMxnmqF2mvDt2LgKulmQ30n/KeonpYNAH7WfXRvwUqiiBLklZXdQZFVb/34C
4vjQiAysX5XWJfKe4xwZGttRRpaN4wHP29xhOYhbcV0He+z2wYjqRKbOOp2XVxQJ5qWD71/+6uQS
fR4nxp2WhPQ4RX0ml/JF8/Yspo0a6MXx5SStNp5dyB79jnmHl9W2TlHYBBhuwE22UB3lqPjDOA/z
iskrNWQPKSiMqXk6g+2nOiWt3jDcb+xzqQHIE+HgVYV+veCJfW2HuMwzE7X3k7SCsoQiwLdNb6Uu
l4Z6DUmL4EkzFovhLy6JGqd6LuxqGD2mF70KotoW+CA5dHIQtTUUeohJC66ocRbVt0oAl03+agC2
iF+Y3BhtbXuz4rPWIS6fila+HTPAvI5/OhInVfHOxiy80Z4x7OuAGNYzmyrKGE9UtB0roUEV0HF/
gZ6/be7PhH9MgEDcLdgux66dItUE+Vt63xsn46JXTKmyWxPfNjkXfXlHcPY+ztbrDAcjemokh7Nb
PmzESWZuoNhI8u1FVuVjPeottX8tSegSg+4KBZrN1k1DHNvEFrn7E92ACsUfWa4suOAHBLtg7U48
R9k0VsBMYRzOk9vIfqzzbch99LvzeW4quS/0yBOFKSt3kWF/WSSRQMfgab8hmAeuDgnS988ffBCp
WHIPqOGpFP2EMsvm7JbWb+O/bPvY55cIeEyuqYrOlfEONVEbRIIq8XhWr7RpJXEgHZXWh2nyh8GX
U6hkgOKcdizbwz62Xh8IRLg2YfDTlnAJrI3aw1WA7RbkWWo445Xs3i4FGj2lJ8lrOC0KopM2xDFw
jKhT7C2zKPbQ+oGiFjJWzTaiedHMnMJ2ZC60u1iOIJyJwEi+JmbLK/djDVXXcqdD6zeCnuRA+ovY
Ub2BAYYV1IJrEf9ky00Qf16AHkt8KuqromDGnG9XfyeeO+CJhx4eXpwshZqEHqPzdXNbXnWZk9uy
ugnxFAZ3yAS/zeufbsKl+93Yjx5ByRUVl11RfngoZx6mBxmFgjHC0Hco0Ki6Ry61SPQkDibBzVPa
r9ynbnug6xt4In2waUlCo2lyHkyzO+psOxJx1WgzkwuBhbNUsV4MvjmLFfnFi3dUtOECCi7yF4u3
BAB4u1UnJKE6UUwMbCwxXsDl3PhtFejbb47HmWIJAHALWGVrOaAUWRXkiFcFHZmY2soJFGjWZWDK
srQxfYFTZqvrh3HI6nJeyAi+gSvopdOJwh7WG7cRBTzyZjkQPlF4U3UCIAtyN6Tr9fivk8H5FCWk
hxFRJzCyqntbpEuE+L6Rxs/Q/jhQcMXb6CakAcJmO+c33YY5uB0slsG6yz5lYXJeZsGs2rZLUvUk
hHzxN7urwNWF5jtXfcN32vC4RBmS+6FFAyJSPDheYnC17unbe7+IEHH9GMh7KNeCanoCY4aBYkmS
7u4aoIYv/4qoC9iEAn7r5Rpz49qeGjR4JS1sW4/9D01ykzpVl9n72f5kGwx2MPtA2yHo7yNi8ISi
RSA/2+0f4U0m+dUX1fflxyHBN39nfkm/9+Fwdtq3L0KxPqDkN/pIcaSJPN86tckcB+nZ54NKWf/5
xNpKda2LslPxUn5tHMN6loy4Ol/l+tdQpnuyqoPsKbjbAe0fvwPOpPfHKWl07c3GLL6lk2NfsPdh
Igy4cXBycrFa5AAsuGYWJ1qZeaCJjCHnekY8GSA7c18AV25YAhJoi+aJahoZd5BpR/aaGrZ+zUm1
u2GfUm4RSUzvWGB/ZebvIRIc9I6b/wvYqm6R00pH01GwAUkqa9cs17dxXzkKv2QAWpKD3uWta1Rk
kfMlLRv5JtWSfrpwnEMr9Hjqq0Hu3PxaEIYN6JnttNeq566ZArEbz5bV9H04neoCl5PrDj0hV/sE
JVEv508LokssxFR7EQOQ8APkcu7vZL+2+TuodJZ0zAqoHe9AAFbNH31puj5T4+J+CHT1K/1PpWTb
UAqHqfAjOVNLYl/xZSERa7bSAN3vtis4vW4dMCHVaqq4Kc8hcPXrdR2MI8WdbImpU2S27SxCplC3
X+Mp6pNoOLb4SFv0KtbcLAO7/zk7sOAW9KEYIou620jPSpQDwgK8APDnMGviREygWR1vggePGocU
dno+XbOtmU8CKNtbDYJEbnEgS0UpZWZvHBbEHG9G0qf52xpRh+1YmPVaMKuql5mbY5AqfIt7Qev8
+PfI2ZLNzHXU0BheF1V3JM5IihmIHpQoEqOsf+XG6vxr4stmcHM6M2TUqQ0mHsTASAUhXJvjzOBn
ltGAThfpjjIXD652yJ/FTNTc8aGWPjmrOD9tOtsktbyD/HhoBKki//2YDuCuZ9R4V08twUczs9R8
if77MNBFunvSQqH0+wv71JSp3GxgSgFpLfSjH3EPX+ffQ3k3LuA12ilY01eVDkAUWNIWjB7umXlb
Ig2YY/AOtFGnqINam08PJTlaFlnEkvFSBcSEUWupugE4Oymtr54CalItGbRZL8B9hUoTzeKei4OR
t8nhe4cuKVnfNfst3pW74OuAQMHrSPCmAjf0DbCinoVcmCRTWAuWb9rJESRNG7QBPAlV6NPz4hUX
8YkUo5SrFA29yFP3+jg93H3rCYtsXSxCgwgPv9tODYU9+rlXqI2Hf+aOBNLzoBbbq/LHv0P4rbc0
8q7Qg2XZDG9jqjvXOub6fklue4zaT5HNYqNNmIYKp8qkQNS9p2tncpveYNXMfBWfG0WiEc4nua5d
SFdePbZgdBO7I2Rmc+ygksyYu57jeUsY29svEcp/PxRZ6Kv0BsG0PlzFd+cSvRcMNb/J3taonew+
WaOytfhLFPkKBr/a154q2v6Qtkpe/0qJQDq0QkL7ih95XwaR2EyFGLJT1ar4XGDvu9rf9hfIUIWI
YpDmQTwhBrew/YcVwoo+JP1nans8r0BTeOFKQ2RhrCZ7oIAcjSXakWk+504ELlM5XeXgFyoiPh+j
PHrv640DcKxOTQGbGp3iNVDYdJ8q3yABE+fOykLZ1Vm0W1MpahzWe7+2u8imYVSIBzFmQHdnnv4K
4Xb5xydK54WmKpZ30XCNF+B5zYH6dV5IXJpSHTXBjcmEBV6A6zu7s4XBq+eupX570wJGKp7mcsQO
6gPOZ3QGtWXgvvqMD2WqeHUHm7CT/897MW9uS9Hri6JMBEKrLxOhHNoN6WICqIKETFWhsQECM/Aq
Hun7ColWRSMdPN009AXDEJZIgysoYWYTC88t6rW7ONiwlR/vOOu3pqa8blDOjl3uON2othCWZytc
KOHEEXOX/9VxKq8aZBfyldWoVjuJefyyzICpZGHznLTaLqWmtslZwx/tg6QuNSlO16/EWvGtw3t7
SsJl01QRO0IyZ2Y7J4VlnYNRjPjElAfvwckoCwyvAbTI4fuEPul29WmfRsU91vi33jG49MWkTPk/
IIlneLKFW1SjDYmInuDJrsfKboSxyzLs3ef1O4DrA6XOrUPi/nPXkX9xjiTKfsbk8SwV5W2t68FL
40lrIdLWfoJXjBOtcSqZkusWvWYwAV9m4PDX+UUTQDdCQuSaElYA+sGgZ7Hm7A5gGG4ewWwoCqMl
IKYAfknJVQIEoONCDlemVFs80DZYvJhsRyDcgBpNaakjy1HezVSCsTvdNS1AE+pMS9EcTZepcrGq
ZTr98Tr1Grme0d72NjjLFFqCKfgacIYYXjWZIyBecaIZ66Ktm1/ihnO+/3tM4GUiGcrVbfLP+zA7
rnTA7oK/1GrC/q73dXXFJ7uhPhvU7oLxApxvI+K8MpeBdhm4iRwI4wMBYrYyJ5IbxAr6nJN4yjj1
M6adoywscwPGD+9yGdTrB7f260Ih6B1g1U9TOd+dMbQQYLEKDJ+tWdqxcnkIW+LR3N8t1luSmxMP
gCcnA88FQ93n/771sIe+dR2TPheE2bF7kw0rbdnRNrAKi0ZTh2pqsunB7qR30QI8sRvW6L3nJjj1
hPCRV2X32BOs7UOLvykFQYGIdT8vYdrg0YlzwrYNodlCMlLBhXPrl5AJT6Znb78ayq3oUVskG0ZH
rCLqCBypM02bn1mOV5R6qImKLxrtD+Xz7J/DAxmo1AL96fFRPhYSkP7W4UH4f0hsJ5SWEdRrCn1Q
YlGZxQoaWhIX58I4GEnRn7WARr7nmisbWe0z/mfuTj41aC7D0pN/C4PTrfby5Pr0o6WjmXg0W95L
nkxqE8bOCEc7RLvg5cBydzWiQfZlr24GeHoIs337NNdsMl5BVLJweOoi33Zppsgxdt0v8R6JizQN
EdT0fXXQNoWrvVKsWNRN8jKE0uR8Wh2xcSQcS5/bs143vUyIzsQbHYDv4tarzsyqEeDcTIt4fPsG
fc0uEMs4HeSu7mii6qFurNJkbts6u3GpGjB+p/MJyovWa7h1AaOLdHvSdqZ8APiJgA1N4P0/rZzn
nN+dpFGPQNSPbw6mBrnvFtBcUaAuQZfuqEooF+YwwFXt1cRPG6WFWsw8ogVvnizuqrJmU3novQhA
HlvTk5f/ExXkXkXaVHkYVw+JmdckpctFshwAQcIjX2OCOpxfJLg9RNNYj3bTGvbtRe7nyZtxGOv4
jjTKnyvQXDrhGvcoPFtxosGqJAfadB/ltKUbaSLdQ3bIUWTFxgib1TaPN0K6xZfTb8bJU7Jhs9VL
jIrAYh86SfBlgwjpJJa5fhh9gJ2D5c4+Mdfm4K3xkFUbD0PctvkeuUbiTf65ZMQK0BqrWHrw6Dvu
HzD7NwfnAQ2SzhOJDkJxm9nBkYfM/vZHFkbN1haCtT9Cmxj4WHuvehVBzPY4FT1bJ2lkDE/tBBtq
T1rY08tk4VuRSgJ0hipPLdY4vC7xZJr+ZeM7wZDpBRAA1uK9Qv9t7YFk5W1NK9aclfTArFqK+omB
UR9X8/9t6s98ycthTn/C6SviYd0JxwBLn9i9f2ZHeZCElxVuy3WLCML0Dn+kNkOR79TPCLsQQazv
g3Jy7VvOygpOSOJvkLW1XJ+hKUP9MkE408QH9UiusMcLqbxAZNSojLQsU0aMf4XlWK3H/BqynYnz
cSxF/qiLyj1tOmQn/ac0T7ErstVwHGQkbd/L1GOmzc3Wbxb2qZLss1LhI44Pv2M4WosV/fXzpYB6
fwrKdnDjpiDUxBAXXzinCgqW+c9ip2A+X7W0vyW/H4fUE2itFeKCDuTsBUCWLKG5bET1VSsu5qDN
wu0khB+osq4jdZfKDGo6qu4hL7aCUb99v1k/YLrmRu5wO1KIGQJtANZgvYwFrPERKtlgtgskerGz
AFv9i2oZ3wGJGwWgZDa3kLh16eBZeqYCTCkXLAWJPPOlwUpZau2Cv4Mq4Tvfpuj1L19KS9mXG14n
Bckh9rH5vTxLvaCqJBdM+Gd056tBCf9gZTISKcSPBUNppvtQV4JQJp7X8PXIUCJJpHPz7ye8YEci
wZrrHWmFOInN+0Q9cCZXs6qvlQbFN6/HpTfLca8eOSjHIE5gQAudITKAsjGvIDbwBrRkNpAXPiVb
GON33lezc5H2vTawvTOFkTRaKBQW0JVSxqpmsD9dqXbzwo4YIHesBUV37QIujorit9Yhzo/PdKKI
fYRjwSPuUKv1aQETdG3fGbsMM9MiJwjZslkDxkeM3TV52Y8L1XQWEYMSZ2D9Y5b+Dt4SGZp2L717
K826Zj1/3J1LtsIPBZaLqCymaV870bjd82iYjzliDotT0WVmnrA5JcwFD+CqpVDUhxoZb7yCYhop
XOiK6K7o0HMJZYVdHvK5upqwsI1Spgk/85ejZpTM+RNXHbKdbedXdysWa+oSob9l15VKtz91nUA/
yXPfA8VtDq8HGNOv8c3RWAYSmDcuDJc0q6nYGbEOAlEIzluhCMy7W+ZURI6wR8PzJ16Tx+REHolj
meazlYquuoXdXQsKmoWx0Ehan8wp53fl/rPNsng/BpyYcGl1gbx4a7BBJZKbaqAewEw6WTlhfnFP
yZM2xSXm15g3vlH9mAYOa/DPIeaHAVawJrhE9PXssKKp6knf+fkaaTiL3RlCF7m91ymCfkjlK0U7
aOqIgbp2Z4xm+QcDA0KP56XRcVhUV7oId0+74/6VGB18Vk7M7BlWV1L/VFz4M3VrnWwtcx3yogNA
Ra/kOF1ohEbPdKI3oJ6POmDiV6CzZIog9zvpFMvgShGWEw5r6u2MspyzomOGVAqqsEGfmTQzLxsN
Slec/aFA/UgeooeqLpF90ZkQ6eE9BLsRO1jTNdkIOJb654xC2W+AqbIZfTyiRBhsun66UL2Q53zC
Dg5ul7zY2ZrR1f/fiNBJBKiFWZlIxAuDYpb8mOmcrbzEwq8jX6Dcw4I2x/vu5emtJs9hYB24BNCX
3SAtYx8I5780I9D46h39SNHwrMgwUONUsHGoVU1DZNtAZ7qbMX65hmRq+cZc0pIu22LgCESgJM9K
0t1d5zVcJpio/m08eUzbCYXmI9Z54kwy0qsyI2PeIIo87y9D6ySQ9+ijohjdTqmsiTieXnMlrn6v
jvey014P8KTLq15JP+lhwUlvfC0EJHy4SgYH4wHpQG69+qxzqiiyNAU9Pba/hVaNXVSAKoyLwYRM
xZvVuIBq2sw5NUeYxQGKf+kRHEVNVzsOHZjzc7w2R9VT7Dko1LC9Q1IsCCUBtOUXJxsZFAmHApQ+
e4JDrdA+srRvQKm7SF7WpQDxI4JNWN9w63pR/Pq3xEsSevHWksoeMdcOVmSIexM0i6ROYqUsp6ar
2jotYhAqe0F5IMdlIvWQOHYKHhjAhpREtpTTX7YKTJEsrrzl5tWATrfpOat1XGJHj/+5uD14CH2a
JCGISJqXKdknR31ZPM5V7HzLVeMl7oJANhWrlzsofYKGFceGrVPGcG/iK+xMZ8/FAUQOwi6CWtzp
cFYQkgO64gC3ROCCDhzFgbYTMc6Wm6/udOOWFC46xDdGJ5Q08heCyEsayXfjzEFuCVdR8wV+Yikv
9Y4ys28ul8fSorGpW5pup81tYuK97FgJy2a8sTGxTkeBwdrttoVbQkPPX125AWlM13NfSWlL0PBG
orrY+cgAgR3W1e81oNCyxr6CW54v7KJ7DAy02aUypezwjJIziFShVshyVU7TuTZpYZu5AHuzAqvU
7AQmzzepT6kwlp3hdUopq4IBAbqeYLyhLNQimFkhQ2TMUCgdTzLPCUSu6Dkih6VRcCYJFe70p6AB
VeiXOjEFBHtRV02bk5dQxvjzFFJJCpKbIdnvzjxcRR9AksS/Fl4zmbNnytKJXjp3v6lnj/ds29+W
FJ75dYe2fgR13ui2bUpg8lf+nZdXJOaLeSeD5WoAv+iD2fMydkq2vk3/rv/yVpuTl2z9SPVTFjbz
y5TjHUHIaurxc2KKovJzhItnimMyq1HzmwdRTAgJs8XG9emS53L0FYj5IuYIaKoyoGyAW7mwlQoC
awrDEcAJWikIcSNDgaE0Fo+dDJMCWOqOvGDel4GNkqZp3LiFgNaYPYL8+Ddco7QtzVQnbimcLzyh
DSdOafePHHRloaud7GIhMf8gOUleHg5CfFlqqsmUhlt5Tc/gPXzNNZALrNS7TscNiam69Z00SuoB
nh7LZBTTcd7VFzH6tIebEHbfjWD03uppNiBWwry21nhmQBVj3Suhd+lIXugk2kOJFfsF+MHYuXgy
QlbS3aXV0KC4g327hB9cHsCsQHSyzhK9rBKcFZLyBIYO5pPfRDQaCzK3qBRNHTEtrM/9Z9lTM1mz
bvNmvOQ2zFDVZ+k/GzlVQkCbAn5zy86iVL5D5NSrT+Aw9+0Tjw543p8BU8DaCalhoPARZpnSFQjG
HbF0F5tpxvuPeO1P6GoIZIbXfUakVKz+5hzT0BRq1HgmDtwRh/0WDQ7b80Uh4iC33JIlviNr6T/U
8QHuS97kK51xBrV1uLDmHHtTOEKwTYVdqJDKq0Pweg9o58T3TDHAjy2KeOZTF38IMsZQdlOkYj8d
3Mb2zTbhXcBKXMucKbgTH5HbcUwdoLrmD1llsMQ+rA0SAIHzhV3X+wvQ0F8/Q3zRGDtDZ9530EqP
vxDbXU0cBa6TDv3WGIHbWuqdXwYQevJVie2SUTBz7+rbBi9XL+75AfRgldUtOUCsN9f9ryL5HG+g
qA74bwtBTmCh5HhxinqwoUHVdyvn4+3dd2AUsTt7sKr6lJJmpFzQFczu2KzlSlVWElQ7V+u1eCIe
wb+Jvv72qQEq2ZIdZOsyzaB2UtlGqSmtrHm4asI6GoHG7cL5eBhMowTMTPz5JlUo7ymTXZynYFwG
29zDpIKL9tQFB5uQS2uDF3qhLP8nKFgNYS3fG/GRHcJKkVDkasAej9lqa9uvR2ONQ14cZ6EDShST
1lIhPjLJ3JdSz/ofsQ88jD5kwq/vW0I2CBqjz5ZkrDtK1amwGZNGk1tVFxTojXH8Aj/c2QiAuCAh
vlUeCa26tQHl5WWuvp3qr1kCHGTNrGuErQbabFqjzvTRSx4KMDKmlBykWSFTcTQOgzgsEpZqJg6G
7Jf1j8802QZL1wQ4dO8lkYO26/kGsiUQS+PZLyXWCCwltwcNbxmjCgUiNws3LTPKbFyh2+SrBObF
DKrIZZR1dN9eLcMEUyP9bcpRb5F4L04fgAOYm0Gf583yACP7T4doBeMsw9o4VDiRLEUGHUYlyzUB
zySJwjq6eYCkk+OI8lwS9rlSBeLV6DmlDmWQctFqO1DWp4mpFXacMA/S0M0yrVMR3lEKxIUsKE9G
MqSn9fv4HJ+uEn5opA3hwtYDpq73VcTwv54sf+3TP51z/B7n5C4w3mj0LuGBHr1jx0aBc7UqwAwm
Ete5nL9ZwVoqZcdvb06K1ru2rIUkT9F8lHMd0430qJWTlqU636gGqdD/cI4wOZNXM7TNsAXBKKGl
1mAatqBCzQO249G9ot1l6gkvEhNJFTXtNdXT8W7etiNm2hPbCald04EprB0JPqJ3anYG9sr+kfBl
lXvygjJxJ5z1www3hc9L4hyBL4UvDxbex1p6LDTaRKYnRK6WZse0H2EgMpa1zKLAHdfFUwYWGY/f
avbR2mgE9eoA7Wmvt0ZnmJn3Qo6qwNg6TgWqteB3ZOTFU2J43CKFINxxfGdfdpNHOeljfSmGF9s8
i+O8ucwp4h8EW8z813nfIVyDcVHAVkiJFfXy7qWOxiKd1dVrKzjwR3erHux2vZBpCRSwqv5+fv7G
rj+KuvP72pvOoyVAVYlxoQ2L558IvYn8lF7MDdSBPm+DdURxccOCHr4D54YgHQLii9XWE9qqDs0c
Z7A/vkCueDAfM6+STdRZHkoEThkXJdVv5eOdChEQbSJhMy2+PhinwnxArqS21U7hOojjfU1dujgz
bF5bEt4xLHnrAS8JSogAXa/D791x3W7zOlzqtNCSMTQubHKfYWK5qR8akeq0Mxl1e37fsxzLnmcy
8w4DXPfEsI4HUb/mCHUj/A2qONVQDVckPwZiNHkNbyGIhq4e+z569pThqsgWaqc+UAvIqIOyUcDA
Vap6AG8lopGx0xq/kOKhD7drr/yS4nQhSlF+OGt9ICD/hAdFvmwu+I1p9FknJjyklj9vVd7Z8L7y
x6i7M31gxrhY5138Kr765Z22QqF+DxEdDKnAPl3BkmzwQhH+2xcdHRWXB8Dp5xG1M74h344KjT1q
CzO96OpPl1cegumY1Rm+9QBE9Blgdw62xpG9qPeZn1RIzSpjeO4hcJl6sB3ms6YS88TLJU3Qm5PL
sSsh0MqlYClurv6fgZKx2QYC2KSzDcpEYmNlIceTEIyEQcGbJJ+CMRp3XzRES9KGP8EMzWg/KP2E
S+wpNmvxZ791nfJHwimLXdB62f84GQtSu3LL4Azh6Qbb3NBVHnkOZYTDmWveWB30RCBSxrSHB5is
I1q6dAoWR/nzWjYTPUiYu+3/mUdy1uSNTWDm6PgBakhd8oCFAfy1MqRmvo8hgPpnGBV7SK3sQ02V
pE7mMHgSC0kLN1U5ZAoOSkpCHvMG98FrhDoyv0GGu1SVBpz9mwDjIasED2axN/NmPm3gPl7X4wm5
dlgZwekV23JKmsOr6+xc8X4d1bxhqO0luJZVM0UrGlGpBykysyKWJHkzhorqRT4vpNuH/q08aMr5
+oKTel2zyLgzrl4y3CzxsANZiM9QlvTPdGsgy/g1C1VutFJoMXJIXUx8yPiDEiUyV8tiWkdOZzq4
96qwGHS6+nRQ3uq/YmTJoBiLcTmrrZrnJdkyC59S3DSfFAJ+WvypykzcWZmmR53YnKOEc0R9bOl6
m/8WzbkQfxwIj77y+t9PEZfi70oVPpTbl6ocyqKWUyL4rYZVnDZIHy5D1GmlEkr+mRQ5c/RPDW9I
yZE3X9kRB/4SHJdDALB0QzBZwEe2iEYSMKbjqkziuRRCkglhctQDT29JqKE8f/aWRHxxCZSt9iP8
Pf0NRbGwWV3pLspJOpm9P0FGI8wDx3Sf/I/TWQyZc0374RTL8gUYF6SzjAbKu19QUzJ4TW6ZfQHR
41HckY0j4qANlu8MQ1HCq9uqV5M147lbJgctFcfy9Mmv48bVy0Gu8jvxsOQJgYEhyAKbqLncgLhZ
SHCK1XpIUjnYDsM6Bg1FhKowg/NQD8OULSqp36iuiG5bTthjE3iABfIh0hbnv1Jo0IO4jhxjNJBv
dbW6AEmYJ9L4wZZO+UMO7I+PBe5Qgl9H0+47xm/RdQ+2w+3aetVgH11uXpQgTkd69jyUBbHlc0Oe
YBhlH/JH6sijY7RN5NngVlsMah4763apNHVCAeWnAmQgKxti2EHmDW2GdIJa4JeSYKVkwR/9LxTz
xKvrtxgLhpxElRNzRfyb5IY5v30PP3cDFy8rPO8s5tkxHs6gdxDZDSmQZKqNkpDDL5oV7Dv96htV
jeOkuQKFoDgrDzJIep/qOtyDJ0kgTSEmG+0GIE5NrfGAAZ1p2GmhVjOGxUmSOoDb8UKuUTybjeYA
fsufYqHrGiwbYI8wGZP+psavMQzAQsHHE16HR4yOoDO0272JzfZwso9l9fbyiieyAUaN2kSNHVHW
/Btblt37BwdMhpNjr/3COi0DpZNhWS0ti4ChId1D9cWUQE1GofNRzU75SJGP54icrnol4RiurqUU
+FIdzUE/moZ9xD2bfW/YedZm0X3LVb0MEG6VaFn62gTEosQrvheOXWGyXCeD3XDIqCJKmb4IknjV
smCeoGLZnc1/NfWK10U5LAE0rlwyu3+gcSaJU5++ZdDq2hmkO7Ba7qTWuhBmF0D6AkwZ/Cndog5S
q0a5PRseZ/MG7uluMjQDDCkp4jTrlRgr2mh1Fw7aTTu+YQooRMUOgWViYLYtvW4X8qrfA7tK7YNH
GwDUAgQHWafAtA4ywSisTYN3ynw+27FcTEYbNShfFWa+P06ldgyjPSWKTenjewlox65bqjExJfN6
d5SRRp/rwsRf9kbJWCTQB+hMGg6yrHLL+PFfH/GYv4re87JJaEbonWG7R/HUEFHq/HZLTBrJ4wzb
quX2fHxMR02dar3UMqY1T3ssh2JlzqIEiJ4auJwyud3mx9fzKgcFp71H7K99b/lNtlGNgfCuDmgo
0sd4nXSpKHxK0sVa8SbYe4jzWyxWUavZ99Fqxwegqjv/iHGvGuoAF9mPE8+s4z12C9ZWRzGCoCIH
O1XqG60nH3Vcib0wpLk1VWzn95wTMRaqsq+6YSNj2uyBEGDjvPr0BkGSyKF75DizvWHBLrM1TKKP
uR8WBx1WV8U3X5tbFK4WFQhJhZFRbFmHxbPMzFEGuBtVAgaRnObz+DL+4TYwYtkjyoI++D6+Md20
7L2AkmTujiRrWV+X9ARDc3nzSdaq/Cdh2oh8O+1dwSzdoQRzqaUr9fTVsjQNTpFUBl/97vtJ/9R9
44IqwV0fW150KtW6tRpHRDtAySK2qWTU6DIqeBsL7f6l8qzBKQZ0vMtxi2TnUtKzsrR3d3xDhLVW
8XFQWJq397yf0jALdgAKRypT+WeOXQIyBfi0QLloRpMtpaMbsJHO3B7w8KpkCqmcZ8yG8/EsnWOI
MezlZDkj80MerGqooWpjAfpxuxAp+75L0lxUcx8ewVqnqwaqtV1iZrXxJuYhNEfw2DI8KxnBWnFp
ExCA78vRWydB2uZadpUT7nzEk5Ax1Avd7vBxKqdTvm/cX7FLqBKojR1zrgNpQcw+U1iRUUFR9eLT
szggbF8c+QgNY11zdA2RSpN4sCWeYzKUnooqzJXMfk53zCuAHeFM+rzte022BvDG7tDP87nCEqaP
zemLsMNFmaieyWZzOfC9g6ZzqJI8Es7CDP/QceBsjXH0ZtGE2r8W2GwlXwVc5F+Rk7J70gEkGiH7
XDK6RTjH3aav1eUq55+CkA/VVVD6sSIhuf0DO+plTRojZkzUY9+w0lw8FYg2zwgKrmDbsIkkRPhg
CYVbzc3UyE2u5C7BPZnj5Z0d3wB0wvfWCzhvX+eu69fm00/31SLtEEyupz3BUzDpuymEzZvcZKyY
ZoW//5Dbh7zrsC4gjZcZN9ppEfmsMSZ9A7u0/l7UrOxVnkbz1L8OkXiuH2pUoeJhOrKfhyDs1mB6
Z122FtuEN9wfeUxaxnFuO6SphCowMz6vKlMeI2gS5pU4I1sG1LTWdCD5sz2yk6ZJzpO7fMuXA89l
Hhc2v0fOzgsYD2GaomTOLaaPiUtD0WVkqbIgn19VuYt59kfsaTiDY4QSH3qX448lno5V1iugaAIN
/PtATmx0OH45g7mK6pbDk0WLjtPNDe6lTDSmf+qQJFOdH3X4xBgGf1fUzt/vJc0ea0yrQzAXCJLr
Gs0qORcErkiNKVVszgNEhAcMpvAc9uwNDrwXwAUfutiqU8q7kO/zTp/gC4DoTdlTnugJFgA97WLA
9mJjtMG/TDpy2GTUYQEq8GL3AvaznFrNEiJouXnnN0/N145NmQ69SKH2WERaJLbRVIGXLxYJYTvW
mUlMx19bD1M2BNzaiOzYMBrUCJd+gJLv8df4yrM0VCeJeiB2IyoZJUB1yBisW5b5tPZng9Do1Q+P
cvVsRIxEa5Jg3B3Rvx1YdqV5n7dhMbV9VWvhMCDVGyVnQOxqBRCR61sA7Rb5SWOFi2laVf89RMrg
xCEub9UNmQTx+xqbSuH00wmWEqt5oJj4rsueST36X2qDkt+MVDaC05L8Y4UVZjrY5FApPIFRxiOx
RoVbc9McYDIdXOlRd1Y3tftFDPQVjRqfkPVmcgfG5Tnqhl1ksLKVlaDQPjc7ZG/YBYhtnxFFtfYs
7dF1RMVAb3uSX71N1uPfvrzZBqh9XDgUHKZYUEa9qpg0SG+UDStaSNSxQQKFMGAo73drbzjVAirm
rrA8v5MHJQJFgHcThyfVwy9UtxoeW8XmF2xi3qW6XrgYIETIJOcWcrPfPWLl+ODLmvugDc+azqh2
tkasH3MIljdG/k16zodi7uOaU8Y6jY7fW82X9vgoIYC0UMN9cWra5UE4bB5IcCGvovOMLA92o3se
MSY0VT3gm/mraREd0D0TcGqBNNOWdpk8js2LwOtywL2G37YdD474ukPxSlqOcIw3PG6dKnaA7bPl
KWrr8l5ZLzhSJe2BwvB7SF7aX6gNcThlaoDouy1OROP1cyHpgPdZrFhTHrZQHevpiJ5LgMDU7C32
0Iw71Cds7S/KNjYJc0reYjIZZ872h+fFc5znDzR5bdF2l2ulah0xs1vE/7nhUw1HpzqcPa+Bmvuy
oRUM48rQImLSE39DjexZsee2fZtdKKNmwKj1j6eiantZhLEW1or6QYDngJUkdavTWCk8++jeSa3h
6Xth99fh7D6h1HGXthP1qcrV0D+zBeeZTg2mJnAWJkkXjh2My5pMBtixQCJ5SZUsbe0OV6e1/WQc
bV45sS4kQ3QrY8hAcLFbEdANOgnLlwMus0xyu051b4/fuYuiw0+dKyxol+Kh1Kabzpu5xdHdkrMf
KbOX8fQWFNldtQUI9MOBya5nN39LcYztPvW5lArxWJmmaCkkOi+ltCgXB90ZxtukXzrO0jBjuuII
omRpRJ4yi3I8K/9nEVX644lvUIHfLifj10JV8ECHGNSqEKcIp7eycfp4Sd+v4FYWxRmHcLMWvnSP
5Q5VKws7RAM1wpmoI+VXR120hwlVYSmMMma/G0YitHGBR0w0IG98mMDdvyQtfPQnOIkKK6lrDiJQ
sDtUP8iMSbE7VhMD75OR3l/7ScXWgFJhEEQUzfhCxOmbMRBqRH8k5cNBIBHqsmr6V+SjUJ1jYRWF
YQxd6A2Xa1kdliTeTt7KXljRXnwzrzVHMrkK+xw7Ju3Eod6bN776mCvAzTBO758Rk6jz7qmN6vt2
u6QBrD6DL9VSmdBiBX1RzutUffHnxT1h0kIMGaAxMR8FPVE8TgxS5gcbrbzXiTLNLKztcWOTaVkz
Lg0ustb4Y5snYy0g6WNV1hDV59zzJXOlw1W5hwT2FWDGAu9m91wFY68E9rR8wKCxN6t6WLBYpS1T
SOAkTmuyIqbeU8DI8SYM1O3ScDaLcXOG8r48anNRG8M9WfRqUjTJ/fqgDMdTxGmGHV71pbacu3wh
4CeCHBfyahw1xJmk7bTIwoQSqo8EH4WLnczIC7VEaLy8Gx/EUeZpxhwb6etjAJxxJvIcPsqNdLly
Tqj03p6UTIkKlwmxcwm5cWZ9WzUfyroyjfXmlFNYjneGOBgKrPW8Iq/58a9DuU4YDu6tOWo+4/sB
do1ue5ciD3UaxROltrx1dFFceyP4UHdLpAArm5gvceLihTvgyl1MFtgVl+irmwyD4NgNvpPtPDsP
Fy9K73BSSm7ELbZ4aRBizTqu+brD17Dp0SdN7neeIAF2ybiMMm4ywQnI+1rHJ0U5RVetFwbMLyDi
KQ10USmTeTJG3Ez+KyasxU0UTfHezPxcM2zFO/qYuUU33aAOPZT6VgH/BTSUueNiyek8ZnOJfGA3
xL7hpiH6QiJPIzbW5pNp5ZeDjDItzlKP7m3M73ANWX2fbBT9+xeDMJM5+zrRgOmyEpT3hTxPllcY
zfVB+a4Wc0vNIfcAafyqvz2P07UqWH6miKoM0HAIexPdFiBLAa1B2ZbvrbEsk+yMZd0Q+WO9Z3Lw
IU8jVthZ1wnL0oH1tJ7RSI7+xwmiXVpIKdDcORJ7x1Lic60U/+N2Sz2Ix1wNE5XSAsbM/HmvcPrV
K1nTjPK0AUCYua8LliuqL2wZZKlR2bqy37DLIDXBai9AlfdUizQ7n7pfIu0Ki2/E7VRFtLoyxGcE
iHSEtFAZdDZSkmv+CE5IqPZpjLvOHWrJHO8lVzLmgct50wYFvxMU3i5FlwMdLOcvhr/zuD21sYzF
ruAjYWhRXGED1cxNANAkEbL8tEeIRR+6ZfoQePOPctI/RFIEY04r93j93xtlYmtI91vSTqQmHKlh
c0WQQem1cpIbiYnox3MXaN/S0fcJUTK3cYvKvB47qN3fF5mDeHf2fDJYQ+YjNrRTd0WKiznVTnIl
LLXrDH79aQcg5nTpvc5LlYgiYvKGAzkaVBa9Kp0CVFexrer43XzjFRres1lZvzSiOoGRUKYFRHHy
Nht9+O+gykVlMw8JxLFXM3YnD7jybDCttFRyz1w78BAC5FUKuLmcM8RbOSjqQ5Z8LTwtICRxoJ1F
3x0xMkrJvlFSfIvJvOMzEktJsS+X760HBg0lveql4atqLOGOoRI19X1f+lVZM3n2WYDIh9DC9JgQ
8VB678tQW9eNTMDJBk9R+/vpeMmsNTzATqsqtApoGEUop9qDdWmccJK5uOHPUx5fcWlIhDegZPEA
4DQCay4nH8DWmuRsLsYToua8QLBJNRCBrJOLPmRWqz0gNx/67z9EV84kg3GXx/wntNnJDH+d62k3
+cbde8wqOlXcOE+UKR/5E6vfP3EX3WJFwt55OBS7pxNWONd1OP2tUzg0RKyUWdTjHyL8xV2+NKzi
nKZYPhdMpnoCOYZQj2mwTQZgKL9C1oVmROqbFMnLNhw+jVkduh3TmtLoE+A91zyo46grrYFvkDKt
OqtC/k7BHdULAfQ6b4nRdEM/iCp3ogd86FvuBsNKKQr9rjx58FtwD2J+LfRnX3/cvOosKUqSueow
w5E+ME1jrU7wdsu7JOVrICtSYmynAtaOpVrd6mgIDsIAPMkmHDxqmxeD5TosjhqzaJ/CVg3rVosN
ElhAsl08PKrUi4QuUdOTbXN0wyFU/TkN1Rw3yTvpKd6KWNyvfkIhEpcbFGDx8kim06E8vK4MP4Yv
fRK/Hy7A5mT4BNNBTFHM/m0MVmcngFegFt3L0ANZIR8NgFDqhu0NKE3QsMCD5jxXyiZ4mKSCpfiG
pVO5uhS6ajhPEfc0NWG5I9gXU2IqSew7BOkHlcEW14TEgmMeYqncg0XWUOPt/JdlxXKZuTGwvV6d
YO4OrN+Bit22R8VRLxOwnum5VGWUIQ0rrqHiA0yw7JyCNsRQENrmbJlev4ynoXBFmSp2bEkPv5JJ
fxSKfkscqPGaK2RDcIZl3qciwtLNozryP0wqq9oYooJrkj1xSp6vSKfLuPJmGh4+oEMSndCGLlwX
i/wbX4k0IWdChSGs2u9Efqa8GKcaWctdf8PZZxZJPykbNj8CNVsUBj2EiEMJAJ33+nSD6LEWxSpb
E9AAcs+QVNqfeOuYvC6OuKLAVSIM11AyG7aYq9raVhjq0HrfrmuEr+u5oT1QRTZlYOEohZ+BkPhd
tW/9jOnnqcMHco41RF6bddPprKyYmaTwv3cfWeHoxe2MwYRnE9ViyuPw1hdZYk2mphZaEcqYsMIw
HpJqyF/+oX02VMcdoFGOmeHFopR0dO8foYj8f1iRUmmTfkiPzBOZ/S7L4leWBvfcVYsHh3zs/gxy
29H/mxjpIe0o4SciVacQfxbmm68thpwaKMhiwNRZcGdtsuYQzFlRQqwsEYn/KShlj91kLa+giTW3
PXH8hM9Cy3h/4+fB0byt0g5yWRaoqKp7fsWZI0mRBUNz+hBoUBni2c7e/awexnGBnHAKkjJp+Jex
J76d9v8wip8SbfdIabyt4ZvnfcsLR9j0SsdwmiLXZZAh/zbUvaxFXtkR7hF7+iDFrOQjVDnncVLN
i/jN23ndLrpc73IQwSCgRl8pT5CrfpR8BNt7cYcOnaVa5oeB93P53MCoBOVxsxu/fmwlKWeC4Jt2
bXfl6Jrz/A8HfLar1+q9u588sfGBt2uK+VzFrFHc9vOIHh/Wh8nAhaw0ihPeLkp7cJjaAzAAC4tT
UT/GKd1Xf4sFqjl/X9W19tZhXdv6hh4ET4guaAowa+6gcuCuLHRSmZ87TmXmBPTfkcBvqTpRlyWC
kcoD9BtEumjBPm3Fm8+o80AolA7z75Kmfpgo7zAZcubGtledrPbuVaLHCfoGWvOTF74F5zYNMHJD
xZRIUStnqsXgbcpLlAi6StyfBqhE/F/EgUiev7DTm3sY0Au6wA4HUojjZMq1h+J5XyH3eJujX/ms
ROT+HckxJpglixayRl3OJLD85Z3iOsXep35iqQ3aBKb+ATscQSU3zThe7da2CDXnDYG0ypx6Ityu
9qVxmA+t/rHjznXzi8a4dVKY/8VamGRvoVrMYA0axGoaNwApDsJEye+DHur2kZJpoDiZOv8Kg4/x
E2DVKkRnOAka0FP952rtWOeMOU50pd3gukmqDr/0mqwAMXugEo5pgxucPR7auC9fmws5I1ywQyji
Wwgs7uSH3ubrV/tJD/NqSWnJOCat1bsgLIpDCkBkEYn7gr0T7/o2z+dneOc47+xK3KtEOZnMkLUF
+WHUR3pJfbfQgGOWFLNZcS2tbFxDVyntzg+5GUaT4Jj5BfUS9RlVQmjM4AQkUqDiQMlWYGcA6oLF
4v1yJrnMEIxwUho2iBsVXO/on6wskbS9IIDUBxkJ/6cWQ/JYM0NYHE5ImcBjlfB/EhgAhozPdE/d
knvouWqix8h8qf1vV0Q+G7MI3aYJqy+GP2tmIfWyYATQDn4V+Jz7Cag4KrKJT5BL4M4wR/8f034j
wA2r5qVdsi7gbL1OE02SsShLpG7aOPgzK4toF3Fz9Z3eRKTrY2pQkX6t4lrZYNkxR7YUgOl5eh9J
auUDe3O5fbUzZ/ZL4gdyQJ2u/7xLSf8U0zCda9EO8IOiqSKPfBnQd1gzautqtrGyB9gDnAk+sZeQ
P9lA00kUTzqSNaHxcHccZhF9djLFRdX5Oqt5haG/n99yMCgK/NHuAscZZb+aaeC7anZWg7RXJUeg
N1vf9CA79JDHiCXp5yNvj7QiSi+846qu+cWSwEp/+uSBsZqAKF9mFx1eC6B/CdoMb1YS+pJDJqip
4et5b2AiQ2llB0OqWHk/upAJKHsVIBuSEHCScvt0UwBWBj4KPE11d5yjab5JL461JXcm66EQx9F6
h+8ZNxw69/LDLY1N5sJ0DOJ1G0Li9q375z61Z/kY4hC9ZVPjdKXuH5dhlKh2S9VnYPU9e1rO6qh/
hyHFOoydiDeCJAMYZSdtJNz9nt8c3WHyhWAHcxZnwO3Eqr34O2PR/Fdcg/e8AApFgc4EvmgcXJjQ
h+AfH6+XE+ZdDOqxK8G6EcSKRx0IwQVvqbo6+OXR9sI9STUdOpqszUNpp/vSKyS8Ah7o7REBjst8
fFZGUt4iSw5hFZg/yf6lqb6kzLaq4fQ1WkzN9L+gUehq3IdGM0PyyRaZjRybIOPkZ2K6q2rgogdG
CT5VM2HC+2V7kJEOA5i1iKx6vwwB5aMuGQNrApaPqwtPuwfmGsXE+hO2n8p6tEnL4c9gBc/oGHEM
6z0X0ruW9dnuOG7K8/b0ULVbZ8i15w0x7fJn9vossQ+FEuBkoWJQo96QfJdp7Hu3iBmWAl9o8JUx
8+bj9jmYBFJtHJ2drBOH1zSg/sX4ofrFGy+1Orx2Faire/zRdzZd+N9DktY6cx+z5IjvcoIY2Nkc
Rys6ZHwepoz/C8DA5ldgTEzMHTYsJgJ4zAzMUkJY/SOmhFvSZ0Q50Mb+JG2iQAJbGkuqIheKv1Zk
LduXyer5aALeHkpssiiBBLLpgpg47cpVjTYGYspWHKOkUtWuwnvH0rNJd3ZDRdkDZpsBBfvLDr7e
ciLJo9nJdC8J831rjvDKmEwaQUxbi4pL/reL+iHV1glNO+LvoA0Nrd3aDNFeomzDIdgBV9vVqusM
wS7nPTZ/fmKcr989ZiaWl4O2iGPRvt1qw/HKpD0yK/h8tF+jqarm13LWxUXcq2GbAKvq47RN9nWg
jyEmX70oQTogRb1ynwpaEvPSGPFSRGiopxKheSSszNO+rmA4Z4T9Siloq/CNl6AEa9tV3cBAaBil
jGyDod+3pJvfHATSmKcVOWcTTt1zS0tc7/Wljc6zwwzTMGUYBFdJ79rl8rcjCkU7FKVXej+8E+pv
xJGMW35Bvc9EFiMZ+j/kiRo7og1HmmbgGbU+H2PfxXtnbEQrXzrdgRsWF9cHbTWyjteaZCwAiJR2
ofHLawqEHhVEWQ0GbAj+hGj+h0q+BIVIf2RfpskRCGPntLdDglS19jjGjJpFP9k0c6JRdTXhPcQ7
mM/lKd4Yk2FFLnh5o0zfq5ydn8AvPBNXvcyQ31JFfBZiD5msjsvIMleHs39YibT4RjCN0KyoqBli
2MXX7jQIQUdgp2XhTSo8tePmhcqSQTbI9zwJr/NBH/TkrEWHpiB6taOjDbBFxKkbpXzH+/xTBVDp
2rUNIu4WhV9FoXPD+7Dl7oP64QIej9FqFgmMJlpY0QFH1aKk8ToKmN/dTRV78zW21xxXXeTT+gMe
Knz2TElsNf0dvLUWq2I/q2xvCQVq+AuJYW7KVSU4Qy7Ac+Lv/PCaqx1kXKq952Sm3a5Nk9WEJe0r
A8c8s+XEzprGTnOYuyDTImOOr7TCEz76+o0ITSjN6LuMIPPJWiCpoatW262ewNE0tYx0bFgwKvO6
XqhM8LML1VhytwHrVPlOBA7YeZIG1LMC029zzYiOxL+ek8uCqyVOtWbO8lScefVUJjf9CDNSAdID
oyCEZI+HBbo7yfjni2gXesLhn47rmDfIrRte+4YF7WCFDgEWNNO0GANxSfoJuDtcVc37CirScN2l
EEyqpARriGqp+Fi5T7ref1GKC45ne6s/uuwpRVTLjqQdkKIWlri1Mibu2cUGUWXf68FKk+WdGxpt
yMs9KZFe4mU1fpq6w50CWRqhpcQgJNPwh5x4kHjVCWnnLBJE6t5GcrhTABIkrj3SXmNKB0tkDJlC
rTBJy79RN8tWlw0vbeyo4iwMxiB4iEMZy9QAFDYl/f/zpJjHgZYQqI43+tKJ+Ytn1R48bK4iE+Cl
ksTZdWNmnhd5s85MEYqYsWogPLHbkHRPyM03+J0QaIDmHpV7yaGupKPtwfBv1zJMNsyrNH6dOljD
BBP5EPqOiqfNEkDTtT1Zp36o6fCn440u+3MXiTtdKfyx5MKIorwVUHWmXsssG4XytpVp3kDIqWUA
1/Uwvu8Gb/8yM5SGfLnE34G/OaPHVOZrxmuGkhIpzryN22tLJFRQ2AH31pdsBrjRAjJXg/dMPrXY
K6pTxbhOTJ95cDF242n7FKklYhpVPnGyIuFxCtfJ/p9R34s2pF7ZjMiKfHyQKcCtfTqkaJGV2Hla
LuYkR+gDOHFn99gvAC+Wa7EbMkQKm0bCTBXhynoNNhpOY1pyr/YOwNqS2mdC7QbytGSOaK+TXLVh
M21scKY2lXlPQJa9IXhtUYM/pZpI4F7QrbJgj4KMVGf/YVsewmmhKKGw+Rprs45JIyNu2qCs1ju2
1tNc354gwBoaTTlMWtG2PUtXitZnJepFjf6IBkRFkS7pKrkoBYGfoXwqpMKd647g6axdmKQA9rhw
PPFbx9U9guwjmEqXxRkJ6fzsi90fdU3vVnnaihPHUuzYIBssFm5vABkE2RbM/gQaZUgJ/f0pA4JH
A4Ph+cUwIRUVU+mMqN3TkcvGTEtDwpqFoO25wzjKCOoaP+e3A3xdkXHkJpzgE10B4ccclOegKQTn
syyC3AUPuLIldHVn7IoIu6dXA9CaL/fKhNI7PBpjau5wOBF4s326iQtEJta2/4lrUGTbsmdImBRd
hpjyjCWykKqXaT0I3Eardn6oIMLOysZAlqWFTS/RzeO0l1T+9SG05ifN1+njPvRCQmRQcit220eu
uE9Meb/iooBJu5cfJHb26SFyjQBeEvNL52ajdPB2n0M8YvL39jr5DsHVzyEDKgT9xRgV/h1OccT5
ka83alAF/mBD7+q4YZvmqlD671pBbH5zXo1bsv+whpGqhVL0Nzt6roPNtAdu/yG/tqQ5IPJLrt9Z
t8pWVY6HzCQzUFk5cDbtcgD7gdgLyf1X5kLvmUcW1GfdkWwHsi5cSZAdecfReuAp8NvQ7jifzueg
n/BtEFKY3Vo5SaAOGwVUQ5LrfYzdtcAe19m50NhNh7YLM0v7ACRlJkT/B9B5bnEQMhAiR6rrNCOH
w/9cr/d8Fq39K6yht9TL8ACVFP5HZYDxAaupqxvl4vdfVGWyOeQaTdQvQ3KGC4UmiMDCI5PXDAJc
cuVMz+bmWeyViXQ1LDSXq6Pbv9kNuM4Q8IbbB85ExYV4kvsHsiB/+LivlHjAV/La/Otzaqvotzva
7Nv/RFX+V0+mSTkb2VuSoc6ncIJINK9Xy9jjD1db2a9B6kLWFeAqgGcFnUXWwvQgDSVgMK4Qap00
DjqsSlmjoBzbHI25CV5dLqzcm5CiLZF4DF9tN7KWZD4rd19AvxqvlxGltdp9FzlB34twNGEQRUeo
xyTr0wrCsvb4ydRK4oIMNVwmoHCiIoJKw5CNCyS2phqnrZ37/vFqZNGtxxfnrbRh9Wqs2W1q9ISS
DwM8QPDmAnbck8cHH8QS8ixWFZKsh53ZCoMwnxJiXRSdCAWJoVe+ZOGZHiKuJiJ5STJkho2TN2vL
c4f8teutit2r/lS5WPzUIE6un9bYwKAlSM6J4Ro/gdzk7Dg0W2IJDvz89iyu8aUiBbQwHudasqbc
cGwFw30MXkpUO/GwdvXwANNSM613JDZQjT5Xk1/hX8SoKjWg9o5jPyiixQ0gbAY3BcRd+SqWzKIu
XTflakxB0cjbZRJ+ht9ZGqKnRj7IIk3AGJTG432AdGXqWCgXR31tIljip0xOrSQuJOfARuviLMfg
DdWmICgVzhZ936dqc0gb3bHTcQeNJYTcH8JFwljEYUFiG3WkGvRYcUSN8kd2Ch0MTyU9Eckp4jwW
1ocA4TvKzyOJJlTksyZZiFhyhKpL2wLq9kYBK10uTm+6s1iH7V7MhhXJXHHnNz7Q/DXrR7dTmGL3
JnFSGHgITdeb8Q44J427pgzn62LdXOwo7TpehUd9c6Cm22eDbOFXoSD5kF87yArF2ScYQRFzwIAS
b8gYuT+Vj4e8iLIGA05eZzfcinLe7XhTOQBnJMLaB6edXT2bw7iP1RtvHWuUvLOWql95jYQmbJmc
1P4V4Tt2ZaWdt9zGPOnW2G8X193Yl4gcoWUAi7HopW7kUbF+zf2UonX9PwGYP+Sjne6FCkcddYG1
v6cRJuW5NVvrwDoT/cI/OcbuPWUkDj6v8qIKLk6Sq08rJaB0JIC5EkhMVm+eCq/ErFcPrUdxvkTZ
NKiV4x6rcYwy1Z/ukhi0xP/ZTIeKVdttn0FmIzPlHsZAUQjHiD9irf6b0TxA1piDNoKq0O3KxkxL
ue9FfpislEz4/slNaluqhzBArfU+kWYppU9xXIzgD0NkQk+ttkReb/XVUPZmPun3GcPzTSX4kJVJ
r2OEOQt7DbN8BCuPEjaJ1BZ47eobTEgvh7AdOojJyUPeOmCPfay88B57nLFSAZV0uMIAsBY1v6yN
ZBTJxJAyP2m38VcfXc6XK+Qxg9JtMZGRJCQoKGbUiLChYIwT94B8F+LUKXr7OJcMiAUR3odfYHOg
eBJkmsU7/lFuve6MIb/qNF8lVagpBj49NpOy9UwUCmdU5dwuAPQOhLvAkltuYq/oEY91v1M/8v79
aYLJMHvU1lCuNRanpAfMJA2Y7XRIWE24qNuDkOJs1mFp/5CAhlUhGC3mK4fmSI8dW7FZe4CqzvPi
P9I1MDoBwlRMT5L8Cya2EBZRh27Efoim5JpPBbX3vac8pPXrF0z5L78BDJcLEiRsyvU5GCl1ZeXU
+10F8PgeIFC60c5WAjAufRbn91GlvP5xjBZtKFv9osPdDloIzzRB4mtkw6iJGhyk6XK3uV8StJI6
t8SeFEa2m270Nvkt0g4cRfD/fiBeRDO0JAWe6RJ5H92EIGlJTlgX6r7R0dgUIWRAMmB5SifJtMH1
yqbC1oMFteuZ0bQoY3XRSvnQwmMX6qliU4aTDSq8K9ILGvYy2kmrio61wPqqsdPiv3KYGXEtZmtl
MwypxG6L2RudrktDf6MdE5pzAnMbr+3e/Tv9AZdtz+TFamYaVSlIpWpCY+JgBbVZXTFPrOExjAwC
JP0ZEr0UEc7KjKsY5XHpfxx17j9uPjPzZlUQqbPH3NRMBGT2wS69RMNsJnRfsD+LgTtRwhKDS7Vb
IvUA/LeS86mGoXmcUqTKQlTqDMiTKEPtu218ydC1bvfLYvp+090Q29CfnrRLAm4RxESIwxKSWXqS
BJ7gAdQ6a9otIt5o80YIA00vOWEVSksHVu4XahPfatZOG5kRSJS73mWrmSL20/9GtUcz+o/x1sjg
AyJD9c7784dz3xaAlwwYgV+O1xTrwDlMmmY46+kWmI9w768xPJQCpj/DiVEjy+3rtx8jy4FOvMIk
FerBhYMeI6N1CgIjWt+cBkAM9LDZfpI5evBNHeVLa3tHzWFDuzV2Yx5j1jVxOZ9X0+Ha7v8pI6YZ
CWT7xGqUb+O7Y3H0cuIhLlTmsBxWjzpXCrl545AAEmmnbasaoyCNbXye3eOSfGcGOR0H3rJ9f0MS
p3Aqt8N5hrCNjfbW4556ldQ1pNaH2vgwQr+9uDDkt2yUefXxalc5MjamtXmI/RCdnep9IWlJzNaU
G8luLcE8npJaqZEq6uHc2kqZuLl4W+thpER7YI79gka/tzTyEbnpHBLgQkgvuG5l4q6sY2U97tNk
xKPEjFR7RJI3Fs75VO7L80/5x3BI2qgpiB/Hv/VHpdCFsUv/so7s4z3OLEifQxk005M3y/e7FWxX
UkjJy6+lJc0vjzU7X664TpAEyibetqVFAWb4BoTJ/lPjUdfeR/NN6IL0nu8z9yq41ucgyDKEk7J1
vdMWr6GlolfE81O5Dfg+3yGPKt0vdazCwKwVI5oMaPxftTV5yWF8Qgo80KbClXrTgJehSDl5zQId
ogKJY58lX/GK4qiaYb8/2tlxeuUTnpCeN7mIDOQMmOAfSjjJFOlnLs7yqs0PuvQmMaDHffSaQyih
uKxnKMvNGVLMMwx+0D+H2Ih5T5q+Tm/5VzJj/YCUF9nMC4X1T8eTuSAL1FJluopjLKxHm/aNZEyT
N49/kYh0N0qO8nfx3sl7pbdnoq5zt6e6dHridJ31YtvGzYwX1fqzbAhvK7izTCA8EVLPkyQr73rD
t4YUval+UgIuVlP8HlxsO7XyUJx1Br8TMb99ZJuuiFjvhkEwbXCu27xZX2qbrZPFq3gicTjwJo+f
tmQK/K/bENvscQDPTf4l7OPpTizg/S8IblfFbcL2am/nV1tu2OYziUnafpkaRgrvhkL9EbsUqHd3
HnwbC8PtB0SgcD1OVyJrVbtLGOvV5vsqtHg9J8vT6sG/LftpR7cYUUn78mxMk2QsYNSjiI6amLxP
a9UBd0DzX5kyBaMSbd3Plow9X7KhNfiTTLoxKHCpZ7sBu0+molTeQHWXlbBcxoGEfddK+2HTdjv/
2PixQt5wQjw1gTs1r4hXobuesuAnqyQmg1nKY12JEu/1ruNTvd2mOBQyraItyTx0BNMltf9/NkHd
1NL3d8K9mwfPLGLPuswdEFklkUBP1wuBOkxwy5NNbSX9MuyvEqQ+P3rpFpKHkhx9rJZJi65ZkZSn
PJYqP41VhlIM20gHbUSrlf8TWsf6fPbb3c6s24TLWKmXS2iKRurs4sHvOf2nxVThkl7JxkhE5WFO
+0wJFxqRRMabf4f9EdEChNxTyVgSWYEPrJCtHg0gPutwFmB7PyeEt2pyYGDhc1gvqNBwR7SW3SH0
mQMOP9iX1kp/jvZ27yxFOq0I8ZCpvX0fiwwOg1aJB3EMIEnpDUwQ4o7dJry1C3/etgAiGHHnmQWL
3pPhizNMOvJbrF9ut6vorF8ZyzcDUxvy4qvcSfmZIhX6hlzdYFOMORFtQRyMcGYd5QNwFHv6vhCv
9RabJDcH79DL9m7fvJCImLYy+xeu0g3iPDMGxnF+fraZjfKxYkftFuiMcAp5Wv6i/+oRnXI0w+RC
Av8mDx9HXly9ZlAmgJnb91FBBDR1B/BmyumrTa6DzQA4QP0QpWIGwcHvITgPf8v5+qUMN7oG6RPb
HXQi9FkGoAZyvXkNBUQvc/3wRIXYX6L6LOmezxOq/Si/CiX8xVbbqYQqnjFLDyRdJZCdj4Rp2Rn/
sjH5ymnWmjimV6vMQcWB7eYP1qZXPddi/Y+h4HwEwW8fFjCgWGPJ54Jzz/6qft9At9fRqN7ZWv+z
k8ZqLH1WbqJwMDndS0T3vjbp261jQZrZOlMfWKYRzvi2GpHV1vzrMkLv82eauqfDZ+8nFGMMDaCb
IdqqRDjgvyNbYQ/nOUU4j6DdSxxTIeg0yq5Ut6mWo07/S7e3b0gtZXKr8H+LcQiHs6WkcNk1iKlw
dbv+ov7C5KjqgyRX9UIWUykfS2CuRT0LJyFlaRShT/iyBs2j9a61UHmaPGMwuEOBmvMe8jH2cbIl
+pcD8Cq84hrQJtNHjyAxvHZbYzAN4QxS6j1TDS6Tk24yoctrlvispC7tG9Pjttc5ZZvJh3P8N8bp
nqmIouCWn3pjsLNioaL5OKxZZODeHuQWzomX6j7BC9Nehodtu6CCuaQ4I4ulBU1BlxPMz0hGvoQD
QXD2FvKcRej1/T0Sot57GIad1w4yVG5fTvLKKbAKngJMFA8ctBbMSPEycNM17kVAkmuuXGi51S/E
jKpl03W1bNOE5lBEAstSZIA8RUeA6u46ecDC6UMvJOQEwRKIwCfSzjrj3IzG0g3zrHxvX0UVfnod
h4tNwLuiEPnPnPt2HOboeI/mOZoA6LXgmKluqbnUlXy5sBWaO0RKrZtCJE557Ks8qi+1Hg9I2AJ8
iEH4oInIV3deLdKGN/BEsKybuP6SlIey9+bN3z7/9IrESlAj4hzVRGLbp9Ybf7fCjfWjZmstmw2e
mMy2+H0qIfzZKpFyx5pdP5zeN1FPEQH84sMUBylRsKs3OUmcxrgYiJejCc9VLYfBKte8zqXG9TrO
wUbtEa+RXGoMtZrdExjFzPYdyoiqg6xSO8DSCMnQzqWwwdJRtjV3ZtUxqOBsELICej0iIBIsl4X5
oe+SrKQNSbTy1k5OXzzejivEv3Xcaipr63XoqhmsXz5xV84psdl1zyDpRVoZU3jYqfUUjkVsJlWY
Y5oyrufKkq/oamOTPKa8Txjt86C1DlCRMfFpzdBIU9cwYoJygPeRH/jibgATgNCPAscnv5Sc9FTj
ZEnVSP73nIrbbtHZYYiszsFYwmmHgcqqjM/FbMiuLXOqwkMdCrEmRo40+WQemwjpsVKN1zCHdH2v
c72xdDDrIH3HHbgYTp+3bcWCMbWEWNTw1Oin/1cQAVsqPSyKXSwkJXlUY/oZntnp25pyX+CFuZLn
20EMHZr8EjkovMGjI0G/s+MzYs6Hlct6jlbS8XyUzuNDhpR8kAWaZHdXjm0gnZ6JyU9nN3Ru1px2
P21UdjDNyhIJtyTy89UGzwacXrMMthjsp/pUx6FRn9k6GCKx3+vNwMkvroFoCoW4hgKkxF32oeQV
wnTW+LW6Atz8ZEoUD3GVB4t/G3wpbXpokizl1RaG25vDzEgo2vNDYtONAHXAuMeUygyLJDSC6XsY
BY9Y4mcW/89jw9OPIQyzFV0NsHcjRNuZMC5JeDhoaxwDLBWycqXB1s8N5PNlnLbDjyxuT7ec6QkM
rHQcsGegivT8xdaBPeWb/fgLf72h2cGIBbrHqRjgTs4DGkhSNbpekwaryKhjqzSP5Bl3B4+SHMIn
h9GXsNGL0Q3FWrxhMAukSQqDkfMPUNo/+KMzhBVPsBFi59pzay/Yx0oP2HQAgoTiuGglRrIt5Sh+
jRrA7X82dkdya1Ie6270sEt2C/Nv3t7e7yt/v2rZFOPyw4+D1T6591GKEQ9277BMLcGZNfCm5UYn
AZmSBIRrSg31Nxi0PNtadjq2YrykXr/VxDM2Yp2DraDRZgkGMqkSTM4IgfPDMO2zI41STnFxx0eo
1ER5be75QafxVODHUWmRn3s7xJwIyFvxfmH6LM5LzFxn7PeYOatcA+BFbdNtaBuNuN1lBNP4h8I2
nqoiYBjquKdwvZHms6ef/2oNfycpdwLJ+SCLsnxV11ML/8gzxrm7qlfsRV2p2Nk70Bve/xemnJaC
UrdZQYZrMzNYFMATjX9CSfbYDVPxzAcV8543FuyYFLnjnDdlCwoKSgZb/+rPD7UhnPxa9r4yocC+
hJhqHyc/rJXKmWRIpq60pTJeoKgPz6PkhgIvLtv/yPIfVS1fYEhFt3x5RuL8jogx/CUA40TuDdm+
QP+Kwn+k5Qr8OtdjYaCh6Nw7lpU4ieJ2A9ia7FafZsY3jUbT0rnO8Ouxqp9Mit5fvBSFKATYCNKe
aawWT2nAfNyZvaNhtKU4IQHWpXTy5AVnz1hj8MJPWKrfuPuCjtr6PJQr5VVVKmstaU16sV0ItVa+
TLfvC7kO0DJPqroB3WCGAwEGY1Mboy5YwTrXHT15z1NIG4xmHwIqa5TPAVTYfi0dkdhaZA9fKlAO
NoZ5FPah8agz+rQrWNWsiXmxHg18cJwyHwbjlB8VO57SJW9SV5Y8FT6OjerRFCq97R1+zkt6AgFi
dmhzMLSlSpGnP5KCK871raiqFkFw7FmCKHGG3bbzBktAiPIh+ihpyNr8ro+dguYwHjFmQ7ju/nJj
+I3uL9PtEMANbZ4zgIm0dTQ1k47fAbLfhacRGei8wA7YweDNmXhNVSQI0z0SWZb3QbcC5eLvRMtA
IlUDMEj7cT8ko1Ilf3hjew9FkCEUK8RQS1PFcXJ65ItV7CxSd1YnwAspakHjufzfkhUCkmRkDluG
IZtcN58bm01KHhHV1fBTy9dNN6bP/eJEZzQevqzOIZMzowCX9LVzFp2sAtGAqg3WbKsHU1MDh1SH
oU/8pyP+cTZOs3P7r8gFMN8452UVqBujotfB4HiW3hvGhZGajim6lfb8Qa1nFDf0LOk5/bcrhYMr
cNYQqUBbOolQwLEyiIjEaBh89CYfhxsVHfEFIX7x3CnPnI43d6Tqg3yz56rT7ip/VWyk8wX39kbJ
Goe3pA1JxIimXfDVkk3I21v2FjVxs7UnVGXxWR8qDZRF4O9yFPtNsF6baMCbsWn0nrsm1Ou2q+k+
c/rOdjHBOrpRHqIf5G4n2n3Nb6AXJVYwHdJIOSN9IoknygU5VjguGsr2legfRDl+V7LK4/QeKsnz
AHsyXhtvZHb7s0dzoFhkoH6E/G4CoVNFUcUlUyQtNjkeoc6umG2XJAIcw4fhvkT21+yyYndZLO2M
f4M7b//uHVrKtR0Zx1Alh7s15Ku4mmh+KfXjbcPV7LeJ8auPslAhn1LROYaNC8AxqWiA6LIYxNZr
q21e1qP79GzHATW3QctwlgnBukfvfmOhZClMr1fbJ+zL1j4hNV6k2ISNAIzxboVheI86n5PwRGt6
OR3nJafgZTUVMI5aa8czw0tC8M34HYsoaW3WBP5KbOPED5OWXM/c63QWAOw2/PVW1pOfyJ7fCxe2
FNI7/9ofNkzrCbH/QJZZl7hXx76SkdHL/ZQtv0D6sXr+zhuzWgDEklxUtRZAXc93hwncGI9AH6Qy
pBDFtGaEl0nRktrhmbgXbbz/HecvIWeS2Ok9ND9ntfUJuBY7rTOf1STvoKBEgTIkiOYkOITvOuyq
aj6bHfWOqMQumJThxiXNMVH3V9kf62Cl8nFANvDTmb2bjP+hBAeqFTyELMsNdfEGAtXBGmNQfy9o
qkuC9NN6YZZEKOqpa5SFVjRpuwy+xxp+iYMpJNpdQohXiIlX8NOsKqN9xGCF0hZ7LXW9NoELgm4X
MfsnI6NUbgDKRlWidjFujrrQHMq2yj3VMMI02fFP10apsytijZSi4LtxGjRQh3oZha8zzwkcp+km
YI/fHwl3Q+Uyku1l7Ph54HzPJmMMTQSL8Ozmyig6nK1NQPWJOX+cMGgn+/W71L7cqARx9O4rLF0N
AbWz04Y7rPygwTvI39eHCQX9RTLJV9qOZuY3W+lswXksUa36En65O6+CJoeQKS2u1F6c3T6oLk0C
vxgpTk9yg2bGF++hjuXXE5n821jJCIa2/LiEJSQQNw5jiBbmWEb79CInwuq973uCC1B5zBsrTBr5
EP3ZXrRwuBonlJrHSoIGl9g8Mc31WyKu/m/DMNrTky5VVdvSgcgnRkNvnKjuIEDT6ZQ1wpv6xMDU
0e/MMq9gK2C+ksqSv8FmzBlaD3JM+F5nwHedvqREVkYxm7Ovu/W8bKzk/XGfrX2Ka6nGo2cNRMIN
Fa82GNrDfegyCym9DkEMH2DE6i71YPnb1qIwn5uXfS3fY9/nJVZPAbyDLi91hbXmtTu6Oapi4t9G
Wv7+IteBfK/YKBcDRbgx1ZRRX6PBnr5ZAVtehN7Xw92Dv/TXFzNq6fs/DoBpBA/SK7JsBi+9SdZV
b5dBesh2hXGhNG0aScd4s6VLEPNXgbauEpe2rasRhZGeBzIKHMScc8N56jiyb5Ugy/4w7cLzPBtC
PnD16odC+hNiNHWMqgZdw1T0DzdkDHivHILILaOzhSMwWlhQsPZ/5dipPy0pb0OhB+uO2rt1zV8O
tx6AMk8mUMyTUsP69TbgP+9zWQjHWPei24XM9je7daqBCXeaaKo8gtkVqmVvgo8PkFaz0WDmaZqE
8GSuCTRlbdtCHEW+HaZ1004v55H79NdbVrLQ9vp/vNTU1obFP/dk4KgIDhSG9WARBrsoJkDpuAdw
FEYnhFFtLTNhl8VI1gXrN0a/W9/5YtMn+dfOMeXYXHmLUdA6/iy+lmK+Qq7PyDXx9YpbpW9/KHAz
a7XfJHRixrhHyOAgni8T5QWM4nlP/NMzVvkaKco/gMoZRfBR/KykTocURsOrORK4HBloea0Nvo6G
qoiVPOcejd+YggJDmXY2RIEJaxQHsTCvlOxVtjUnD/nOVsUcoRl7Y05RyzIE+VKK/tMkEc6y+RmA
mtT3RnMz9pTz77fn7HtVwCpUWW1kkEW20dVD4efk2P1icA4NuUrRdP6Q0Zm74ReMBu+U8xTSGWPy
zpqDZlLsHFnrK0eyJKo6/WqVzi5OFcE+fjzX37C3kqOtjCSxk1T04SSbQhUzRXInbZ5HCkRzJbQp
fxCNFtrG+0JnZtfn7+ugRoi9185TRAZWSS+OspeyJ2eglQEjYhQjOr+sdPZA0SuzAzCovJt/XD16
LiHNluxWmFK9m6/3cYIgPxNH57NCmieCEu2Gd7DH/gjGHIil9mxcFdJf4tzTLNYap7F8iomdjfOj
lxfyjW4cxevhKxF5QsKzsJJnBDYPL2FL3c7qji/ribwRra4MEdiJa4RjYz4SZayvX4Hh7lYC/hf+
lOt1NIeQCIxGmq7218t4GNVUbiurXlOsC5gdJzAgLBA/h05XUZ1/pTQsfqyjmxS5vgAOjuvx1PWx
e6+905ihTqFURUDdhELhyF7KvoU0qBEpyHdpyVn1fiTsWQE5GScx2xxb/bgBdc3DEiG2UCrZmf64
cHaBZTSFBPpUBUV1Q5kssTOslB36mglXqLECozeuwlGGzrdqJ0iMUjn69AwWqi3nu6vb+C7WL4pY
3iUISyQdjpXklWvslTki67dO0seWPW2WRB5sNmzqQZjDOISsUMe5QFkvnLTNSxbQKdqgkFc4gum9
O1BOonTP0B8v79uIcKgQNAjnsL49IKRkDu4+cushIY0xq+4VLJsr0bTHaJrcbZIyQKJgnrTgmgyY
7Xs3M4cOUz7kf9/WcC7URdVQkKUlGr1LXxHUJ1v2iR7/kga1w5RRyDbV5NmvbjYyHSGRzj3WTQcx
cJio3oJCvxIiKY0e9I5xtREdQW/uRrtaGWgMcfoUt/JSB7EV06gRM+06m0U/1o4Z91+U+5d7Iyyt
aPkLKmmA2C476rDdIS0IJ30ROx8taPrsceSjvnG0x0pplrCAOQH655AomNT5GhQWA9AKhjOfPNkZ
apgJi1Hwy9dMS9Pu+welKS+1LdpED5G8iyk1WSbyDlBS1vKD4pIQCEWSUSqOqPOdXDiCc2q+anrq
ONiNA9F4aP9WfAVoqFGs9sEw+LAuu16gChrB58wbnGSuxlIYlQ5zDoAi4kA7KrUaqX2Po/q6MsOR
qTG5fze8KzlzOFsSARelDVnQkLjOhnx4K/zecinAG9lKq31lInx9CluEAfws2QWFEgAmKC9ve+H2
NIvQedkhNh295C4X7edPciSZXultcDg/amFpooZ0LYLNoMqcNSXElnB5GOhLwYAP1EIOBInyhSVt
q985PRuApncld2je43Q7vNZXxZzHC5Q07JlBxPGFHFbyxEzjFlznImXYyXH3XSP30VbP5EjljR9M
Fia39W2w6AKoEgygAi/7IaiLItALoZNb0IX60BiFbstQyPKv51Vn1ORUGW/ZdBZAi/ftI2rmKdI9
rYrDHKQoMv5t676AbDlwmmfKrSNR7pDhKjheF/7R7RcreHKnuYBguOtzp1ZnDs5AAJl8bjhexR4A
5btUYYT2aKe8UglxlbA5osM42SIFpw0ge0VBQCv1sORD9W2MzQbQoK4i+Hs+84/Au9Dr7PX3ntYD
WoIN348JUN1mOqSXM9Et3fCQ6UT7F/wstgmBN/kXtPFXA6RNUwvZAhj6AXNH5E/yki1HCRShbZg2
giUHMNM3HY9azKTqO4ys2XCdSV7ioLPo2sB29ITHrEsOCtlNO6H+I3VBHatMeiwecw10vR4BiqP9
I40aAReD71JUAUa1EGJwG5rH7r4d4mtd0nyyUAgRgT383nIe0KJOOIChcop4Llok3PFjlhQkArqm
KwddnOmbz8Stkq7AUJl5+i2qSx632hJ7noFJWCskd53BD90Sh2VASBbv9baHGev1SG8I06hr7T/T
Cn36bFB0Hi1EV+JZuG5huZboxmxOyawmlbQbhjR18qB+ps+hATtLUP45PnV4iJP6KdZL7SfJS4h6
x19/WQmtPHWHU5/V7Ez67KBRBVGuTtHtYwVGlavXnbMNI50NyJRrkgA6LoPh6rukLOwM7MQyiQpQ
b+JALavwYueTuCNqgFy+n52FnUXQyR1LwF4gCryN0kABIBCA30O8r53iuSrI+rZv7jsp+wRBLGZM
HcPID9HME4pXonTkzXX9TubPfoy7pm9qDKenz7nAALeZfFOt34DXhKgMGUN8FyipoMelxdxffJb3
Q0zbQe8lcVvsK8D16qNrYgu+fE1G8Q88qv5OCWSC3F9t+6SPjkyZ7//RPCTp3YoAn5Ba+o4rZ5Is
FFmOzjemrRWirEnjB9qR/X0725FIRrY8o6p9KEWgVQBHQCr0FxsMQWr3zvk5qMmdkr+suwB2m0PH
GyM3s93fdO5ucBTv21pTeOkqdDXDd3pTF7M2uAjCiec97kvU2QRO8cqZe7DOHNWBKEzaagYj6bth
Yw/kw2SK7zuS11cu87+Dwd4sQUtOQln/OqTMtLzEzwPLCNLwrnEy3e6lLEfrbpsQLOjlQYVQvsR+
/TCK2B8ND1ZpJmKwoprc2KAqjAN2yug3VfmbyYQcX9DIN+M0UlE/sHKKGr94rZqyXLvVPfuRKqSE
Hr54mCR6ZzNlBXd2+TI84lC9DOpIVpOd2qR1A1Zn+ss88xxVv25jvTRkYa5A8HrEwKhD3ZMA0JZc
6nFJxpRt4b0s9kI4jRM8M3Hqn1ma9Nh1Fs0BO3G318oHCsQqmWxdyfeFWn0Oq1sTgBtzu6u+DEX1
b0s9M7GDNOXF/HSTPF5bOy3+rHaYuCNrYGAENxIIEZQf9paL0BrBLVyRq2H432p5Oqk2B0IfcIN0
Ooa+22Iaigh4J2bruOBq9XQvZsk8D7XXUvsESLsSU5UQd3aTAHbvLVarGhpgL4a5H5siXCvC79NM
yE0c0ORV6RTfBQ/RnCqlmDQMAn2GdGWA67HQdg1nlHn/yxZPTSSQMSbf9TEuend4zgQ3O4s0rXRV
2953t49VAmM2zhsPMDhZogJVJdFHupBKY4/qckbfQuMx1/+FHoQJZn/JyCG4eDW2tVYdw6zM5vr+
++PqLDQg+/MSTSzUE6JL7FldDmjRukm0Klt3XWHIULolrHi2AGmkfiwie1DHCaFjgvCUSIFvQrLZ
D+z38jMZmQEA7/QssIS1/P5YRAV8DrjpQxGRsFkK0wyymd2T9YAWrrT52oKWVX++YI6+sChl8RaK
jZgCVyQlWfetpaETuGIXnAol/EvAIUTXj2egFguNrKkHVsZdyKaklIzCRGadJEQT2JkBTZ2ra9uZ
WhflGml3riJ0dkLV/6gw/ks0MztxB7MsRmh6/+ToNgUs6VsnUol5dh5NhDblFrI0PMHHWXvr3eDY
q1Wa2NkiA20B4ycXktAxALuKsyG1LaoTVKNLH1waILyMEhAZTBA7VrE/SmSh/cbPwHaKSH2CRl50
c6wGZHGUO9/EcTZt00LUzGWKyHJWPPgiW/eW9o1e1vhmBkvLge6q8hZKV6WLMfIi94fYq8U9E2SD
Hx2LtI7K/8d16se9ZQUD/PzQB54K3fvPwxTbqK+PpgDlfjGrQF0bIY7OFc2Spaxwr3KZ6LFTQUc+
2HG6sY/o6DAcnjWIQLARBEXCFLpjT1YUFs6LHbd5CUYMhiu8ofUaNTuertp7+SKWxKFERRhVGQhA
ikfk4N4LXozFnfnP3XpsJKUH7fniEX4Cihqiiu8O6tsHW61GoMiWa0evHn0FJYw2TSoQHMxw+7sE
FEe9BuuWdcGCIramCuZY94+R7dV88eG2DatL0rOMyhRLTRrdgcw/uCIiZ7U6V07SQf3Y4GNI4CKy
HxK3HSDHDrgk8Un5ynBHHOCUSxaCyRQ0TIxstgEhPY5Ry34qn1WIPsH7uhAm4Nhm5kSoYscBJxnZ
eX8krTop7bqkUQypUHy4+r9hzlVna+jbfCVGPb7jGKLh/2FImuMrzu7U3fU88P47anfCMaRYw+AW
jMSBHwl6ZaEFojKv++3AMQihejL/1jGnrmAVRF8F4AsUoFE1oCsjJiaB6eVQDow6GnUQFUKNDEGc
PAxAA5vIELB60ThAw+B42IWhUpCted6sZYf6YiEwhx79hzRRvMKMqxJJqkXSaCN9u3HCAIoLHYjD
SBz2wBWwkmbX8MHTII3/tzJOM7tBRC+TuTNYW7SzBNMKK/IVVBOuIuQFlkmObMpgb6WpZITd5PdQ
9dYLKNRVhtcKFT/Uu+dMT2U0SA8LcsbIlqZ7xdjKvsPkRjYu8eJAEcPGF86+eMxyFdhXxcUaIpFZ
tjDTlhjQM6NQEISnZMxevEI9LRAUPlerPBe7ELU3YU7jhBHhhxQ+40seDgseqhiE68b6Is/wegoB
xxer9SO0NC6RzSOlPOpIpnGGTaGp+KTuS+nDp5R47immwVJLquWvGCxjH6PCs08cU9+cHjetW6p/
suG4Kck0uSTISO6NhKezY01gXvheyif6zrRS1EpRD/GR68f7gTsD9f9Qh8kXswGB/8HXglD/WnCa
Bh+SWrAoE8LnZ6rmsAeYFNxn3v0fnNBbDfwPPPt4AQzNv06SZGTgHTzWxBGSsQ2fVJcEcaoQsG1Y
GJtuqATzLguFrhfmdF4KPv0mye2SPscVm61EAfZigEZIifcFexVhahz7s3K5s+URRdYkVzMyvNGi
YLKf1FyszP6kV3h33P0MmMGv74pAa/znAzvG8Y5tWfGMd6LqIhFzSjR1RHHyefGSIuXNNUznpeNK
Ykb6IHFPnYY1nEv1PpTW7po5S7oRDAiN1/QRoONxYR7QZUMIUKouN/xEv8e4rZfQBeU9FQpjYVol
ZcaagukbtxP+tIXYKa9X16crDLSlGWfuUzEnF5gBvfPrhvknae6I5G5enQRe5bDNnE33zkqN9ZnH
4ggj6/juj5WbJ8Cb8KL5XOiUduARBWatso8qn7gfVj/iNWuOpMHHw3lMaOm8uQjAy/lr4DM/YLGK
QHpn+ZXxJsTZ8nivp/m+bJ4CmKsV0o4ZmJpYZOqvQJsp8A/xq9ISe5vUptz+yJ1PNwU2xmEkUzFp
c0XeB9sTs41zJlNOrpALIS8k4cit8N9Ri0hpOyTeRqt9nf6nBFP48e/iLVXTfF/FDPSX3KiGQ4ra
fdYYss92Rh+STLVLtg2HHujYru7xJIPkTpDcP5LVeChrt+wBiTsfw+tyX3MjPRyGJ/qO4wlJWsLy
K2jdLaHiP8kFWiVASNY69V3g5Eu++FdHCBf+ItzZ7HANHC4aApznAlU6u5yMilmUG2IK/NaSNKHe
Q2fvU39cTkm1d8Z7rAw7rhqF6hm/u4Zur3nNPs4j7SjdIiySoEcGtmnTqn/VIWXlIF7Z6wbMjv5B
/tWQoM1UiQyJZlJXlRxKalVXqUSCTkB3wJngyJ8JgOi2aNxZnLGYRYHAV7hlpZu7/wjXolLujVt3
K7MP5FS0D6Yr5CoeHtlyLMX+MbuosSr5CVQPDNb4Dd8tsn66FJMozQ/+Ng/7UZ8sQN/oUsTzFT4V
5NktaflVU8A4foC4qj+oedsBK+ATXAQlFEnI/GvwmqAg2s8SQPSXwofG8Ba2qih35UR2/bZoOfGG
mmLc84rv1P5HRs6A1N9TWdOYUsqtZz5reBmAvoEmwh/wEL1oJr/Ube4PEEMt6KFlmF1GqBjdzkIA
1ENemT8pqbJBC4ztTefPg/mdfo1yusQGcdhheGKqxPI+nIpS5fDp1I5R7ZAuOgNx8pbpLHeGxCD6
3EOjFQ4uLC1Jd9Hsb6vfV3Aifqv6mRBCGjY8pFTTH92cSThiXCmNYg2u84R5m1FsyRKQwpTCd2RC
Dx3a+qcPQdcaOfsuS/WfOu7cRs2mEZqenz8+wwByvcLh1gOihfC9CnfzL3zhM/hLSDZtit3/wh58
CgvUsQclrd0NbDusX0/l1Mu7Qu5iFk5DTUcvoCvLtI7MlEkkK9OlmyJfWxWZW+AUCNhiI7ImHqX2
Bs9VRMOhquJNL7gNXGLVcCb6ijQ5ZMDAHC7nIZXY0IAm7sjy7iWrSaQKLspxr3BqJlFM/akKxOpx
tnkNe6aMmpcSRWCtA7KsdartX4KW7NQX3EI7z09fmQnVGwtNnX2hfLNxuP3y406pXMr4AaIHeWmL
BuWOqqXpkcCXfRqNjnoUUQYmbf7PRcgUJTrB446/wBJo5f+LhvIhXExtjofd1ArHaMhUEMkxw+gR
EBjXJSZd1942zh9pzg89KLg9bUJcRO28QqfQ0l5gnsMNKMiMysKGYkHWsES516+hKJs5vc34ReNo
WRwqt2xFfKZIGJZuzwTJqgK5oM0CpUVzuhHb64cwWzvg+8THL5Xoj161p1OYBwDLSB2R9JK7QrG8
6xnWwARzti/UE9BegCRIxTRC2xFCTLYAqZ4S+U4A+W4tdHUCNEkfCoGNalFqTf+EQcxeEWMIANaW
TpFt0kl0mHeBEz83LWTrhOOuJOjvBeKp9zn/zVBM5OUUmnwgymdh9VNEHsyYvWdmII6WCI81ZHuK
re/owcqyWFCUA/gGwC2+q0b+mI8AsNRHLkc5agy6CSMFxd1YBJ/fqb2c9a4vREYJPm2xdWTWA+Wu
SVyxCATG1f4HMgxziUrtlFT7qby2KKmxLTjs5gUTpLoh/7Cc321XNnaxgGNP9wIVZVhDpLlycvmy
0MAExZIKWCL4gfjTiWKOiJggM6xpLHE/KTncPzKOesAGZ+EjFObuNeicvhkIlgTSQAuf/ItR32Wd
qQdR8IFxYr/r16fThpsENCnAhEreUSfAlmCVxNccuR2k+EWWTTIGDSq9O9nV0CdAO/bs0TcqOLm4
SmWR1N6PsZrkmCbuyejSWv9971k2oE2WQimGYevMrCM7tK96kujwQZxves8so6N4S44tWQyAbFqS
Weq1j/Uq2T3D8Yca7X0TFtAhrGd2fs9p8fOJcv24F2BOk4nyzJiV+qa+9IZp/2htOK4pkRY5Znx4
/6/IAZeC90MMALM1xoJwM6GTljlY8HnViXtyyPEVLCcyV0BsZpjpOrP0RnvqtaGW0oyNyZEKE0um
1WO/1nNyv49B54nTgQq6YH1qh+3jfyX/ir19cFH63iEYhv+LtFOCxckFyvH3/MxCzdzyYqyieJrC
HAO+Wymx5XTYMiSY2c8AGle+Qlvk5mawXGFdl8MQU5KAAEpXTINEr1jsJ3Q7boiT9aiXVaXrCg6H
6kU1O2FgT9S00NBCkUIMHSqS6Ax/wG05fP6fAeUmAa4poS24nQKBg88Aglon5xOxWawZWqae9nbd
P5vchzBK6h6k32tuf0CGq3p5kHppUv8rj7Db3UBbWC41UFWyZxDHSKyxSQ5zUNwuxGfWu5G9YUeA
U7XPjHXCGE5w53atj0nDAk6c0TgAgC/Lf2BaGmDzZcKkD9xsEgQUodVlyomNZd0QR5k2uWcUTpqx
6c+wIIo9Y2Jfv3cf+k9eaUNGKMHkuadqgHMCzwBrliSeK5FMlkRBGXWMjC/KOc1v8QLgXR9eTr23
88PzJ6oCIuwIa1RKvTVn45uMI5ixAL46phKkf8f135PzhvtLnDs58FlgoPryv3XTSQ61M38wX7Iw
Nb5UBKvgdZMHowgZeSziGr2vXjg9fWZw5HbvvBgdW9ZyoIjxjGEifMYVuGDC5DxYfEWa83+StogV
Gotmvi8woXLeDTavyf7Teeqoxme2IZsi01z/P13XtAgIlrsCzd31+S/qZ6nX3Efmll9sa2fAnwmT
RbFQVFjRLSluy12gbPgy8xr08tUR2FLmWQwpgu9+x4gNPs7HXjarqeFtIzVJiWnJ9f7MKTex/lyt
f18drISR/jcNMj9/wYG0z+3XLgzeFfxTkf44A+P15CiuEYDoSMMhP4OKoz4e/iHyqCFXP30iTfaM
uBhNtPnplwZSBiWG0dEfwD5Bo2LMjZBt877U+t733OmbJW5xjatOyL+GRZ+RY1RH/LbjkF/geUuu
fEmvgKwpdR0mHqt5pGPx7gHaBd+TgzBXuqfxCN5RbQrX9TAI/QYZFWBYvImgCFTRB+XDPTo3pEd+
o+um5w9hBqpdh7XXoSYIUE1CAE29kZVMatbvz8Y5p3GPnS2VbS1D89pVqc4462oShmnsAufQM7z4
9422b3wacLSEs/WY1UTOlZvKddFHNLCmtIjOjObeWZepBvgOgcBtZoYcHODTTsTaqbVGfuSiZQTX
FuKLQYCnt4oef/rmkUJwdsE8zxraOyj6PDAnFHZUBiaLyG55GbOyiCc/uvy+gJYU0Ee8d1f+KNXP
V5j/XFW2lMcYtbndSrWpIPGQtn9NuOWHS94WjBXQ4sXuBI4Rcj5EJEV9h7sWDK3qE4ZiFbHwlFFL
Jc9vq78kBLElgbyc0AFlGUyeq7QLUgdXGg1aQbRNPWhW1B84K57n4af0FxOLF4g/5hBCk7OKWt8H
/9UPNPAHS+bmJiX4PJkrjiHpWRHRUvuvq18CWqDz6okX6Jf8Hb4J5KaweuPwC1tvQSHmKiKVS6He
nbUxBolDXDYvqIZRb9Y7tVqeEtngQXBP0VgEUrPwjG5LRwpZTQQseq13AnqGCs0ZE+qaRwxjQGU9
gtxf+HLjlfEaKV9wo+1kXPoiiYyj58npOyqfNWUuC0ZYHnsyYJf5aKn4BbYkJcj3PLKJyRseH59+
1oyUPnu4AGEs61QZYW32IFGv+wZCBS8tH2LWMuprzjbAIk8uXXiMWZW531FbX5KJVUjAy6TXPIkT
2P50DLmKGDGys1m3gCWkLbHHIK5ZFX6ZXIsX8CDoJm3auYp/X82hefqiB3Ii/Kqr/zHr1G6FakUI
KsCnoJrZbWqsC7FAAWhYYVK/YDKwyCCxzQmujC+gVVyXfRaUetquKGdzqrIQvwf8yJdcjjsyN00w
nLeOkVn0Ui//YMQLEuexH425XuehRT0bSBqecYXnKDqWeVpx1iKq5LOoVwhT8n2FrLw26hXwH2fT
WQN/mvy/6L8Uzv2LyWSRl+aA33WVWC9bCVp/y1bgReWCznsZQgSccQ2CR1s6Ue8kSJB8KnMhc1Sh
3fX4/Qa1hGY3trtkp34AUl3omwVo8pyRrqHVqxopu4pcSAUBKHweoXvblqCazGE7ouJBg4aYhBao
Sk21XfV242IirnyZvBHvLA3JrCCOVS4BTROWQEgIJ817EuxfUN1VMmtszq01cF5pjOGI3fuQyMJa
hfaI8L6BIZUpq0cxmejWqvgD4GA5x/MIOX/mOP05tX06TZmAQq2HD/wjUy52hVe6zDrFyo4qZcFV
Vg+DsFsdU4ReygoT599b2JVdxxbv8Sv9fjEZQV7YkSO4CUzZQfKcJKTogULgo+DtHZuXVpFkS03g
diwiGhQu+/gTtqvIcul6Lr72uVyfbIrZqqQzOCMERe+MTCYhuApCHby5gy2D6N2YPoAdj2hQwwEi
1YkeJ6HsoShJ2R2Np/YqJ37H9/uqM/L7nLmPBYt3C2ULPP9P6XwIdrXfcjb3xjgcTdgqjbrQHmC+
Rc8vLvs9Sgor1tfnsUJ9caYAKSQK6ULdGNzmXWJDcueM8N7EF/zwrXOSKnHJPgJfLWFUz0tM+dxm
0KCRHzUJlpigfFa6Y8hGaBA6gA43Ahd+YkJG81wSW6uZo53btoyAZdA3pgeFVb2wgrSybWV7ostp
9uoH9PW7VRUyUqyIiGSCNurx0igLlh5/0Z1HXUmfwZgRfOF+gppAe9nCburQGdc8nxRdxI2YtvvJ
7+k4bSth0oKd3XYIdLDVW85xj1ZdLXClQlI5adiuEfvc10RxDg8Gp6k4Dh/a60DlFxJyjtjBZw+/
wTOIsZ2tFcz8qaP2XtgYcOvIOojVULhhaRY9kL6hREF1FH2fU5Ww+vWP2rSSLijz5T30GAld2OAO
l7jXQg5M/o3SNWqcGrgi2vBuNwtHsSyAT4gfMRDPb4hcjuzZcrw1UTtMnocZq4AGPPdrnY9qnCuz
45vMVV6Ypcg+9pxTRYpcad7lanFbFvRZ1DYERHa7rhioxmydsCJu992OU+sdINGuv59SRI81gBRh
SbnWTfpZaMDfksHwRm2E02i2nsMy5OpCnxlev+cmAf8KCh29TMlc2kI+9P4Ull4brtOlylt4R9rQ
jMMHPo7DkrsspZzyFJA9vRq9YiAg+dRj1nhdKSkVaVYUk/KK0NSqKEsj/O37Sl9VWw6lSeukUWr9
71C/366hKDhyTYtFJl4XQTW8PeGT3AEE8Ukf8ytp3b8GMSI20curzgXVlmGo0DcL6UFZky7/iDDx
m7vPhHAAFLTBx37PZOpmVz1RfFcJa9qLYl4yZPe4rzPEnVpofDHM84lhoLhPOaHfoDC8JlzGM7JC
a2Fi6Pg7bHf0gNbnGvKFObyUM/sQeMvJLatbHCVk+oeTUeE3LwvepAbDLcecD/WZjVixfYTpOBaJ
W6UprHU79eCK0O8hXCTz2ixNH5CiUomETLSW3b+gJ4iqUQfbJ8/3iLVjI3UkkZ0BYTDrjIjWX/xN
fF04c8FWC3KLLCHR3Tqw7eUKhDLTcH5xmFsbd8LihV6Jwx+7Y9WN+jSGDQHabrLk+aMgReNdHfrM
qxHW1LifyNfvMAogo98pzwNLTGLnYo8UWScsgxh8MV+s10B+9dp0ASyWj6S8youuZfz0Ee56BsJP
FYrxTc9aGt89BaVh7Cw7pvbZPtmmGnzJQqrozP8WPAfYfgGTtzNyJUWxQeTugmmG2Kn7vqzYwPjT
zK/sL+hRgU5gBPmg79Au3mskR43jSf6sprcXGCjhXS18mHBq5gy7yUeEqHKnXch4MMUlZkb8bhuI
DD+CKEkSC9C69CyepFKpRRNatBI956j20L4TXtPkieN1zxTYQYXzyOHqgjhR3gpt/YT0k0JboFkS
Z3xMKGEdkdIDnelfpb3lrU8f0SivroUm+mhKT4twWfrzciBCR/2mxI5vkV6Jx8m2zChdAzsciFXf
717rE4HRAsvWaM83fGsDSMSdNSU/eks3Fv+hvXUcMYPEi5n3AmpPejS4kExsynHJKsHBCdn5U5ZP
NRWl0N/sxvxRAxbI0gwaZHsFfJXfWzqQbfsgtMRx5nE7iVjEJtPJUjErxziDri87Ddh67wKS8KWr
MyS3Hwx0IIqT8tBB01yanjswG5pKWZdAjOWLkesQbmpiSZGr/I4Wyfs07ZGHUyyHEyiUwfsrP8HU
i9QGeukoyEwDgKIrk8jsJH/Sd1lNdMul82Sxu3p29fg+PtM6PrEwAgvqyK0Vbw7h9Dp/X96a0EsR
KfNgkEXwZFDvFB2O826pw2qNalk2yK4CTY69+tIXKZCJK+xFAeLM8z9VuC5T/rsDxq41/Vd3bloV
3uTDQcJyL5vMSqPLkK8b5FR/CigL8JyeaZbgypbIytvtfnme2lD1YIkNueOv6VMbPscbNnCQaKwa
zS+kplCnJ95NovKl76evKAMOSZERzK/MKN6cWtoMSOfKZvT4cMR1AULAUwqvkJ40LzDgx0rCoGww
2dW/iNqRgGr0pFVuP/24/TxK8eRfaLPcQtfccKgqCXDiewog+WslW16lje+B5r0FTaXiW/vtDxBS
mKT16Rex4B6yrnHo2WSjt3Kyg6vOH4F3cfzXhe/7X8AFlQ6KcJqPLYitAqdV0kW4IkJY8ZSQItee
IuPnijJ3iWg480Pc7OpAw2vITPc3n307o9ta1hLC5nG7s1aTzK+JZw5qWXutEYbmZmXKWSVjjtuO
Avr73C2ftkqoGaLyIwVQEJ51AfnIntWSiqOyJh0Owzlt7e868Cz2wU5dm03dPUZbOgyNVy4hX2O0
SKacA979wJ0DI26jppX/Cg+4HK1QSRgMqU6tu9HQprmzbhEfDn7zUOH5/oD93wL9T9dEctQ4kRDr
7v5ZBPfpR0h19PAiZTqQA4+LiFCrdlUYDwQnwb6i3ufdq9ufinP0tiU5E/e5MDQx4xPmMDeQD+4s
s78QedRfgDq5tEzEFa69PRSpb3UtKEbNWlStruqJqCnSEe/Xy7sz1e96cCHgPqJSpVzBKTCYsM+a
BpJVQD7hNRIb2PcYfKZXkdgSTs5qUaD3EZXjfVOVR2ss00D0pCtjfNWifmDdOKMDGp+l8a4lvDwZ
PYpEcPfVoj4zMBvnubi9qDeq0ghXjhV/5Ot77qip24rE/yk50jmBQIAEAGmbauufBn7FVWVdm4MJ
CXU/qrUclwRv2tTGEA9f/jQKe/kgPvQuaXFkYq5ecKfDsvmhdOEXafqN3TS/PwCRbr7o96/HrZgZ
S0IsYOViMRczNaDS57Hr+ST1zcfCi6rWBe5/ZzpxzwYUBlDDv7ToaVNQuVPp0ymXEE5c4u/4djvR
tPGoXDcM5jupRKQoxF4UslNmxEAd7IfqEcZd+bus+KfX61OgFEFrkS3m5wMBRhd3puHwl8jc3cej
j4iRBSUQfjCvTu8wMlYWFHKHAmn3vfSpzRhxBgidgZlWwUFLOHgPsc1Fyhy2ZfMnZL4kZSVEyiSB
OcOUBhLK4ArAXEa9MnabVjguCwCchEPgxnJ66z78OJVd7lI4ap9S1rNcQExhQBHpRI4bgUb38Lpg
Elak2kozbIc3iOsQ1JpgvXlRbz/mOLkNMgwFOoUZK6tXUl2DIvXEF25IdujBZNh9oIiHTD8b0rlL
S2d5CHbHKR/pstSXiUBMxKNl2OcSU04FcZymxGLC9gWktDe3c+raWXe3ww9skB0GPLqZr8GWs5OY
2w7G/akRpHXBr+SzU088rP0ah6W71Qv7FqXsaw3XP+mi5CrvKPVrphMirpcK/Xrj+6+iB0FUl/tD
C8Tp6LLXGYAVZksJ7Ky+AcTker0Nfp/HsMq8mdPaGIXfQUdv6QG4boiU0sPHwXn98hlxoWlQIukI
usWeKl8x+1M60PSfZI1uUoUfwkXt6fUBbPI+ttJv4Lihpa5UWJXaMF2uIkK7aNLK1frQWBG025HF
OKN/UkZVfVgdzqGGivM13DdOSRGwMg8bIBUeizUbJCkDCmboOgQGEyhS1f8fh/CKNxHrI0wROu9Z
j0fP052OyEhelIfqxhf6bb60Fkk6xe1EqruYAT0jcppeu3HUx3G7Z7TLmneCTEX33SvwbIaFbbhX
NOipecpsKpJXJRXzpJraAynAFc0SXuojWIdQP2t7Wchu3MIcNJIX3PjZPnolqr75gITM/uggra8w
Rry4oKVdvbtJe28cIefOp0FcqJR3vVGHW3X49fVNXOcFUeULjkJIfhtXvaQt2BAXxvEx2p9S7o0G
SMCdmYUzO6txVittASy/RAieklpWMGdmsrwaFI7xDRZH0wsQ1IrqXbvviQfZRM4Hlg1b+IZwoLkV
qHOaZfsXoNmuNtzWgKeQ8OjnbvudN0M2OGvc/GbVSDnZ106Stbda7CLZ5/72PoaQYGjckGnw78zy
eBU1K1x+jChshV3id4or0fazTWwt6YmLoj4iHZJOTq2jqtR1LowMeUSXcvH7TjHeBNywpdOg1Y5w
f6PXMiqMKWoCbkPfT6QTQawMt1E1a3teUtNq9qZddjG0hu1TqnYDOuARnhwfO+0YOJ5dg3BZolri
P7Haqv+IxkSdXxzi12h5B6tk5+vjvdpu5Hjh1bvO4tuPgDh4UNNw3KzDJJstL2LbcuFPReztZ06l
IVKQ8PXYFsSpTDK0v1/+aMZ24bLeq1f9gPiJMxwjPEG6tmq2uR10ss+NWgcALOFozatj4I8jlSsd
iFzwoAZ1TVo4tGUsLmTb49/9l0ckPpun1Smd/p2zlNw2ZNwBzY9+hegNUkk1zN95mqNpsbp6rCOZ
7NTtKgi8ufjDLRg0lU1mX0mXn8Fc1aREfnH7wMEem0QmlrrCmVvK2AY4UtpFnmaS5N3WMXn03Yib
DuWnkep4YK4ZiVRLwHWNu2pMrjh30HLx9wR/djqZi5gLD7dhnL5UMSyscuVQNjczZfng77mdX2O2
a5aHo5wkpOMXT5KSMu411nH46cwNFEu036yk80e2OQBLwuhHS4C2gG3p5jlsn8ZxRLLF2bNBAERn
fnQrDi4UBbGmVsEzSk/WsWITe7ZyVQ6km3+eUy6oVos4Kkhd75xqhFNRYRwrfyXJaFit+te1QcXJ
4fWRGDdZEUFQeX+vm/uQAr+/apwRqqxGWW2oCqUB4mRSv0JBKiS0FBr+n41O94L3k2OGTYM9Dfe1
QFdMpI32OoBy3tX9skM69GPeK9gJ2ErM9GHEaOK1ktm52fpYG714Y84apvoggpJoZmkbpZxhgbt+
p0F0zyQdxb7Y3I6u3M6nRhJ5TrEVxwZTb5y+kEMO/AwndPCctvWsKNNEHLcSuWjuWnkvRclxu7I5
aTGC3Fsb5QG6PMaax4VlCwogHfWNeeBK9/9S59HvtzXiCho1gAYMr7D605I0wlOehdiAIJH6m6ZD
5X6KLokvw7JsKEbmqGB8eON8rO8whH9m4uOSpucscGEJ/ibyGQBYqI73bjW75s4jOR/sHWjywQ4t
MZPkrhyg3zRdfHWLLnEpp5zsBmKw2MOkF92Fq4/z9yDEgYTiS4hzFvyeZk7nc2F9+U9efHEeVmmh
nCt236SuST8l6q5koq2ukpyHVPj0KRwc3KjozcL7IcHWbV5jURSImMImjUUx58gsbn9J12ag3xR/
KS3TQTAWa+ayx6/a1e0kLjG7qinDMD0REe1yOlZKdRHXzeKPHDLXgyI93XJO0lE/gxnYbs+FR1L7
o7qwwj6Y8P4DcF4NqzYYJzfwyQiFA+TBqwyU+i7wxtvFp8813w4XGoNNiUr3jSJNYptGtvd9XSa2
S5Sf+xhLZJwkqHvHjTRSSdFfpIAVKQqz3psNH8rMAPP4rYAVeWuxnvUYh6geVbsJZfFCyjxde8r5
gdc0F9TwoXIlQ9lac5vHXv+FyJVgx4HEKGCr4u6GuerjAwE6E3WHPk4dh6cWkjWP79UAMXDHa8tG
XdhZi1msQE37YIxiAW3w6QktGucl1QMEe5izn+8+v1ilK7bBrrbyPJqMITA+zms0VCOZmZLwnQM5
fMxkTxHiCgByG7TSxmw/U/au7Jj5K0J4xiWlzhbY9Kd1qYQqkb9TB1u02SBgcERYEqDVkKliyW/A
9JgM3DglL+diuakvKgWk2x9X4gjSp9X6Udm4aw3JGxrHTW7LXynfYe0rETsD8U2wvmJHsns3TzKG
9fH3OxrLjFWDjVA22ZMTmcWL7fRoPjvdIqlOHf474XfWwvReNqGwd1AIpMd33RjqaupEzEg1DHKi
zVaJtjlxaUMMreUN3eeyI1ObwH7T9mNlvS605fzrUNsIc3s1cJqIW9Fqw54Ykb0qZzEFq9aufoOh
YGO7oTeVTh8l6oVsY+kFXlpV47bluXHzkop4Ov2xM9bVYB6NdccOH3EunhMXgvZs2tUqwyoQZAqx
X280X3XxVwx+wLsBCkAy4Nvl2HElodrg550YxT448YqkdSBgDVkuh9tXJVKy7UdqN8QIR+wMbBHu
cFg2n44t0q/MlSOUAmpFHTkCrCCeLrrSzUaBGf98H5RdF3OpStK1UdTkGIdC2yrThZqHADLM4NJS
QghqORyyWT1+JLFBqRs6I4JDeTAxBmp2/i+9v6dY6+njK6cMBOb8Tdniw0wT25zErxmSarMK88ab
0vk24QFcxhPfn0F/TpPBMlz15GZV4ziyZfgFSQTmFL+NVS+Fev+nWL76VHsFIJE48RuVMKctgO2C
SLgNUwsi9oBTsIjZ/Vyk8+nKGICka/9JK+picu/JDoq+xkLZBWXJpOPrIy0o2HShA9GCckBZXRJw
7MbSgJYgGv0gnQ2BZyUUIUmUGx09Y4x6WVMAxLXQ81mXflli+8j6NMtHe15d1vyE/du3c24X/UBf
dY11wOHyanB0bEKakNp5uowqSei8acwT3MdpyboWiSgdveme0SUYn8hRblZGQmqDbd1XI3qwNnVo
RPLylPwdL1dXPpjclyLcWrtRzMZtp2l+8QC9vn2Y3cdkfwXdu6oklCy06e3lIVUsuUqbGYiJSd5I
NIphaR67UmYSOmKzAWXwm0MoUZ+Ii4r9jky8bwRL0gdr7JyLbqzVWgAJb0kvduxA8M2PM9oRoXGH
YV9vnmk5SYqiM/eveCdpuGLuPbs56PSEwGHqPeAaRDJt8VmjRrLBJDiDZAnqAY2EHs800Rm5GXAc
sBwckGknp0aVIY+bdrWcmc/WVn9ajeirWyf/0HprHG+s/kQv/dw79F6mhsqQCpdhwzKNs0BnKPBR
0u3tmA+lcBqZIEjaX78Rf78yn1ekRLn9cXmscoTzlWZtYjFw6vlJIzJGRJILUzHyTXpMeF4KSYuQ
1Af81d21HYHy/Cb3ppdklG6B+INwLmZqD/OS8mXNsH5Ckobm+ryCYFK1Ycw56MgM/k3AhpDBV/CG
eVoUVPKWolxx1uU0bkUIsYPAggBemqtZVSUUOdupGm+ndeR9xMctdfO7hMR8SBqvjY6Pt4EYIX78
2+JfXP5llO7LXIaVZmLo10E+vEFehG6HJikq1tlUvW2Hcgz9b9nrDN0FCGAAv2WtE+0mFACJADvd
m5d6fNWHqmQFm5C+9rdxDxMtfg0rhuYlDckAM/5xhtnHiVO2haXax0TVL0mjENfv1VFdTM6r9zNW
5IRwUQGmf5TjR7wpWX8sX9hBh7mnsL+p7MZeBOphp68d4CRo23qrURuE9Tcvxd/pkq/5GdaaTABi
jRFskKWH9lgj1UEn0xmmyhrNK1ANPvivBMaxaIPwJBwLwAMIbZQma3OnNNXhmjNWUXz3dn4JpUC3
zeHg/js/6L9MYfMEJfA/mWVRrUMWzOIcfH3zIVN9TLqUsArSva5GEuHISvyAU/EV/Cc3n3rIxdgp
lGlY8y/g3YUb3Fow44U8VceYl0yTNSEmLkOlKSsRgbkSrTlCkL7KEbN1YvSrjd1vqRZlAPALytdg
kVqf61aznx8i3EDVgYQLNPPUmgEU+ZYh0MUrjfPJZFELFFJ/ImOe3NoSCys9X1uapkJJAGS9uE39
iWPjOXdfXOut70qaCgAE8hs9mfStDNpJkM9N7Ap0YKej6fwkDroZ/FB0ctKZzPqT86Gphri/mxL3
RP9BKJ6vOR48y3SEAv8ThOMFnQ7bhh92mcC2ZTsnM++cH0s1StjxKgqkaYNVe2kqbb43s8dR2WrU
mXgBSVE09T/IiEiNGb+2R8mjcpk9MvDftS+J6jl6JPf2VhOjO7MVtla73hB/PZUnXr6kyL4bBsu2
wGFlwGtD4eXqyux8AomNyd3KNiSj68xXkxT/YNLpssK8h/uFls1mKwRt/zUak9BxN0C8BVkENUUx
c6+HakiBr5rqDFiVrgOSqWuKu1ewMrvRI9/f4sRQiso1maYSUVuys7xb3P44XaOtJ/q/Wd+dKKG9
wMAKRgahdDbEXbN4F1Py6UwVUglRKkopFLbv6Z2//orDLKn0ZXVufIOLqw6XineB7SM2Je2nYKjY
I1ffKk/UhwQQgm4xHxxNeGRzngKhuuRSR91DlGjvf4Y+dq3BMv89O5Y5bChzcZov+Fd8IP7/TIHO
/oF35pJp3NA2IeTnZsshydA3+/ichApg7G4ywwSPtT7LR7d813sy0r9ubi9KjB9YBXa/nqV7G8Fo
a7bVWQFyT5QeLKbypbdPWp4iNJjoii3qsqPfVU2TzqdySIv+F6mAzOYiCijjCBebND0dbdgG9EPR
SxOhpy58vRj4ebNgGATIrmxJW4tR9pHCY7Dnb8P1ZcaTuaV5hJI/NHGR/8n7iTEWr+RsyTPQBy5M
82BsGzIhibTkc/KvG4kONi5i1YXzfPpxdoSF3L1xMLSsk9ku2xPtwYF3DaIJA5ChaoU3COz4O1vJ
N0rzHemX+Fwhej+5n09K4NLp7/tFwWfo/hM3k8maNi0Eoy8Hum8r5C2QQFio0cRvJjfzeKc3wyXA
eDGUV1EyG2gcOkiHIMUIiO/JQfDps6XWR7mrMWUXfJ7kEFFy+0B9iGyH0aJdR150ssn+6Ezwq+b8
SLYYuwLIT6A94g5v/7CIA1v3M7IExJmZYXFAF7teKMmX2Jy0XG9uFKicjM/wVlGbfl1Um8tZ1Mpk
W4lL0e2ji7PxXIjX+HA1//P0mrBLG0r6GDw/KspNyVpZh329dtZP/OuadUIIogA1WQviXGovJfVt
4mHGMSPGJ8DWbCJooHWNbqUfohLo7sL3uND/bXWtQqjryHlfDNYxGLSncgfBkCFXVZuk6sB+mpYX
KGizg56OyiBkkiNsfm9dDZ47FOUntfDnXP9aJx7835PHtRGEgQ7wgorN1BwGLxfaGYsz5I+8Iw3S
UArq+2rhbsft3awupPuL4Sk8VLXoZfedMziwqExfvUc+F4t9Ow4P+b6R27RN6AJdzMXLbIaEc4qo
CC0elqsWW/e58a6EUtdADO/6rZbwrc5zfLvCV0LRuVYZfDo2iCEbnzds35GqD7JBImTwGODcFwwn
O8oD2xSruPKrnihxHHLVjzZhb0ACi+WvpaovPKrsSw+XyyAXZYfJ7G7SCGf2QE8IV93UNBr4Wc0F
TEcxQxuLDyLJ6lPKP6EXNbYZ2QMH7jhXrrCVVXenTm61DcFiBrZLscTuzkp6gqu6F4r82ohzImkW
zCmfh9Rk/wHr8HpZJTbI9P43LyK4m1cOoGfYrY2NpylGd7WiSRAgkMDyOFtCqDvEo7WQlluQJgti
voWH8qEudLHnsh4fsOAdpvxC70w4T7DhlKa0KKqItTgVUFPaIMwOpURGDyJy+wJw2eqWzaMtr0KG
RqbHvvTkXLzlQTE4NeSb3Y4KTAoAaCFGGdyBDwKnzCam0sHGJ1SIdwNV9QfhHNwtRxGDe2N/tTPi
+ryvwc5dsm8VDPsIHNsKeVaqtJMIg8HjRyYsqvDv8avTqHLBnyWeqIRGWmofANEPu0lfgCrESYMx
dQK9jom4XS3td0NSP6x00sKVpFLOUxRoEJNa7T2ODSBb6d+BzupTsDP61MMBgQQL+c2sJ/sFdeXJ
KcQn0aNKBnv+/mmG5itlUaHNu4UqOSbSK0FmxMik0jKA6rB8o+TEg1+6qrd/1Py2FVSn6A8/pQ2X
MMsZyGrjNvgXNSfh0TzjT3EPfNu1t7pmRDuy6bYPqmDw8Y4PC26O8JbZi8WkXyKdzS5RtB8eunac
T5OjEszKp/VBQitxxUG05hIYr+WhN4698g27cb5TvMAAy5U2GzhF/iHKpmHTUz+BXf4oW6iGEUDx
WZeYvyR/w53pTPo8OsKS4zeSBCwb78R9rEzgIvStG2cm71uhxTnPEw6G1hKsjWZJU/awabAQQCxj
yCjWk3PQmRquXSDw4XrsPKXrUMTW4YTItAgPIq3nCoQ97S+7716ORPxmgUh2vma2tRhfUxPUGQSP
9VKsrLn+8wQGI4X9/sT0Q8qL/GkxJHZOrHN18R+SheRP1Ku2uelvHhY27nlsUxMsSGL3erQgshcl
2AEVRy2yXQSHBlWYgvgvrNWpdezXhsAuf92jo/zFXYBwVXlcxpI6gWuUydbJnvxcGuGMf96I/NLF
KmycSwdCvEPIvWG4vCZXurluhvqmTLGOIfeIzouHpzsMcGyJradBcRX80ytJrvnIV78CmfvEOYlX
5xMreMVWLqWuKLsOarcFj/UllokDvpmak/ujxh6MgFh/yYTa7TMtpQareTIx03pxbGL/kOy8QFmV
Fsp5YzQv22XUbm2XFhOWyF8CglHEidN6kg3bQPLigriNnLdIfWR+jsbORvgwiMoFfNTdS1Ehy/ct
gz2k1KwIN2GUzFP5peuGojQL4/0ijsUwR6M180r/lLuMHpCRr5mKIvQapIz0fpkT6X0hLQ1jmnk8
zDS/n1MFp5YXvg8k0WcBqwRTh9sX/SnvtzHlbruMFyEpSiEAhVddk69Ojx8qSeuMi2vP0o4F98+K
riw6cQZXxv+Y0GFV0jZa6qtHPoN1wFwkd83NmKCocz4Rhjra8iUbmpLaG+JFvQmH4wZTpb82kBoY
7RXy8rlbpgV+uUlJobarZe6zp677nrjRa5UmET3Sup4Hc9PKJNKe19xJd2h9VJ9HaKgDp0GmjEDg
evlM6SqjFfoL4szhpoUt3VgqMsHp3zE0C2Rt5qiKAo86xMwHMfZqf7o34ZaJunBcjBpQEr0zIuYe
eFrbfa5+MRL8kNjDYL3rAIcT8QCh1fV28eHZVadgPMmbc60LTtQY9jbZM9UnBlsmqWFRIWA7eTjr
0jAYbmY2DEuhtK/U7CNFlN1Gt+dOULyql5bnSCxJyOSj2V2/ppOafedscjnPu4qigBA6A5gqyfma
a8i6UXGjJ095y6PHnbZG+PN2Usc8HNFi691qwDbO/TkGfm1M3lo3k2dn5GH7xnCqf8c3UGe9RlDh
+Lbypdxqnc42jc4DO1+wIcll0P3SUlyoIbzUQx0A/kAvSdtCQP4r/haRhvdr6oUvA6iCP0NXg8Jh
nJQaCNr2YpATkq+C0BMdmon2sYaFPZnYQK9shYp0NuSyPW0OANeUikOqSbm++zTIWRJ9VlyH8alU
IfPLIAcSmvZ89E/DIAdrSyojkPlOb4Cb4vYkIOLwif9hKGINwgpRMKzaBOjdiEzmwxNZlx/ehL8F
iHqM7xeztgqXFFgzDT4ya9y5CKOqjpA4Z2wuY/fjTIoKVfhf8UoXZsziQpy6yiSQG1pBsqTh5kXQ
zPk2ePsYOs2cr2w5vqcbmkl2wZm3VRo0UmUc0mV1blc5C0izBxIRaDfYC0K3PjwgrD0IqdzTxZQq
zvNDo4fkXKoYP7WN8vtLh2lddybc3SPrVT5RNdyZTdlZErZNJL2KP4p91wIXhWp0tXEGRNZzoO3x
bld6VeT62Mh88Hh70I3+ww8+4kpTfHg7s14E43cYnVhQpuEKRxSkMWdnkVVERoeluJHFg0uWjH3A
BdpmcTrDsEY76seuB4HppWFMI/hgEdAUZDdRFoyc0GXauniBhPtreKz45NW1UNt5xcEoPYwoFzjM
4JSvNQoeNEzg4VZHuq0/FeFCllA72vfHafbjlvUwtBevfaVbj5P3soqb+hynxpcj1QBYoi1Wr1I/
CAvqUfcqyg70x0Ni6T5NVb9iV+LWyuP6wroeiNGCw1dNViMUOaczzgFzQ+x5bExzD/mk7fJ2cdfd
nFXo2BvI3HP9g8b5qw7uAUBUXIuuAKDIcXXf099e0cZ3gEabzk/kbpfuJ6M/xlrDx3D1v7YImLmk
r3S/whTS6JvxfJwtK3lcxYumIqr3HH/bafOmsfB2a/ftoS0lrrGh7Rfq532kyF0UZWRqS3RFKwG1
DIAzMTJPAxSmgllOLIZIy0L2h4Q98hboYIG7ApmOAp0DgcS6SF64CJ+wJMZ5M6HrANhy1c8gYu3Q
vpA/8WKvKnermIQFx7yqW4/XXom+4W7UQ9+32PmUlXa3qT57cjaQV37aYc6tDJBD2qKurpEnVb1c
D0/mNA0BmQSjcaDoUNHqovGN5rsOQtp2BNR9DT7B7yUTJw1+hNWZ222CuzepOdCzwk2FbIV0QFmG
KQZ2A+9w2gqk4m+wtpWlB6P8R6bg8+CqqN4I42hbbcCD3Tp7gM7vT239iCjTFLLuV8fifYK0mtlM
5nnSqFL1C7qxgcGFZx7uKy7CAZUrflpzUhxjsvIBNtHHNAnbCjZkDwic6Sjc2kDJeJoeasnXOcXL
/MJXI4mqtZbUn9U5YAiMAJewnU/6h4vjcQsjCKIL2JZYnxjcjGsWA8ajr69UjNmk3xMm2jAb5fWi
EHaKhtF2ju/Dwflm1qx1tL8DCJyxxCd195WHu19mYddGyBmtzumWeVfLLzSCrtMuzGQNRr/EkmVT
WSVUk2KaL/hIFqsTfsJooaAF9Q1RbSCKoxEPY9IGpqD0Zh5mJIUJ0vuBaNM9aj6OBb/3V8qwJjlU
h5P3o1RmdvMnuJ856agjzJYcz/CpSrx5+DmcYoov8VeP/z/wsAcO3zwhgj4rvNqJRJGdqLJwvO1R
XuwyBddtVcHyklE5/8Itg4tyjVi/G8yF5qPGRVv2GJFaev9Mglc4jv1IzxGWjvH6OeMh0npXhyS/
pY1lTCf+IcW7oTtDGUbB8lXD4zN6RZDNi1ltQFJaMhiVm0XZbUn6VPBv6K9EcNcu+pdTMO77HhS4
iw3oOyIaVXMgaPBEHFDc4Cgtc4gBOlJH+AurJlpCsnjExcgvd+/3f/ARs7ih8WwJLk8EsPEQcIR2
yfeg1jtQxC9QXvvldCnTF9q118q4Z+4cF9T8tg0uQ1CDlN3wuRUpCcPEJoLR7pHXbhisiK24WyAK
2RZpYGHG70afrzaIsU59eTwxn65whDi3bz+fNT/0y2140bt2yxbcrIA9ZjJhNVL/UmmM0Wkqtj6Y
0806FRSfFVTAZmYblP24ETtZPD5CY7aASmrfoIiy9FHvgFixIfOhN6Pl0NaADwHVadZI7g1WHxLj
OhYHYhLG/O724JYu0YoQ73nyPhy7AbDuL/ALtwcrjG3EgABHzRdVkkXn8cg+wQv6yikkPYSNwv7s
uUDJBvcWEJIt/r9hWwYlDJXwEbPMJCx6qs+a9iVRz4ma4/01aJsXsQTOIpHZ4I6o/LteuNGsLcxh
tSNDQWO4Y7V+wgbWaUHoeXRcMAE7PF6Y1RTHhfOKGCjjWY7kxLuFPwndD3TCwXCz2RsLxDTv4XkW
pDs2C6htLQCzcM5mcHd+qwiyGCoxcQSAoMNgtJeJdPIVOjaktbWMGGslBHhIAZPMdVX9rdPtsaIv
lQ7m89BbkSEMHiQDavwdzsQ7ZBSMv9qgQVsJxExTeoF00q3HTNXqqvkzn4YAFGlE7Yxzq/XFYbG2
EmYEG+JwJ3TQKuiTCOKgvzOrbfBNfJEJE/sYxa25XG8h4Tfkf1Gf2hZX8tJy9nZUsmENnwAOmlUe
blvamCCtuwvnJBh9XHngYt5sciyNDK3KPRixyPalCR29l83FtxHgqbSU9Nx984WLLcLSu+hx/ppp
ZpNNp8r/8Y/6jQmb7ZbF/rsHEwPRAB14VaOnOGi+7TYtN6fsFiLt0r1s7LYr4CgYfae2Kz60xPU5
ncG784C60RnA7py+T+mP1hSGzN90bNeLcWacKt/1r/H8MF7k9CSrwFTaYKpqy/J63chIRwS69c4d
Mp6alQSnHlkx6/Dg7X43rtY8J+1CwzPZ1mopB6DKx7QWLYlqpv2yX+xV/jErz6tqAqLEMe3GH56e
K/Z+edZ8JulFdT0QmPB4VC+I3qj6aUpoe+CkjciOiB9FnuBT8n5zJe/2TaQqcLh11QqEKrXlyyTd
mQw2F6bJHn6cISIh9NnaqOVteHgsp7Tp/luWklr+ScIoHBa7LtUWeErZU3RPcB7A95LgRmkN28pL
O10U9BBcEiCvtH3urm2qw2d/1TQchtB/5d2l8RtPsBMw4k0/rXWGhuVIjrP7Dbu5nEBYYtKIhpme
SOhpaF9AquzV2CQVuZ3lT42e/WGTDw+NU3/7zAxohn7aThnkwoW3E54c23Lgbx9LhpdQh6919wd5
MaCMQ60q9L3vPQDcy2aR2a1Br1HGTCqetUbf6lLvLt67ag02+lAvfvQaIHmIxElSLAVCXl0H3yf3
hpwqj9tlh15mOW30DmCAFrVHY6EaE+0FYTa4Zx5BPZ7Jy+KuUPu2acaYJo4d+ctiWj/RwCd50TBR
o70Hg5E7inYMmS1BoC2VACNORIs5Rf07YwGSYVBqR7HcK8dl36jjyC7Dn/G1ffJtqFdkAciDXM9L
D0mw4p0/WEIWPmOghM8SjReANq52GwImiNhDWlsJxMcvT/sjj/TeTRiIxwRb/cCjbM38ZJqCd47N
ae02xsmVtKNgDTY4hDbIxfcv6j4OkDXKircYIuFqlgRYY9JlMPeJCeDMKXiAL8VPmbiE4+CWQS82
gZVDdYY7goymxx6D5tyEanSCZrH3ca8IuMu7gQtnxFYZdfTVZpMsH5uCCs60Z24g0KqEV1Mi/q+A
/xhjmgVC8UsSkVXm9qXtr3U+RC5TRnVWTKtfKhGxrYlsRJp3uGZMHnyxC8f5AMFMba34KDjQ8S2Q
IJno8hy+wNCVNfz3XeTMDqnJa29uhvkDiDimD4S9mHKt1zj50bYhvXhvo9DKOXdgaED3ifEFiUJF
7c0mL2RhcvqYNrMuNG3vXIgfIoFKuN32Ft6bY5Ed84uHipHSC0BCYa8wo2gCGoI1r0HCSmWV80fx
cDUWWp2zEczJBEPmKiRJjZo85P/6M5l7OK6VFnUa2r7ccmKyDuywQmA5VV4O515OpZ8s4cblB5xc
bNuk5w737fQKf/kXlHyEsHj5XhuZbsoExjG/SsUXNko8Tb1GtFl0IVWODipccPCGPYC1NbEdPLuC
cuqhR7zpVAVR4OeL9r1744W9uompLR63TtBmQVyafdJupK3brwStG6mXjqhUD/78E5Zwd0IwUmt6
EbLB7glKC3m1JMED9W80ZhOTvsn6yuq2Q/3dRy2gzMz3PGsTY2L0kBEhVOkkL+ZnqhcRMlNTLTQ6
9F+DPrCVG8XB2w+pTcQqorjoN8AYtF9y7zJzLszUygx5oUdirGzg8C2DIkldOG8JwGTPViUglb51
uSzsvE6HYx+ZmRo+HQDDE4XGatdCLddJv5ryGN+NINhrniyTaKJaTnPqCcRnv2A0kuAoIgStcjRW
q5PEYCo+v5QbrmcKY741UmcoAxrEyXKLDCLYK8L0LFw9FMrSfqtfc+Cq4RaDUxkstjbPFZh8hs31
3xJY+zHMCFgWakqxYAuLhdPOaqr7y1Ns56iCQ64YcCemgh/ffc6bzNmj4IdvDUMwg2O8SnzJULSG
IVsYCcKmXbHzMZSjkl4NChyHAmleR/W2CHX5DflwH7gpNUejeipgPa0kZUX26Mk4Ywlcr4d50EN+
CZMHTl4VKm9uWSwVPEL4OJKeqrJK9aA3DLHPciaV33vDKyhZX5TOKQ+BYxVUqsxnrd5iQ7XWm08o
74oSDoVrEjhcLYuyo4kNWFRyBKL4NiIA+uVgRV5usjjtovIIOqMbTQgxXWLz26m6o8XjuysQZ8Sq
KNSwnNaUkhONQwdZ6f/U57NwsU+htiRmwstMaD9Z6OTohXtuCtChqeMLRuUFKSAuYM9x2cFMoUuH
xOgV318/qThBHmK+N+dmO2e7dTwlaSDEg8xLbwaAKV11ekx7CLKC63kK7PWXF5a2fb9h5BwUQm0h
wnF9A8PKnTCglipEapcxVFhTtjulB0ROcOqDZlvorCj4MTuIg5BUR9k7Ir711w0zwDIEg3rpRl0u
cxyqZyPy5Z9GhfQDVh+6T3r+NCXqS2I8EWWe3PVAD2T5tc/gCiSibIwdur8KwEijlwUsqcthmqlH
ipOQ/Epvohpo0AX+WZyNsxGxWWC23DtXPraueBDvxrYFS9Dl8uor/LKdhk8RE9jr8w9BZEr5y3xH
YlEJDBMA4+Tq5AkJYfYdyyLSWpWbvTvEEFwjMjXnH2DpfcOqHGPhEZN4yL18kvvNsuGflKkVN+NQ
Q5Vo+uQm29+EATDYU3gd0AmnVJ1UzTPAAmUwCLLv+VJYyscjcO/H1p3ZqkWJfJehJZMLJ4ud7mri
e+Wrto5K4bpGy6iL2W0a9LIg+ZAa841TOAMziGdAso3TfVg9BmYcOLqyT8i7dJIE1K6UXyoG50QA
FheWKjUN2hVdP4Mr+fWus0Z0Cfl/HkXL9vBq5eswK6ZeSABNvAn6y+jJHo1pmZ4v28ftvnQd7A80
SpO69gGVFJjOC7uJ4ED3ixEMQM8Y0v1pKX+SyNboYXlTT3xZ+dbqA8qeYUJDe/gWX+nALcWGg1U+
y/CHb8d0tyjgQA5krh8Iq1FA1Gzx3okhK1U+YeR9cp9xAy+GokMzZizulf94CxdMt4WMdF5fHVxc
mjjFRQ5fml4lxJPwUxJLNppd9WlHLoYD0FVptvxM6YJYMOUGeI+ABRZ53LHH9rc+wJG52ABuPE79
h/uhI6xMQ3qPiBDeaHsIvEd01EGDwuUOlTGZBpKLNYaZrI6Ez8hRENCHLuWv+jwLaIRfTPclHD+S
Ufn+jx0JYKMFr/mxTRoxYnlzwG9kw6XlrurOMhPSS3i0+4IrrDaI4Mi6RfOiQ+CaVl5OKJmQ002e
uAEDyWl0UeaasKvLUj1JT4Ne/OG/iBd3dpr+WaPTm8vQwd/datN6h6iUcHjMb1rIg+DM6j2XGRDN
kCThIMHqB50T80vzHazjUia3AborV3UFt3YfirnfsvB6OD3ZNoBPBd2ObMJAJlyRf2Cvnfmc2eec
+4GQvnQy9iNY74yEFZqgk/wCs3gtwnsTqqE5cwWZ8Xoa/p2e0xgmmCOzAPl1TMk/AUeVD1ykE2jk
gs4+gXO3E4MrI+m1DfH6DRCxearfwFuvUeqqFCwJnQSBMb27ylzM/FVSLrfVxg871iH10a3d+jRw
bhIHCUcuu8ESHCGWMMORmXz4SPc4h4qjhPQkoW25dZh1QhdeM7xi/0ovr/lZKltLFyiCP5OjTFab
/dIYkMD16OLDkY35gr3HO2waRQhY5yjAv3iVNvLpjG8LUs7EtnEueO/QqSHKFFEzauv6UqbRWxdW
kWHagaweMgzqatd7DwpVaCyVCwJZuQApx94Kw1kZY3mA3JqpkVcIefMJ0BMAVcnXhzoIl908Iag2
oCffto7QROcpyA40DLqVJHMQw00lCSzqe9+XCLu7esbn9FySkpJVdniIfcYD1l9t50/q0GWIMSLN
cgEc+eFTAg9Vkuc4lEK6IY9G96RggToFnLMRHP3hErLfb7jN/lbUW7JZelNidcyUvglsK5KYxVs0
v3+CrE1rHNzHd+7TfksJpZT3B9I191G1XpxksifZdeSqJ5H+uyZW6KYh7CavlfWRwbm9rvTD9HmE
WLHQyEgf/CSAqECMTYXvVr77fx/xgLiYTILtOZVSM5a2BtCheGYn0cDx2xLEYleQqL2i03JiZmk7
HXRJjB/p0ks60anHH2goMj29ZFZWBOaPiyQennGF8XA5gZZ0e5b+CrNebDpi2XOZJfr4ViboTyBB
ggQiTeESCBYs26tLnP5Ji6VAOo11iUE6azzsA6QVgBdyeWnAquIQojyP5KzhaZXWKOZh9ZwE7hoZ
I5cpoXJ/p6MmVT0fnV3SXFB1xvYpFEhDAce9nVfPe8T30lRn2E8b7Q4xvagS3yOMCrfY4M2PRhkm
MpGf5sKD1jP9ZEuW3Un3J5feE7cS22DeP4/lQms1/or5irErqRgPRHrKuwWsZKLGcLdMfmDf9LBn
YMGxvCstR9WPa9PLNaS7ayZYiB70owHPZ+LA3R7qgloGndGF+rfnhxNUadnt28rdu8vxQzYoUlLv
SmFnOA/nl8VmJ8CLTpI9+0MukkTZ6w+56hdDlByUX/G0Y73WgyjjNUJdswJu1DuK1zRXhoA7pUAS
v1c9pnVOlkfOn8ak8MRFbjaCrDXEG7TJP0IGAi/GIXzTd3ReER03DdvraH9scjenpTHlomGmwPDT
yKzBPldFn5i1tmfwjwC0hvA/kSHSevvDJQh5J+5PZoPGcvfHfpehHjfF1GT10GnHlPG9rv2oOVZj
2Q/RMnmo7uZP4eyMFUGwl3/ig3lJ0ACbQI/jdu+LNizsPKwR2+oXkDnP4EdZsDkRn/3ZXaO10dyO
8neMMh9gCcrJU8I664Kqlh+CQXmhBkTQ4HjF+SJflE3yn2ZikXMBe+BeoIXw39JiQbK9h/eejm6/
Hf5zD/LioYgLoUZCwVlqsoXBVQtavv/dRoqOWBlbf0dU+Qn9c99EKX0X5/yOetV0jVXxoO4tnehL
Xtm2iTz3v5Mnd+akGUlx/Fz2ekKMIIvBuG5QbGI0jv7fEwjeSUsQ9SFyX5PaGvkJnkYppoMVpdcj
MklTLgsnIT/ZiWlbddC4/CakIj6Hli0pZH+5VTnsLHrdoBy4amCFDAibPhZs3Kjy88lEIbLMoBO9
etUswuSu9rxo4LBCvVl/BZvuEzpAgUsg3id5NESaOLqxPkSq8nb6wxrFTeF6ZjUCZh/3fPX1tpqV
UdcX2UzU59VfB0do4oNYmJPKlUMziVjUwwb56Xj4kZcUJ5duG64ca6i0pc/At+t0Bxx27kv2nFIn
gKKFVqR9Ro6Y0/aJID2dfPCST4uhFJ8Z+ttjjNfAAd7x7dQhd9V5k/mcYmgzFIOgmHPZNOhbNZTj
yJcqXx7eLQnSs/4bLDusE0dOv3bhZFjJkgx/LdxxZ+bQVJbX34FjBNrfOAsyDMed3N/xFD1nxClj
iYrlgUJQ05nVS6uauOu6ooP49Fy+GDb3DShjGd3ZywSc/xtdgo6nbhdrbrqagyrnrUeJ7mcUcPDL
RsID6AXhgd+t4oFlbGW1WY+AK45YJ87Txb/UOPMotg0xPgkq3sDQuKj3egNAlJ5EBSOnxp9XeUYG
foZFumLkmA6zw5sZB4Titm5U7dsAvxCTp0nZoulaF00hnKeCOHitEvnNlDgNrv3avKUfy3EKLK1L
jAjIs9AwIp5V/GieodzoQR7lDkU2Mdr5GtA59VmjMh7JNndhlf032N5o1HKXhJf0h/AQy60swmB/
Uh9roZFQwx3Iy2VSzl6sJHdEkRyHzCQl4YM5bzTSmbGCa/kNURh5erck/F4+jU/0Pek2gIaIDEGV
W4uDyuavfia0EWBBZst813JxfZruj7YKKcZDeOW8wQzjGq3HVePBGe2bconc04wSGqO1Z1sEGhek
wFnK0wAl95uR46V8+OT1r5RfVYDNJVR+LiR1bWBtagjB3QihIpHEi08HmJshLNwtrp3CngJBKEzb
XLS76xNjWFz8LapB4awPp/8It78+87iy8yUojKm3OfaFjlpEfIKv8pbTdAvZXvmllW9JWDCOsNwM
af1SxjSNJqdQvhrrYdxng0p9ld+P1HpGOASHe6o1F3Mx1+DmUknsIhaDS+CclXGvggUvEJvMvFaC
YVVzP48UfDwYd3LoZQI7PrIrBo7SaXiPTiX5nSVl70wdv5Dm3FK6Cy6Pji9dJnOaWQSJCa0sSdw2
QlN4MgCJrfGbVH4Lm1z19nNK/pR0DwtNt/5GSELSyVpqpVYDuR+fEWEDZwU2Pw1Q77LL8SmFYxQ4
cn0TGhiKUZ+0qBI2h5pBRp1ceLUFs/buEgkLYaMObXZRJAQghKTDoCA8nJ13ltO5KcofsuLVcSpe
RmT4f+bBlDgWuIBOcpS00imE0TjbNmH35gvzvhWwsKqTFlz1rb+HItA/+9UbhM3SZJhPnwpmAK/h
jIwA5oSJvreOR41ApPIgXvu0qcy3oZ3mSJzmcPEKqhoFs9uWSdsppWDO4/143AVSyViAVOAaanPx
v/qLkoHzy1RmQjvCjQx5Es+KWo+lQRglnWycbmGl46XkXtr/YkgyGvs+BE8cEowSNMiEMzSD5u0b
068Dqr5KAgyXX6K3+NvCOhndDR5dhbItkmSigmdMvjYIs2DKIALchQGAgp8kbANov6gp7TFdNpaP
KkmK5RQ5XCMdkyQnwAbN6pYQbHKsyFFWQ55qDh10j5i9UmZ8ntrY/PVXeZIbZEmnjeX9xh1W99y6
pyGbFFZRsDBuU9KfSvLcZtIdbWClBL7FYdd9xF2jzVH5YDan2DVkg//xBtVtPsSLcRYva5Uoeh0f
Ikc4WbVCziz5nSgOSrH7/4MNYkZCYO4cevWAuuOREQO4R9ONsuWnyhiTTyVjCe7EtoM23G6YdgBl
eiZURchmttGlAcnqcffD1vKtY9OK4sLu4QoMFeAa7wQqHaOgCLav/cVytTtpSD26WhYlGCGh49vy
0wSc5Y5Ehl480Ywlas31iZSv2S4FJ3szHTY52Heo0Le5BIaKjL9MgnzXioiN7a+znfAMtbsZSuOr
/kn9NK1+0cx0ebw4ziwvM7RkeLkNmjEBm23M8yuKDUcto5hHWDecTevccoAtQf1mZEJA5TAw2r8C
Lv8ALEvQFQp0dSRFqmpg6TjZ1QXocXgvohs4Co3kfdEyzM1H3589ki10TVmDLAV8pcS5CFY6GbYb
8i9x54BWn7xoBLTzpSNUpThBqR08WCeHTXCnJgl/JF0f2gJ5hOWTWjw2oDbBa3il7ueh0JUj0jSN
qTGO7HjDWYqqmtkSJ8gcieTdptwNzP7o95nU8SD//GWj9DRCNOv/nw7B5xOM3ep+cLv54tvKklhz
6FQgzfNrIQ6TalIi6HjnTcZ4S2HNsr9Ik5U23a/n0uurii44+U64WiGeXgkSB42fqdxrIdltHJuH
Go6YExRUjpvqJMgiQoGWpdMZI9WCu+pXrF2WNTL61PIoibGFTq0AZf4n3FDpmo0rywX/LtSjkcAy
ChMGU5locYK2vc8HVeH++NvrpNS/qamrary90O+CXgCLLspT3QePYvrdk6WhM6OGbM4w/GMLQ7ZH
XuZhhf5FREVWjc0wcLoVaeq/Aa8MUHe1nW6r/ejQoWC9yMC/t7IuxSSlicI7J8ac1njY4abOBzOa
fPVG1x//akBBQl2BOQp/VrAw+JqiLZi33dNld5m5a3YEaZjYlaUI9f/+aJK9UWO69r1S6t1ZROaE
/90qOESbTPB9Tas9SxkHd8scxoVu0SKpeLmfe4MwoashjJWDAVvtIScSvBgKBaPkeO0tyStNVCs1
a4g5DFP5fjw8wNOwlMJrlZhUmpJm+F7+2S7gZ1TKeO+rsKzl/EozNeYupjQeq0BZN9cV2f9WsNUG
x8rcy3bOmdXJr2+gwJ9EFULlGedBDxcwaXLlw3sNXBAe7QUigjCTNH44Bm9QWRAXzJvl2MOOfxQU
GL9Dpt4dT8d1qj/ffzEcIWMFr1gIA6j5JebK6qoAS+Qw3aD1FYnM1u6Tz+yodmUHTdq7QfmmoULH
KppXJzzh+s3IvSUnmqEjppx2sDolfeSwKg9nGV+ZxB5CB4hXYvZZkkC6WIUFzZvOo9J5sd3psxI7
K7CvTobB/MJU1XCfrN86kE+qEqpNb65a/l0QgBUOI+uAms6JsnRjraxOZl42vDHTR/bEPyiw1VGZ
s4tquWI1dm2pSdguX/1qTAVC0TXg10g7P8v621EH7+XDJFIgsPvQN9PRRtaM7IepKD2NkRmXA0i/
gWaYXJ1XhVd2+XfYOo4tLblrog8zKflSGzodRo4xgRv/qUg6/WQbk1/oLUkY0SS04fLEuhnVy82o
4Ntmp+8YZfeoE9onVlS/G/iVM095VzxTfBt3VWr/hY2q+toDSjTHSVvWukpnAEwjz2nrOif/x3Uq
qDh+WklML4ZT+fjoWs1zXMvBEpVQ5BHodo5zjUj+gWxO6Dj/giozIbeeL58X5a1yrB86gpw6+Qh9
9rIdJbjhs5bN6AcJrNT4AXGghAvezGgQ/STFUV2tKovudUq4TUqtAAM9tl3v1Bo+dw74M0376KB7
UKoRxBUHuA8KfkzJfaTGynpGwzuZiSYKma3PMO/F1cd6PxLwio0Q6M6IAW8EvAO1vojB6BRRSF7/
oAaUsK/nR4WU4xXF2EDzNcd9hnP+f8bzzsQWMKaO+wlImFFRjkHwlVzk/xbnBQwwVaAjDsmjbw4w
bOurnlun7i/gUisv/rfRN1afOgsi+lWlIsK7Les9gbjf/fBlP/fWqaSblFcWSn/7JLoc7kzLfNjv
EwwTDUnEkqDZ1ukyKKqdRBQtU3eQT6SSz4OB+UOB9paH87BhD9qmbUl3TiAADfvFwoBQfwxi9SlK
R37RGpcju79NmrrjqkC6yDrewOyN21H/7Fx+W6+IBVGtJOScGRJZjXb+JABaLOu9soAr4A8y6KHe
/IZs6AbabSkJjgFAZj6BaXLm1XPyYq2/rBjBmGoOZnqZ+E8egVvmdMHqYNTotA45Azec7g5/ZtaD
c+84YiX84iClpRoLXSdgIGzzCOvLQ1ACKWfnfsRbF4al37pKidUN2IUt5z72d83LrKciq84B2dsq
1P298fWIq03Wdj2TijdwqY3J09UDAb+HPPPbbpHXIYa+Fz1Dq3av0udeROTBXWyTya6YyT/GTpSQ
EuzdINz+g0WY+/Beyoya5WNOs16Yotit06rLFqmIlUc7rWEahUI/n+9hsaBTRwdnFd3mRnKJr8Kk
XH1wxKh188nj+QCbK0VKrYASDFqPVCHqGGv60yDMIP/nXws8eAeu16Yfb6RSjUuF63HjQ6NIO7zO
JLMQtm1PUJB2Z8kN69v31MLp/IOxsg/SP0zOZR1xy3rm7mfVnx/W8DlhjajtxXwD5ponKvopbJa0
l3AYcQ2wYgr/XdrFnpy7zNnPIeLpfB7eIfLWIsxPEAHRrfHNa8lQY/s0EQB+fcNfrks2+RSKBJN6
ibSjitBEnxE8eQ6V9RyQ+8R4MRVWYxTqwx5JH5v1GVFkkxxgHQpl29+xQUtJRiiRr5QBMZdKP8/f
GyiNWQQR0+rt9x7s0xktX764F3DlWHzQ9ph6JjmkTLooFkUotS+ofFD+kqAtmpm+fEcoLblx+PCm
z9UhqdvWdA+zXWZnqT/7GygaASxZDUCKw0+2wrplsW7F6nmLdwFeuffdT+PZ8fZBDE8ZOeaEoszU
JvPY5LKb8aRimysvzre6yiPW9upUs/lkX3vXnVysDGiBVmRSBLU0LGAJycQ4uLQSwpHFo9Hnzgbc
/gPOtINbjPCvEiewibD3Oap8MmVJ4NAcVISeD+ujlzfrkIBw0boanGzxjRE4regWxti0omkVp4hI
CE87BGjBNEMWk3xGP6RJbQw8bQ8HHqufAsTeIN0Mw8gbNsoLjZnsYm3xSBPXDpiX34Wr3jr9Yz0z
2XE62urQhnw42Nha2DbRduZYLi+WmmlVVEjfVas7gauohfkIYOPBdT0V4ox2ix/tELKYgfA/ME0i
aGOsJpSn5OsVjS0K1x94oYBCljqAcAVnfXvyXSczKtQhFiNMNBXYqN5N1uLRLyoT8W82cUpHI3nu
GSgosIMsTGKWvHy7q36dfHsj+VR495meQiV5ltHFXqgF88r5TIb6wHS8DTY77pNny9hqxa5l3CeH
hzgiUpl2QNt96zlUQUhzq77KOX30lOx6XhUZIaXbh5fn4iE/4KKm9UUVOpBe+ZqqPWUGOmKl/7k2
933Ag8RYxq1Sb9phGXlhZF2PHdPTnT/pHKBYEvHUk5cihxInwn8mBNUk85TwVThdZNSJN/w0iFIn
QxOwgyyirhkgOFLPVJa6Z7kbqy93mxmOBVhS9/b68zW/7ClCmJFDjDpWVX136jtXeGSkKlT9njsR
4k6JM+jWu4wqEJPbmJNcgR1GhfJ6lJaq1q1ZitwC8S/FwSYbhDAfLuywS1tl8+MZfwCy76U/zryF
jdm3u4Smk61GK2YfWQURt0yuyID32YppGuC4Vi21K3ZrdVwEzAZ+8PptgoByVd+pQ/3Q5tFti0ar
H6SjyLgSYwIB0lQba0XbD2mCP0hce6IF5v2pkiNlMb3p1j+A4dEkHs0lTDVNAlhbJjuTBgOZx0qf
RvUaSEM8FZzED9ddsLlcnIQoKve/WgXnVZbOmevegn53m0COVjCj34Wsj70FYVsj8Lt4tNvHcUkB
FQ3iyslg/KSYrfZI8l/D6PUynJCmQ1wEcPMMpTw28QrZQ0r58LL8UEYfwIL/QQ48Hxa4Xo/XSxH1
0xksRm/2gOMcld9W+Y6SArEjkqB45id8TsbSH2RvpH2cW8ZeDefusArS7el1VvOLXlXO75c/f3p4
OALVh9otDRvI0BV8yyhJw5k5LXj8P6grQj3K1fQxc1WiQ8rx5sjsXfXlOsm3QsWhSZc+8u4sZdWF
ovee3Pk0xNUemzk30J4pjiRFgBowWf8hF+ROyHj/Xxit/C7I45ZfDXCYg5DFbCdDLURZEXNCx8Yr
FYd/q4ed3p1w4AH4Ngd+7OtFwpaewa6CuzVfHSlasAk89SR4QB6h8UENN8aOKgvJfYs27UGoUlZX
d410ViKSMrxiBq7zSIecMgHQgx6BGWS+UcgyOzrQK7P59D+Q/EJalkmdxawAmD6bVBL5rE84hE7R
UfhvbEe7yiohSJUxLTsiOHeeNjMWL/eCj8WaK0skPE7+ox4AaC9h1aUEgxasIuezeHoSofEIy9oM
oRgnTUbzauEpZsjK5sIOwNdnEZwnxbAWFKxA5GJAjS0+tgQnC9WYTbo7WQNTKm/D05l9vp9B9twX
WhPgl2EJJthh++i2DP62HMphpR5lEOe1OT0618tLwZDYs5hbT9X4uD9ffWKHtO/GuA4yCgqELNoN
D9WH0qQc1n58NSjqKQtb9rVmvvrxOSyTdL0QW048E7LnY65Ii5I38H1MMDhfTp3lcnZ9GCXvr5au
v1ODS7zVnZjr+mWG6jITGlFl+SzE2ZJCfRfk+BiSiYYN6kAMGM5uETGZQBdX91YtHj83/0Rqf75C
yyRPcYHMrzM/ixjQE8gvi2QWDcroCExN6xYOGwqRqqgghWD4VyVW1WWD8pDJShm1ijI8emYqUSIx
oSYFFlOrUHXN2+QMZjDn7vD8DZmusRlNIUjzkqv3dbSApYgFn1aCSW4otzCvQZkPeVrMHhkxkLXC
N76aj5URU1LN1KNFC4rI42gdHck5fpq8J1ZewzCmrMkvEOuc8Ax2pqAPoXtzHQCO9iePs/sfcTwY
C2ulpg3ICD027ww9zwwElReaZLrp5mDDCM0BEaNqSPLaAnQxkJEOW7pgo0ysBQvRrPIklAjSBP20
tGsO62KH5KdPRP0UooHHLxubf80xrmqOdVUn+HistlvfSW2YvPmtau+qX3EByMwjarJlGH7KlMIn
qK2MPAU8To2gchS4C6y+2tJC92E7c5c9uAqyL1ayoE/Ss2hPWLmRYPDCZB0gJYwfR2tdbkkDZST4
T7RW1PMXf3UczMpdc1RJwyAPLpB8FTR0Pn2lfhYQpy+5oqAWYAVLrimkZ58y2an31Z80DBkGhKS/
nmhHAaOUeHx5wkbmyw5I3pvHcY18bJQ+rqECGfyVjA0v9mxuW/BEFp5WY0+42l/5qmD4TOCxWwLG
cO9XzJJfdukh9VoSwzEUhBKnz3wVnnf6K5lssyx2kmC5Ya0MhETr+7DVJfD9x/OU8C/B9kcFe50k
7x387181IkWcUW9EUGW6WoHwcrQBwvsQZY3oJo/2YcFawo0KQ+zUz58GY5OwbpjUW5jvK1qHj+H8
1IhJgNC7bGz3iNdcwiHu/TWKjlDsy3r1GYUa+XLzTltc+6/p78k3/VIKKnk2lZenKnvf0SJiD2/9
wDiggksZad1sP+WhTk1lCILN6YX7Y5i7CDo1ra4j+LcfNgv3AlUhYJOqIykbAHlviwXJybTURasQ
BywaTz6Qz8RTDat52tu4LDl4oEY9WeBkJu5StMg6U5Q8i/dTs7umLFCn2xsbuofqz9UdR3ZEbC9+
xa6+E4zgTCSIh8Pjl6laahXchMEntx4SC2omAKuyPa2WxaESKxOcjwdhJe61Q6vquh+kERlpZoyK
f5xoKF9zAlhFrhIOLahpUryB8p1xAdRooV/kkcwdH7E25pR7UzcqPumYToERwjt2891QBQeifiKy
OdXRlMVcP3NzbeOLOr6K5d3DN0M0RmzK+xAl/+0i0i6T/GRqj5cUl/fd74r4WTAKMMQzJJisUbHu
DKYGgHUJY7zrCFkTxgzmckT9NYhXd1mYJHTHrVM+amTr0/0hJhrHYyX7rVu+qibmMytQLFTyz/wA
T2YT8etrHJi8CJw+g+4qDncmfWMx4NlQkZqPnPthNKyO2D8s/xoBQ4Ekgn1f/IhShXuOV4gcTs2v
yr3YCOrNeLdYf6KHJts1BSMiIYnwal5hFiX+2X+C58ER4V3hhHCN81YPGTRTjQG3GKYrxRpcCRl+
6yTV47IOBYKmNgukCDPH31WCEk+7sVsNbWekCPwgaUcyNQFQPOJYK3j8xOS954cTbX+tLs4MIl5g
DXl+cWVJXHxS7g78+wuOg1P6RKq+rVV40jTxHPb0SbjvF3t0wwFwmM8E1m5l/etq8In66hdEBhtw
shWcw9pwD9rOjqP5JA80Oiu5zvw3wMTSMqRTWdUjsd0a71CXClmxsYkqrEgFQkXJ2jRw8djaQkCc
Kqz1uJL3tXxUmRw2M/e2RNZSZ3aZCkKggaR6zss541A0IXvImB7WqOZslS0ZdzDmsTaSiohpM+n2
r8tShgz2+0l4hYUpUop7CeHSDZBtVmuNyIr9wC7Ai9x5X+4Nomwzw83d5JoGVUIXVPa7DvnGAHAx
Whl/dyh8wrbAb7EMiFj1plE3VzsL1hQ8Zr4NtY91tDQ205mQzgRDnQnM94h5GXQ5UhSdS5DhJGyu
+mXavivHM+X5ifQmeOrD0OcAe/81DQ3lvuom8DEQW1WIukvBe0r8YB0jo1xq8PiYqEpJTWnTjoxL
+G2KZMY4P6B+oQLQ11lQYkXGYf6oZ//O13q0jFCyQxDdSfff+bl2V+mCo+s4RrKsG6cOCnsgROCO
DF6Vca9x9iOeKZPuv9rz9wmILecBwuwYXkKEi/CSd83OmfCI6yHEjsWXxgDyr5/I92mq89laM22l
or4z+ORJgKTsfZZnW98hZ6iRZWlWmVu/5q1zw75KtjO07NitP4ioaz/j8x8YlI0FyDqQW2Pd3kzO
ZB944lkw1jOhZ+CHzqPQOHobYJ1TrsHakHR/qE8lOdckpN8nBo621c5yR5KQxIw38+hXrehnzX3b
bGY63bx5PXXkYCv9PE4ih/wBxHBS3pY/7g+IDyf+5bMCt9gyeDzye80XdxuQdNgoUTHBEQEb8hbm
V42ZJSg4Zwxu+ljq4wvwgsyUzKwo5g3McDUx8zZ8+nn29mfvYrhijRI1wvYaXw3mUFhy89G18dP8
/VkLAb5rMfYxk6xOpIgDmAyw3Puvt1n4kXImD3vkvgNl0UuxgDcS6eJoE4CyKJ0reTt+oP1VXvtA
vKW8gYV6+ulCftJsPTm6GAx+9nERisHQPf++/Qu+MAfN79kyYnI3Q3GElrXBVw1zGuCX4NAAnlfn
seVbDwsJC8iL+LjwAvRotzpZAHaMJ4qu8JWe9pJqRIAjetUAJTCpCIAqxC0eA9b30NKM/Xzyj34g
P9ELyHoYdtoVk2zjoi0yep1k/64HLCHS3zktz9Ww2r6tfA/HaH3OHgQCgBXJmIvja4GJ4dyUL+Bf
nNc678no4xvpcbDyetvIb+u1RkLxzBg20BLaSmuglZ6zLR3lqCjD/SnCozG1kGAqK8VR0134V0u8
QUDMCTcYBbaJ4amk8/1Zk1Gpe6xx6pWpe4Ej12OhQkfS9cWZXHdH2zT/yw5E/U9j/lvFVLYpsF4P
+0c8bsWYsdv68NScNYzAFpqcwkGfVC549HDj0zG7uDabeVzJ8NWymxcz7Av7YwFZfkBb/rWUyGsP
8eKWroIn+rK8QaogqW/gGZpYzpFpqxErMtf6wmVfnOJwyiTzHmMSdwBXsFAgWTt3yEkDFiyE+D/h
q0WK+BflwG/148vND4rYOOtMLxSk9wpiqFbLiuzC5Rsuj04TznaY3WWyuGXzT7+T2Exbh2cqtqcQ
UrCqN6Zn0Uq1Cc9+tqT5xX750CFv9zIl2ODGQc6ORtD/mzt8WwbAyE0mlFvHTMTN8MAM+g28dUTx
6dpBeb4ZDlZneADIDhrdirNu3vEKAcDfY2tITewHslSs5Mt0RlfpKfjfi5GIEgADa6gyOTTOvYhH
ySilVq5W4SHxthgeFnQr/xgDvQpk1LQeaj8CxrmYOx1H29cJBKbHUchrDz23fhgvomqt5Acpnqt2
CwqLm/GzR/ZKjOwzS8zj6d4gO3Th6XSXuOua9PLqTFnAHnjqBj7Cv1+dwKx/Yp7GTon7MubbpmSa
TzbjPCPFmyTLZxjXIfFgwdJmPo1Yj4agRHvMgCzF0/w+AttwvRxWKw6PnAa8RCrczClp7G/Juhn5
IDVIkhcF9UxozI0xMSXt4YnKu5Kq0m+E6apga5GaPp+WG0UFXdP8ft99fl6Fq3EGuWGcHAV05l1t
SNKoev4N6qp+8GTMb13m8TyRiRwE7UpOjcoYtlhPU4MDQ/5Q56kYe25hJpIu+qU9rB9EMzVTIqGl
v4+8B2+QeqNgjvZJDQfNjaGKcV9PAtEBCwNeLepdQUEmK7gRhJgDHu+UEU8bdXrSS2HeYJHLuQL1
htYDKlnolnk8x+YQO/2WaUBMYDNIeuMOBZwzbeUCPjrBN5q0Uh+0+hgoWLlmwyXsjuYPdh9uYmhd
JT/9eJWU6LU0gnMEpAorsx7WzsQlu8NTUOQ7Z2cP8DeFozuuimsXUb2SfLUd5jwFGxOnmcdNrTSG
3S3xEwe6eXVY4iqXpsiu40UG+6Pu8tAx/5zdmr8SlcWIQNeOZRFFPFJfqZo1BqFuE28/o/99E/Iv
d2HnP3sfGZ7HI/Y3eCV6N6IJ1DZDVi/8rYlYyR6cQumfrif26i7kNnGJFqOcLfpwljtGfIPCABeG
n+673rHcLAZpdde8/5i1RHZ4r5QhGl4WxtFv6Z94+Jm/YJin7nBhdsfgOmMkZHBjww/DX6XeDiUi
Nr2uP2qobR90Tmy5ReJsK/TITInuvvIq/bNstjyfZb1VrDn0yHEbIcQfuCjElyxeHmZrqZO+MBOq
66Itv8u1411JZbet1Kku4vMOKqTl5IqDLvsIPNxpZxtcIIKX41R56IHIcHQelhlC0vho4Z/Tzvro
8AZVnwFOYtoYZQN0fmJmWBWHi+vSd+nx+pYtPFvqpgfvDcOCB4G6lkuhJigVkbi9y1DkunRyGXYM
1X2X7MDJFHUYLI1Za3luCpjgd1bTqN4i9wT1B8im8PvNRn+2sdpiad43EDId6YGCg99lqd+62dW4
qzGWe5gmufkd34voMavhhxhsD1wqi2J3jhhx+rkUr5eSlqnq9m8AwnF4q8bSBs7lVZjuDM9vefHH
6xMbrqioVDqfHlIZmH+xSx2Sm5p7IgwEA+lxwp9o/2lBwmdTxXobkA3gWhkVs15KnBuGa+1zHugW
ysR3R05RinlHK6jrRYYupTAbbTPHqSo09N+KjfUr2nssph0ZAQSy0J1c0Txzi1xpsacAXUoSh2PK
2YZcOabpbUe4UbA4fko8LI6WDK7i2Uh2KY2C40eu8i6KZb7V89ED/wnNU0mtt0zwJfy0ApoEHtAe
mtl7JCrftVsflL8lFObwabroPjaStAWoDWsJHGGgQeq1AA6xr7nTpvtqTU2u8+9bGZ6F5sL6enG8
EBkFy371xVUsvatMUKPCKBLlUbpFyv2p+cRmlijLC+dxwymowkXUr7ryMzOKY0Sel+kfMvDXATvD
mkF9bwRET7Yo352ChNwt2Xn8gay1YJwZcUktgxZi02M1gCBapLaTBVQFaJAQPyHDK6vRs2HPF57f
YYzt/zgdKMAqqs7HBopXmZKNIPeveM6Jrd88ALE9oxs1pEYyGR8bjEUDSPv4FQJ+3HGvXjL+8bMj
xUT/NdSpB7xOFxTL3walr4vxBPOIKf7s8YnDMaU/iq4FFQvalJ/MnJ299UGFpwcoRpVhpgOSi6M0
Nba7obkiewVIlYh8qH9ahl9aZ2T1lrvfpldOfclVxrge5Ul1HkuU5y7H1Pl6IzOL3mCD/SYEX1ir
PcbVcG9M6AjcxGMw4T7swBJxVBfRngMBw3Mu949IdtqQ4lckETj4aOM7GCG9aatzvJe41letOs3S
lnHg75waZTWuhIgeMfDBhHhR2CZjnnLlQeABK/37eK9Utj9EJ0URY9HQ0fc06N01e5++BfdtAZYm
Uz1WuO80N83FrwqIVeL+qg9ICEkex0lwzOBrM6gcCLrxjLIWy7lOXvWbd9J+6u51MWivH2Lr2f27
cokMsf7Tk14Ce6tP2CAF+puxQsH3+3ZMTlIIaZnhwQ1lHYpPS5OFaOGeJ8YU5vxDCJl7k8BVs0V+
dhhT7P7X2St6jNIolqyQYV0DUP6GDWtzuXxAsukstg4EZzvHzO3m9/+eTX7lu9n/yc3tXgU6q/pW
PjwuSgDMuxM5cLTvqOlXVgJ3o7d8AwMxX81MSQDg28biGJVT9RrhZYk/FeKNNm1e+yvCnw6ILl/E
E3jyXdmJVNSsVYoarQ7Al+Y0pBt5+VZmBq1NHIidHJ8B1nXAF+hBHJc6JymuYlxLYt+OCSyFqGoy
lW5MFXD36lrRGvjJ+1mjH52CmeGMYgsMn/L9G7mWK0RZTRHh+ugFHVEtDbn/JAQVtdwwmljyjzTH
leuyUXPooeIU/FnSCoW49hVgOLOQrvjXsPWOIKmtL4YfornQHJoQ7o7Hn5t5YvqaHuo3anqG5uGH
QLz0SQMcsJmey9+cl4WScTgnQFFImJZ8tsRF1c6OKfTm5fm1Ijhl7eHz2rHGlAquYjVjgw6YV/rc
h7oyIk8UZdwyVcNcfJnBTw0ILfvBDWBducX/bHgAj5CfPghxricvUbAnYg4HPurnlOYi8X3GDEeM
Bm6mHl8BwnCIltUx71rjlPyF5PjRDVrxl1o5O3SEeJHDcR7I5ja7YOUx/rpObyBHjB1G+/KtELFP
M5gqH0hDsTVEj+2KLFEXM2GEcNkMocRJCzYvNcxIivqxJvVP0ZQAQT9KjrDFQW1gF+/6ssQHk95h
Dk4TVNw4J9lfWavkNJDJH8aAD2hD+68ZG721KJg3eWffyXtbbm4avGJQp+g4zw/p9U//aoQwr/EM
QoniFZNLEg09QzJSQNCg2m24u9Oet1svaszlLqaVF7y3eg9OvhK4ZKw+3ggJ6LcsSE90G8gyIWwG
G7MMjiV2vvzYTNGZehrSKFnHz4b6vyjX1H6wTkxZMFsKKSKMVQQBQyirxeseyUufInKxea/JpaLh
iEp97lYSxX5OOVcg0rzXJnhEUU4vjzP7ipZ38jImjUhBNWAJy7TFXC6HWJEFXue6mPCFe+SJmdai
tfclzNwIfmcSfQUdDvXXTGeFNmtZFn1zBQOVQ9qQRePSFXvpUBEnlamBHkO7IYB9UsztImLWCGCW
gGpO0c5DJ8A9kPtQrneHzzVMh8RZTUNDKSKmhW3qIydCeIfZJc2QQT656PsIII9fPiCbkAsUTIy9
GPk0cq9UyhdmvJHV+1TRt7vsw2XUJm140UqAR+Ml9Bw8gPl6dEiilyhEiag65jfvgEN73wi3+PGp
Jn/QM2qqeO7sMNjxbEwNm0QovUlBtXzGWt2U9OWWj/CRxTG39iml9rBtxjucnF4WEeI+nV8G4ADy
YWrLSJc6893VV12PV2cx+LN41lM6v7Lj7J7KWkmchHBmh86DWERVpntqp77vaLudEh8NYiXA3NbN
rP4pBNynLSFQCGdtDtB/gOdkmbm0O06QqOSu6j7GGVFGw/2sD8dGXypQ6UjOuJqVsHynzQUMa/56
7sC88XO7KKtGp7i05YDOg0DH8zRHlHTyRpKwNQm/MnFqPxlhFkzDAQ5xdAcfvaLGz5b9lNfXDwr7
S2Q1P+DvzhVN17FQe80FwSzmmFTeesM8n4BN6CUB4ll5LwJA6c3C2MEvnwjUTIxjUv2QuZQaHrwv
D9CNAmdH6/MtXf0UIyEgSaijanAdQhyj0Wd+hChwhF0QK+6YT0hNP6cVnhm7XZPEk353veCCmCuC
iNe5pXSe7xIs+Wxbjl3JGZ2fzFxYlVAnQjHVj8cKaLe9M9cosALyyVEb4J8BC286ZJYAX4pDG3wJ
qL9ib3psTJG+rZOW3nIIS+83xdLRIHiBvwN+oKqSJYNDj6/6VkgFgDHjlzlH2DTA//URUm1p+Bp8
tdv4LUXBe8YAp9Trbx7NhMPdVOcftmCFO/05VKaFVgiufVemuOelPhc+XZEsbBg3xozcDf6yqwFn
DGSoKFJo7ux7utASrkAajaQ8WAa808GGEnF0E8uC9SUoZoPLb4XCe9OsOLJANPyjNiGDcZLM890E
RQ0qok686DfnxrlNCyTtWo4sUiz9dKhJ8F1T5I2Yr9DTRFrtOJEKOR4O2Ft2pTDULrgNZw/1hsj0
9NF9ACTsASmUgosXGkaw9TeQEKqni9TtKlm5IqDtWVka4BCUuBG1DNB8q3ZBUZuIpybkru0irHUk
kMEVbge9lYh2PCX4OQyy3fZaADupIC7mq3ab2PpPra6uDpjySGPrENFNKYYfpwL4kBTv+c5EzgIF
vaHtbO22wAmT4Kz2yGFHd0dt/xzRZAIJK4BGFLDskvATo7jxILBFM2A61uMiW9K08JG27Q4NC9jX
QvCcq6YTuDjVBNe8jRne6HJjxIflYWk1TTImSC9m4ZKqgUfT0kLKrvAIQAyhlR+A1j0Y07X54Qk/
nXGBjrnJBI8dZglIUBh3ww6kWs9rMRFgxHMpJgafqYheWDz5CHe3PZ2gSyVep9eTAH0E9S/4g8F8
Bk7aecAz1+f77e/GN8UaoAR9kBg0FNa1YJ6JrSiTPGlRXC6g4ZdyMdTUG44kg0S8ZfuvuX+o9nqB
WO92/81B4EvTUagqtknG2CF4/GM+KAb88onI5LS/oKFdvzKV2meh6NXU4JuyRAu7YkDpAcZX0+Cg
6KunW4JBjKoYB5OBJKUBx3KlGEA5Euzcs1O1NYzFqG7t3eqvzNF0HGkWGzzLm05xcyY5RJoaYuQ7
7UyD51tXqbXuUlUkIYv0bYdrgA3jZf1d7J+8JeIzS2cNgaG6Sbonm3aLQ2uNkq31kMWsHkDaEdOf
GAJx3VSDGXbH168SGqLSlP6IUs1ipdkjxZqid/A2urIgRvQLR16W3/RMcugv0MSIJYQBN0k5gx6G
RlklnORKKBTIMQwWYahMB6Mbv7I3NkE0GWPEqiwwsedg8nGBd4B0FtUHs4bSO0pPZpMiEb44nR8o
J6Ft34OBNQ8pvh/hPWwWN/bJodmDNYvHT+juqLwBs3RzBKO1DpEd5jLJ+gihg0fNdG3m/euTT0Jq
eAX/9Ui5tFcM+Jj3evUOUClVivSVWIQXxZHCoRjrkJoTK7Dybie2OqFsECo6+iKxc7wH6R0/Plle
jIC95/1Ads5yZujKZIbheFlZd3fqbxgXWAS3dcpg/veLZd/mQaqMSb0PWM8p9EjQzB3dlpvcA/wF
QKJSx/RDBiEO+OdwmSHE5OR1cvpxhIgtK22PNDOgJeeLh6HmKhpvjYZjtYQhNk2JEzliOb+MIwHY
7nSVWahAhAUHOHL/B+Bvm+a6iKA296uwDC5hWD7QZUzUqy9m6gO+1fQToDXP7vedylYrbm1XfJaW
dp98cF21SLlojPDGbbMWGbaDrh9uOHXFksS9/rVaQBFQf/HFTrqnljTyOT4HimPMGyXdsynol/C9
/rYc/d1BERonqyzgjsDW/XEnKCJ7pPNVcH5UDmrNQXJ5R/0flbPDssF0uKl7czqLVZoxMdbOe2ql
ws6wT5W6uu9ACgCO/nu/u9fbF/LhFmQLjGjvBes2TYgcM6x3vPWFJHQ4OJhycPBJvkoNG8GO755P
LyizLWkl4wPSVFAAhvt1i+2n4Q+NrHDvajCmrgwsr5AmSFlEyygJQgE268cIts/lGGN1pIgpdRhQ
OwUTUQVCbHv+3zC7MfFayxxanYwiOTjhG59cRhlDNfLOPrGIex6pkhZ9o4o05xeNPWGxSwm0STSx
r+Jk3p4lHo67eY6iKNbNRwhcIuzv/kIdsaiNPmT27mBmMsu7Z2QjJGVx2gI3piV7R7VdPjHmNUah
+5EmYtKP1S4aanaYiJoUJLNLNoga1qO+2IWWClQtvDKZBOAbM93wGZJeO+AX4TCRahscvVLsP8pr
XW7aXD3LO3+m0ttRMtaSDjiGLN4FwKRLOnMaDbnTIJWauH+9lNDt4nK7zH045kEd6kO38svaN3VH
Yj6xkfSnPHBjnLY222Z5uvH7z/hrd3OKrfFcbBwj6TInbVVgDmqD+pXKaaM5wgAX/Lh+QHmV0lad
2SVE9am8QqZ1Ffmom90/1p1jvhJolqyvcC9fO5cq/P//x9bweMwQSPxRV+d64B5Apht8Qx+MrIz8
6Wgl8itRSRvF7OzDMYOybgj4ZbG0bMoY9VrQZGLL5EOHuSxTJfh/763ewcZm9GFWXHU4wWHgFaNk
Wylt4edwkeERgDeqxI2EcIhYlBqH+QgaV6KefJfOQUsU/C0KZ7sJf9LykvXjYl/Q48AEK2hSLDpx
lJpPqKoqfGr44F3phpOU1EAdp+XSJW6ccnNxIIaovnOql4V7/UBWiKzUAkkfL1pIXxmPPJOH8eel
5bi7yO7uOs+K/CTEhFIzKt3fSEpfrvvDQAN0ydC5R7WMrRhnCau+xP84mr3Dzd3g5n8rD629uFtu
c+KQRD8IQ0Dakr8xpf7hLuZZK4pn5gcuy44/BQzrS7lpKhZGvdQWt+WnEqPzXJyv3LKT4UYyN0M2
LDANYMVcNFgTfTa3T8okKVhhepQ+L2YqAR6tD/eEfl/0CqGGUC9P7S5es9MM64QSgP0Sjeclj+tv
z+n1ozVjeS25gi3P4cL8JZl3cdreR02nOSkVezM5O+3EvwsuqFTuW6SXLN3Z4LfD/2PIkW/ZbAiz
9h0WY9VoUilVpuHMNaM6SJLeoDnBK6wTSuaDmtd+WPAg1QcIeoWlw8vAqQMlTvFChh2ExbRVeAub
sQ72kOPl0lILC40Sg9e/NsKG3qNbyToV3raNowAmKe99KYdTkgjo99aBqwNWsqZOrjm68R7aDt+C
GCyRAGz0RyXeNrMd0/GfMy+H3kKpzg3g/YZJsMQuFBAygUsXNj8q4ajCgbLry0v1WfB8KA930oiu
7gFhaZG3YoZBCrwYlQsXudRSKUEnp3G13gtRnktcxKKbwrteELLHS0QY9BA4Vuq6Z7C3QIKETH5g
KFfXB6/sF71jeLRAFM5P3KXc8IGTarmwX81Vov80Z8SfgTxytlC1riGnUPArSyEE34T2JUwEKd4J
reRILMX8+N+ZpKpBqRpIJ+yvq6In4kHPdhUnpCxSfHUfGhxMKqrx/iUo/VcdOsGqP1qwKYNfyOJa
BQkVRBTxLG7sH+gbng4MKOceW4TnbrDFvoJErf7Wgeg2iqprGf2hCd41LEr1cdxZweZSgy5zaKVN
0irrSag+WeOiwOd1LCyU3MVsb3WkSZWBlaBvd2z9+aTsN9gaIV8ujgnLdOVKKCGBS9PuIqWskqSR
hzhSPlygZ1wmbrfE4qYsF8y5GFbOPdbTv0K/Ovf//lqm8UGKcxaEm8IDir7COV8m+c7Crmr5w0ba
hQyZlkmYbl7HcRwOH0sU44YlfG3yrNmLJJe1Fjx+2LyRXCJwFPSpha3tB4VwBIimLbre8bctjoIB
0c7QG6+2gjXJ4O7+KLplakLG6tZ8cfOOK+6EtV+9sv+VbkXuvw7F54Xq7vtvN2vU8+GTW7eHVjl/
QO0z7RnqleoIgROigqcJig+ukIym7EIoaD4nUIwazp9Qv+4iDQ/wHIsHAbyIPNel21Cxynmdgaxi
uSuys6FTf7x5QJ0csqKRc3i0klif5ELhQoxEoiPiC3PD+gHw6X/2Sywl2Dhq/nXdYF+Kt84KJPi2
Xb3nzspOJwe8bBwjI2fM3vLStIyu8rLXAqBhNSbNX9kCACJ3D/cliLQPorI+LGlo81CzkarGVGQA
ZAljhmJvXzxPhbOCexarHgHS6NoQb4lDI773zhdGO7wE5nBCdAYemu3PrKFTaV17HS//EDhD2vH/
gD7DGxYeLmcD+fmZF5gylepA7VGFsddIflQ6RqmGJ+x6cDPdsT9Fh6Sl9yNzu9X025ArdGnRlA3N
rOHmg6WxglRUPKITsM5YQoij/qChuC/+Dqxc6m1FuYlRKDxQJDsS2ARsiNrj+qyDXwbuF2D1Wk/n
GcDt7LKwfh/oiVNMVQOtWqDIUQsPzg0dlvb9Z46W3m/tACTelebUC4odrJNHpD0FOMJB6JdlTgZl
BmPF1G+Ry8TxNC/bHCw9dE82HhR3a4DX55u9BrDLMCXd/CXcPLpAihswiSAYIuqg/ZKhV+4lbvIX
oNMxloZBLNIs422K11FklDtkysU2KlS507NVzhbDDK6J5w6afRagnj6lCp2f6cXm9hzmiqRxdkUT
qGXpExPaeLTiQu1+8y93gh27jZTpG7ckBQqh9rmCrLMSur8Mq7ZUvdFFa+gS/8jDkqzYJCoyqIKg
P9RdIFZ3vNgVT4W48Tn4ua+59Gy+WHpGJvK+QRDNMAKfdXbCDAUxuy3EQJLeXnKxPPqHI+7TMvt6
RKO+wsLsn5T6WyKFj+ETTdleaok0kPn1pLnTHIbiyt7J68ITNq4ojk9BfFQlQhaL6nOzcZIn7XJz
qsA9LSwdN3L/bvQuemBDAXeDdLG9O2ZJF9ktkDoMZkV8Y/trgGhREmt3bKCJjRa9ZNE86mp2sEek
g2ajreVO7yAt+uSXn44h6WYjE4Qoc56P7KVMMNrQHJN6Dmhq2ELZZ4wmC0QPRdBL+XBcRl44J6pF
YhEVHWpQIaciAp+wJeqQf8Fdl4n+sbaeiYtFAC/Jc8FPEabuXMmkKDj1daOvn95B+C8WM8lvM6kR
Rdr+Q9IwK6FOBNTKKiIATbCsWsJYzcVOEr0VTBkO5Mlyqdfn+lSguBCyCRKU2c0wS+BVwK0Si3LV
/ysUTBf68L7FTnFtrAnZqQDNB5zvsxZgs6F/cAiR+1kI+KmJoWgXXb+CZ1IBLPg0oUJVLINXIvp2
aSo6sYpNirEY010MEEL86Sm9rQgrJmoaUc2EWPlq7z7ZV4YMezvErNZQP+DYTPVvk85rvrUgeCpM
q5K/KOilnJOgS7Kyvobf2oIES3WSffvD61BU7dG4CjdVzqB5FKFIPQYQvdlkRopJS15m4mTjWorJ
qjyZFsN2gM7SDqgK38oX9GWL2fKKR06h1ihYTgeryslc1J4to3l2Vk7LL/TfF18a8jfKuF80Z2Tj
k32oZANLFD/B8WAAGPYFtXmdNOWqqYNRMdP+G4ubCLNZSdVQwF9izOFHn2pnRbtKEyAUzJj7GL3T
z91dWiwSxzSXU4grUa5rHguVD4Aq+Dbch+EH3oV/fOBDpFjkNFdE308Il2K5fRtwdrC1DqBMaB8e
7YXodsOtyeH1WRQpWrgWInv1+T4THdcN9SwU/p3RyXIFboZNKP2/utL3AkM8EYXnlxrdD4D1QyhP
tFUqKpXqwbI3A4Al/Lvmj9S1vqU6yXTiXruK4dkDJA98jUdzLAWmWVBlI03afHVBLOdyLaRMP7BI
N7caomn0yUygNXDqMcyOJTwJZtsTTSCWOx/DeZud99VCaozflDo2EFLyMry1wuzG1TmE3z/Nhl8s
tejeVszZ77o0VEdbSl/IdOOMrCPed/gsfB3yhHDd9i32BuR8wILvwtrbaKGxcDjqyCBc4ZPr9jwJ
Wh3ePs5Vg4B1rWxLkaXCAU5Qu59wUxw/hIoE1km1H2u9uX7Dhw17/Ld2izrCKLXNy0BMjmLeoyKq
Xfr3Ftgj12uMv3ehSLV5zYOWCBSguqIwxFiJwXNnq79iVaqwtdHqXB6ZrfQJud1w3OHDGOiiYYBu
5Leq/pnoBb4MqS1pE3IxvNtJiLiiXjefxGQ3qF/V1uPFyKwzeXrAWiCEI1sD/VtO1oAuzgc+tiI6
aU6oCGJkBlt5gGB4hNIQSVoJNCAA7cVVJIAGv7OYw0v4HZAfYUo/VKLfhDmHpCabC/krzY9uta3W
yvosFIVA5nNtjHQTRyVpa8x7L1xWf6LT/+vuxjvYmhjxEf79kOvXRYfeB0iyusHzN+iGBVIiaZFs
SCC9mGGM+BBRsPC05PU4THcUJz2btd+uva4TL+/XAW3duPD+0meYR9L4txMWhRDDOu+RYrjMC0yS
mLwkGvVJMUG6GAyRk3LR0dRDApnKqJvxclyNq2TylplBnlLDcLWp85iE0WkpKG7iK40VYoqQXmD6
vm+iiU6YHu6sbU0l71ZYm1xo8L3k908lr5i+4xG2JEuihuwzYlVpFa88eJKd8VRBqtLG2QsAAMGl
fhgsS8V19NY+tno1qMwhC8Yfzcv3czKNUShyKDdZkFpDNIke2/XP92d0EEEXqJVDPLWQo9siv8ra
3S840R139twqqc50VhVl55+hppLEhV8euL1PjzZzDDgSe1pwDZreLA4s7CT5q2Z3mN83jT8lmchR
8m5gpPt46z6b2mkUu73HuiIYDAwMVyoUZm9VqNuV2MJnUvox/ZfhyzbzAWBLpE0DdvvE5qVGk8K+
CERGnXO4x3z04XUF2TU6BoG28XyoIL0p5Rg84jQlMtVTZsCDke/tBvMd2KPEuiE2xNUvrO85RjQF
LM/h/HBXpvSNfr9BrnPJpDaf2SEL/JrSDswCshHMWzSBz19/khtDf+e/3p3d6W0XharxQmEieUln
pSmdfVqMDWmnCG83yVpZ/+JOKdKNcCcUYcKu/qCqIbBZSLwuufADb6wp20fa+I7nqa0k80wjlgGA
S6N3/6CfvQ4OjQ/IIGSw1ybQssKJjTkmR9FzeTALezfx6Z9s032QJcaKd9D096KGPm6MJeszDv/E
J6GKm/nPWu1h2CcTX/egccD61G3vo+5nXJFcweQiMBEcSG46KcQvNNPOBIylU+nn8PNCan7CZNdl
cQCrT/vDtAFQCnu8y7noOVJstEXzfNTDl8GCEivYuZwdJK1Dn7plR3VZVhrwzMJYUlG3VRtluFUa
K1lFuBSK3wCHsK18s27+CTNgScdRL0VqvxFstS1/4UWw3qQRw00xWGhbCc2a11WxMVdwWTuIx0Bn
dZi8KW+0rS3dAOipi4Ih35NWgL1n79P2LRNcRQEInFOVIr9iMkc/E58peYzDsI1DBMV+7WgfCF2u
w7Fbemu8Nnt0jXi665Y5DiY60J6/NpwhoDZmEpTF08vwxcz8uY3zvk4TQieobfYbiouynJoKjqxt
a40NawJ6Yg966TycTo4sYt1NpSUOQw01asvch3wyzBYKB1KQenMEMr9R6GeOLkZnsafGsssmMPto
6akjm+fNf9r8hQRvwoWtivSUIY/gowq6ehytd96et+X5S8WVkQ0LLp4jSTUBoLo3Ux6nEHMj3Wb/
/l4U2/J3Q400d1EIssOHLOi5YCkrtY7R3tkLUd7fpynMlQIS0id0U4h+3QFHWodHZHgqCxQA/Kx0
7+zP3tew+NrhtuRIZ7XHP5Tri38EhmQuaFeFu3moevykvEY146LfPKUqE1pAw7djaqO5ixdtICOl
6GptJZqAgtWwHUCL9dD6ILiJq0QG4a7b74835oHNrss5mMgw1ZWb7eBxWJn5bfA+hs+cbIeAAOpj
tGZ1nMZqgE183PL4Fk4Ds2rPYYC8g+N52C138uoS85dMF2NaOyCFMUaOYCkga2eP8GxAYhvyAtIX
G0GSH33+sbfWp/7hfbJNfo+J5Yp561llNETq8fDMTq0+ImchdTjVv19C0w/zXTnqSq1cvhvb9YTu
TXEvsqHLpyB7EotIcokQdhhNCAf9Fta1CNy8uKNswOkW7cpcHLA5idEA+22STuXxc7zhKMvz/BpS
K9jitrPDgY1MqbuYifD2USOOUWa8zGAal0gaqioHVx+7LgyITy+QVDe4m1LD9TXfJQT5WQgauShC
xk26QfmdIBBfASMxq+q9i+5AxixRQhwDRQVwzONakJpEuYfOlj6KIVeKE3pRSCNrZ9tr1GyDfJvh
btnu3Jd/BDuDsvZOyY7w6lGqEj6m75bSWlfOEaPkTxt5h3VX5g47z75crZUv22RyuKo+ha/4JM52
HCJpebt4NXI3o7x1B1oZiAD0mDaWUOkA8x9peV9mnjpo3sdKj1ZDSUpOfHhrfcIiHu9ich/68Tgs
tDS0XS95MRCXxyIaVKTAFspYnQfKZ9K0ism3xVcKqU/sQUDFX9leD918M3rrQniEiM9eeSLjozQo
seRAfA12BA4sbhoSMgktu4qq0v+CK57FuOJefHKUYz64dkQGhthEUhA8wSCRn2twGR7n/6jBLv2m
7iUuTRM9uWDbApKHDKpdrLrNPvNE6hKCNJkyktosb/YLzLEFmeJeewiFSUdptlo86xIwmTCi+V+i
zzpHn22UeVOdqMm4s+p6k2ZGk+JigpZxNrf1BN0N5rXg/Nq/ha8Nxl0/meuv5bOck8/gxTCaZCo3
yUfZjCiJk6G5JPHjKo2K0I/GmaqpzpcsxOJXm15ZLQMDsa10HbYRT06ZXYazPI6VkItwS73lqJ73
KH0ioDQM6Jw1pKTe3el0aW8DUmTu+tHR3WvmoDTyZKV3BGfCPHLCIF1HQIlzgBZj+p8MO22Ptsj5
H9toh4jtnmnIvt2jHyZgxyISYdjpRTm9O3LvzP44wsG96L9ELuOMARKJDIRQImbFkmk5E1+dyg1h
Wb2fbzStDKESJSnicFZdA91QVQ9Cdg0Ua71bK3vwnaFsBw3FwPX+Tye224g3eFHDf8UztGHq1oI5
KcBfBvlCwbxdaZtzFhcfKfc2zWBLgNxfbRt9/ixNH55byq2HoxaKmg91eXqHCLOut5lDNFafRG6p
0iVuEWGgeHpjZQ6ART30ni8zai15RgATQvOkjwsSmRPH2KYWVZbd/yOCWIv9PC+VoESY/qmOvE4J
pbdrautnlh73YMv+0wPINzGmamEX6FZjrS/ORBGcHn27+m5L089aVvuibRmc8hqQLdLgXA5kPv9x
XyoPscF91faUp5rHeIdFM2Okf0Syd+jTV+j2q3YU6MFEbcnihRanXRlSpR0YB7wYSK+YVUXuMGND
nXWZkpzeLeeuSCkBIkoPUQlYvC1LDc3JNhbPMsh+8yqzVcGrckUBuKy10PeevLvY1UC01cBfYT89
iQLXJVrLNgbPVcy8n2IYWlRUyxb65rWd34NIx3DeMEa1ajBmW7FyTUz5ZA1worhpBYtkfp9Jnq9h
UpWA3V+WuQQpyDOqKLyFD7L9/B2u8mRjUvnB133nRAlz15obfavZN0fs4YFwCnYi6aHsDErIwLz3
oh8HSSaDe166TQ5mtA2knyzu3CNOg8mWKbsukCK/WCnW+DNnYIC77HGdOMllFCf9BT1ZTV/m5iA5
ZEz556K6bhwjai6VJTZf8NdtCiKMYGwJwotMPWX4eFtCEHT6D4fMjP/2aAfdoGy6/E50FqVAKlR+
2tiO2tDthOUFTdwPEgs5cjGB5B84MlNY6QZ3D2AZtZtPKOCFfEDwZQswzUEPAPT8XU4xPwhryUoL
LOoJSREHk5rFOIHoBVy2Tl/434E2XB9GtEfgbs+iWmSIDUK6zxdrN+VcV5GKgGmLu3eKbucQXaHM
ByxRajltnAZuAoWqKh18DSJO5iCgHE/cXhfBq/6AOaxNO3m2Q6EPdI53xwh47HgtpUoW6zKBsNHU
tsFPDMp8PF4Xhsi7GSEVF98Le+mwdnRT9dafJwIDcl5Ut32zoiywT7rW0BHJzTX7ozPLUZk1iQbU
eIuJHBAEhPmQOIa7oFm8g8VzVziJqtRSrummobw/CtWsosQdkc3TDSA7TlnIVxEsSVZ8LEjGTKmC
ZaqQBY1ZMAN7QZbzg5wM2PcpbdeUW0zIGIerVP/HP3IjVCQfOpjj12z0TIvbeDpZMQ6Lin+l+/zK
08qUvswLuK5+QEqwTs2YGILMwETLMgE/LjbSGjYeq/DQCgJ6L/ZxlKKWpd+hhNewQojC98/4SPoo
/1nbF09CW8cGbF8/HNmFK5C8SvlXe8FT21wXfnRuzU/f/WtXWOcrOm0AgPhX3U/hzmzWtKbDE/8d
qiR7rOpdVFeJGMMeQ612aWWUK0t7CscOVO2+o+6XUtqnDgewWrUJIreE/OrHddwMdEbeBE+kD5zC
po93Obe7GjCxvFY5D/Hf2uTitNShploxq+CpINj2Z1HKPnEmkSfd6XYDUNeUNyieFVbAvZ7ST76u
m3LnLBkemvTaqYv+5mIv+f8QNGzLZGUYZXqLoXvq0n7jNd+UIAqJ+tCddjes+XTyh0ajgSbWF44u
EQR+tilv6JUyoriOLbj6ogZQxGxZAUzeniVXST2v86cJSWEhXa7F6AnUokwXwY83/abT7j3JC28K
Jl+SyLgv9VlrllD46i0znMWwkD2jxYs06+qJvurBx54i53/ytKq0JZV3hBhcid1EqRMcaXMjTXJv
v353TxdGFSp1kPdXLn203KtrNK6jodfQyyDR5Zr99IA2WAL/wKHCOAEb3qRPp6d8Io8dfhDjKI6z
qWfghKgUpPpwLx4EHQvJNaG/z5fJcQMtpcbUsb5ksDxKvhPSkFwmWc/dXga/woiKoY6bxM/gF9iJ
AAyV0N7vxYg2ebU92t2Tf6VgaQQ6vj/FRfnkgRpDItdL4r4MjhregTQ3SpiBV+5xveA2yl8Glp1N
IhAqVyPxORMAp+UWGLjC5wjsosQWo1+ljvoZ7jGciB0cTxVLSU+5BZ9gcIgeKWn55d3gIRErDzPk
bv1JeX2cAGfWIn+ririuirHrZcHA1GJ1OZtKJpJsDKYgfrzLRLfsymGofS9lhaW75+KRMuqz2Ua/
wuNwJhux/bT25L2bS3x6gxeDNtwDuQbwXN/3D1cOpHjwr9BrQiRGL9Ivw6NT25BKXzIBIXN6eo1r
1ClGCtTs8AH4GQpTC0AsiGPtgadR/oL3s/nKb8Rm1CIzKLbmZKHWqkYGBwX6UaJhh6gO9xAwq1No
3OoyOR7bzXSM4/ZunhxNQc49SZMbNMFngwkemUJdDrEYJK40RDkM0Twy6jyR53NVcKYUMFwTYlae
5K4gtf5mF8NQ75gbMViB19Bgj/jmVfWqxSrVz5che08rO99ZHdmVkxsdKFWSv5l//uPe0JFE7svS
I6Y188GCA3bgzd77kLUnsRWCUY3wTxEHuVDgKKQDbjtOYFoThSmb42h5Cu7u+yXl9tDORia8/bFV
yNDNDU5XrOhhL5K0/pc50ZtETlcWX0a/e96vaJlhUPkLRgsfQtj/0p3Obl3U/QKe46x+2pEQ7K4z
OTeDUCpQb36V7UsSmLkrhUxz+NDg5gx8Hp5CieA8L5lcvWMLALPxL9acCeEri0Km97SAJ51eACep
2L91VIy8Lt3GlIFPQTWqsZaQa8TgemT+AwcHq+WXLrDl2PmdJkrZAqkQUb65TJ6v3TzCMKFoVU/r
jJzS0W6q9dHX7f2T5hJZ8OWCXbAfL5mkP8mTmYMnbFU2zsnHp/D3kLNcQLdac8Q5cyeRzkABHUgO
9BFMafLfsBom+N61ucfIvU1dR4Ly4kxqbqlMApbymaMczHIIDBEdMrfUphKFvyrHQKVSCLsTOC68
lWtRG9+X+6CJA5FKRAZVGt3vUbxeGwP9G03liHntvVicflMUOuydIFl+gwb1oaGYWsudWNaf4jel
q45Au+zB2zWHxPvinCiPvQcDkNOGNIxidD1tRXnRwjM8qBeyakc09aaADW9W4vLDcEJFGEqZYUYK
f9YlOnPGk6AOezv+Uxnhto1zV2hRy3gidu74CBlqpOlDJYkfXZAkP2r1xLRra3dukL+hh/zPytX4
cwPGcK2bNRrvkOPX2t2Y5pEL9K7+GO5I5cfSjbPLaHtvbFuzeWQh7tdOU0etDp7rUu7WrXJt3gC3
6IRmfLDm/MIyI86AfAJk90l7HW0CxzvhsUOZ4kgtbKmqB9JYDwDvLhXqxP/SLtGlGgsZnmrifMZt
BFoww28E8ZhVtzW6THA3q0aFGxgq8GGUmViqrMjDva+R+Z8qsBhDVtxULw7JRidD8irykqVz0j43
P3boLSwbQ1SeaiO6PeEcyDTja4hBvLGcnKusWR/ABPdW5xuQAuF327+iBZc/qVrtp/jWPwNyHCc7
4wCKWSYhwjc3px3UkzUeA8+kHlbNwLCr7x2kzaBs+Od0USCFB613WFmSAyTLx1SFz//zL08LY0zl
3PgDJ8SwlYaFpCJGoFqFPzJ9o1e1nYX4RF+a5UA85R3OXrZssmJAd8EsNNPvM758gkeQ3lfy0Pfx
1RbofsKEJrxRcFdLCXdkbk/k8Fa85DXd0h8riYkQeOSjP9/llrEoD6PywqKBiRlw6gid6d1+1I8s
FGUkkIypFCcGOaZFa0nk7+XfBqAeFBtpBLVCzptN1WWv+Orefhoq3guoqVuYEggJAAbdhUvXIaYt
OniNWyU4R8lbbUYxWJ48w8iyl0M88cTaYlCeLJmJ1qdmT9VpXH3NamIR5LZPN758c99+5Sa64kQN
PvKc9zZ8I4z3il+pW/iDXKpi6yor8aBxvBAhC/E49tVEcCXcip8rp+fIjOTIGH6HUzEocYIddOHA
k6tdsEPqv3z56mdts2kAZleAvzvno/biycqQ/maWCXYgWSVzcoS8wb7HdLxQ+1gGmcJPhLx8zOOi
sokFd9pdyz9ezHf/4XpPUTQS/I81LICoZRYErQRaCwFkzkSp6M3Psuy+qFhqcnWGNxOChlw/ZT6H
FIdrre8KGt0MULspiV9P9cJ/TkczmcqgCYi38suZBM5Jd4/Tm3ouiRIqC60n0rk6h5tFBp0ViZ+h
rc1dMis6u4XPmt+ypBvPycg7O9RchPkyxXoYXleuKtr7Ws2nt5mXzWNx1f9gm2Y1F8StyyATrUAG
Yyki2nTpg9h6/KnOB0eMit3NWNFFxL1hF9zZLPOsMPnJdNsWovsSkRZfwZWaC2Bew0AmuD+klBgp
+iur6pR6UGHQHWoD9fAajCyi6mBYeQsdYHzCUYzpxvnDPgn83dPLJk73xCVRm9tF+4JjwYUg233G
6aou03dPO3q7cRy1yEHRj9mbrnK3HPcE3n+wsAr0mKz/k6ivohX3zh8jP3PMYjkT0VvccILnE1wz
4LgwgEK0ZO5AuUGkDt4cTr5mk/5l6QT1C5ctAdY9rEKgVnZhNxew2NgnoNjufjejr6oW2PWPfIlZ
TAZhNKnMLKz1cVfC+XK5c+DprCBatvHQ+Vpul0rh8WrgfPS6Strf+TvMJv6bC1cIwOSUaFPvzCDX
GVIBnrAxYvZf95W+H32DWj77au6b+8K8gOXs1dm3rbqqj1R7k7FtCbTRe4ekhQt6R/YbMVJGpZaP
2rSB2ExmzSHHnVMMxfWB8qAFb3IeP3PXIFMrg/MBUDLb/cgFcZEIQkvy0092sW2e4FpTJ3iQEE1E
EI+9GINJRfmyZcDZMvy3czXgXhRoN4DJdPM0xsJUbiqQPM1DeyX+OvfWqz9MV5DekHV7guxiLcuy
avj6YV5MWks3RFJ0bZbLPwdAi6IlGTQoQVxz8dXs1pu+Sgyx4j4qaPhZ6XYevSvGcOdklmyPruEL
PfCKBYUEV18W4QtJa2bNrhJm8eBJxJUEgcHanYZx79IjIw3VfSudn6j7JSuox4Xv6n71EpdYLzA/
pg8FoDPGUfif6OPk8pup2WWpnkDWQnZ1IJ3lXHLG+7PtMWigwUfHyMtZ4tKZfPjd8oNkOknwTwKH
fxnQUWEHQ+vP0J7ncXkmZCSHd68X8RPqpYuNtpRGKsXez35kR3JRTRe/COXCedmO+8PvwaSClxO5
9kKEEHjPt17Fnx4syNtQ1GDkELlMIAAhsV0KsctpSftdyGw0QVKKWrnZPjag/BSIGw5TUQN2GlP5
c5ztJAFKsZHBYAqDpNk01LyR5blrOj713c85plyXaGbd0NzLJQ8IbzCdQ+QgmrpF2BtTp724r8h2
3jeUF7M26XNQ11ZlsA8uINvou1hu+e9DtczgJoO78WWF0S4bydGgC7ZD7uGCgz6+7yyYUAVafx1H
Zw1quBC500XiWYF648POaw8FnR8+M5LzsyKfWd23Uui4j/j0lY7f5LS3ZnbzSQj/ghq9lrMdkktO
CPgBD6FQU1tleB4Y2GlW3kV2wV6TBmvHYMswOPPgmFU7Fgch58cSXSGatMpdYDtT/gZ6H2H5lLKs
2EMww1fant0kpWQ26D64TpbUzvXbMErDYaj/pNd6ZIAWWnXEWfhZR83p3Vz4qhRVomHgNn4mKplQ
uGyM99v6OjihIFSTMOV79EwU3hFazAuU5fE4FfNqqfH6kdE6EHE/5G4xGzbYOTGigmhmGcmaFq5x
VExoEDTFslF3/yDjDWVHmQiyB76vnhqcq5hG6PJsdmt0guc9fk0cYi/6bQEx0kTFIGarsj2bJGmf
wmOf2fvIn5NiPVoz7pQ/j+4DNDRCooIfIDiRXezSoBZeQE091H2dUtL/OFwYRTh06r30iKKJm6UM
0QUQjXP8Sd3Hh8Rp6wwyVbicZnvZi/7leuKsRfdtzU44ZgzXEvLa7/wcqaDLwWO9GjHwXifMzsyK
gkGdeggSSSe3dZsYWWAgTJ84oVEb6hwD9jgZEpNJa0TFMC2jVI8bTHk0CL1Pc9eGUROHe4h0le59
KlFXGAy4aBkjvQFSkx2RPsjAsS6ZUiwyKIbtMKcz61FD/Iu2KxGGn28mge89Iu5/8ahyp3u3c09/
On8o0aEb9c+VpJUysSk9AN6BC2pFML0TIWOqGDOAY5QJI48+eLsX0wzjqKqCSag/danaMUBzXwKa
o577KK7kIUwTbjv52neOJGmcV7/nLmDOsAimNT2kGgegPxQxJRLIxwhz7KIjsjr3OObCYIAA9gRr
2eVvQ2LeQbyLBWyYZq9CWB/GrpRa9W4l8JVcaxcNL4/oDXazBinfabvvQQydl3c4PvIrh62RtKdY
dt235Ym/FJHSalVJOOZBvIczIkdU2NTdParcq5rhPRgTBu1vRCopUlcIarx+Bk2tF4syztxLBgMa
FZo0Tl9j7+6dwDdbUmuR4i891QxwK5D4xnkcR4IrMqCPsv/DPWy5wLCQG/nudBLG/XwqJEwFLpiL
3UUYr6Cam/7DtZS51/TkgFrirll0ZEynyW7MiHBt1JRgWPo23XHvnyrMSv+kL0K84KGh7ar3rDwj
WpdYAV6aMoscqyrtWXXVrDv6SebnXPdCdxLivhW3HEOYx46qOe8r06U+/uSBKnbJ57ibPAPuccvo
2DTKwPs9b6W0lQc2g2UBFetsUJQkHnCDZCRovVUyFPEYUhgqF7tieQzBTTF+GJrE6stOXQgvoiaG
lY/lrhIy+158dilJVFLEI+7SAHVyRT5gfZXcEokJqt6bB8ZMDuyujFkYEHQ1qCB3sprkXSn05StH
n7gBYHWVewRI3YAN9ucJZC2qrXBs2j1HQqSa3ELRv0GvSQdvhd459GEddaFtDwni5OmaJ0OVH2g5
f1i3FazuCWpg0fOIYWkUH4nUby4VKkdK5o6+362Z4lBJTNNAZYAPGU9+6887rBnjCPpfhm4cHrHF
e2m8FsuvKcfhxNh7+LJ0Pp102cH/ZEKxphPKmwrLX8z1K9ILaW9w1qRgzKHYqe1bq4Ym63M/RSdZ
Ug5BigxBY07l9M/ljQo0pLePeZop8pFbPZlGhS9HbArl5Mqh0UnSAFtiQHpk2/GnUd5mGr8C1uvL
wrTNcDZpi52PgkOWdX/PLqiFh+M9EN7/M/rbqmFOnRAfat6UJZIOsj1nUK3NubSwnIbvb/kiJ8Bx
ADY4zNess5HVRhYGKepNQIUuhHpWDC6+bFwjxAdH0JiiEsyfgZujZ0RAA3daU8yta95FcNlHbFmq
pGr1/+s3HuPHMKQiJ5QOfwEmTAakw6l7khdbTFmOmzsOSVduUOFexqWMMFokGPmAjdHkou0uvqEB
xZ/yVUzKZE2mfcG8BNlSNxzd9/tMpQ8VgWPiHcZsETSJVljQFdrk2uOKLmXBvUrKhygMYtNtsAVO
cQYKHBSW8QGrFNR71G1nTTfMF3ViytHTSKab09p52ejmHpjX7jN4MxXCTorpqJEKsHbwAFkDaXWR
N22oyNA7FrNf1eW+xNoTSxFwnVRn/S7uMQjAqJE4vuURTaFOa5e9Y1fC5m1QN6F3a6cxE+dZo4fb
/emT7Aox4n0OopGc1JXkBO5a1HUtTuUvshU7ipz7nQh+SOlP0qv7qX41m8YldR3+EBK7j+reuOVl
ffIMnNyN7sYBWSOu86S/XK8fsag6ok95LyjHXDIv7pdG5itqB1Ro2c3GDsmrXXINgVaMiYf2mA+U
Je+VAueiW0g3KaM5NNCWN3bDf0LGtormMkIkjz7d5fOmqek/2uMj57mChggHOrMuWm301PS3lac2
CZPsAY4z7YjnCTaszH6jAQslmkCjkmMmAZCzglERR3fRfir77iCkXt258jbqeR77PR24QdFeobbA
kvaXvwic0BQrUCzFs2bEmp06cLK2cukVW+ko/+qxyd0eXaaVzTE0r5fyLcIAd/h3yTUt2Ss+zu8I
HW16+vOf30CdO6fOMr4bJOxZt5gJzuqMv8QWWuOTMwJ58/VFYXB8SfPTxkY0Ko9Q6fruMRk5VWeh
HPJMC47gLOV2dmKjfPkv3x9L3Cv9KuaH4WBSqPEHmHT3PPkqxVNiF4XK7sXTDs7fEmtJTzTgLFE4
yt6y5drTrUfvj/Je+uHt00fCAkvy/SjGcdslrI94LdflN+AOCeZTpx4TUe7KKqVxipYjpEnHGS66
YC93i7VO0hIjoToReyRWD65vhvD4UdDlknx/tKSWYCaxqKfGkkTYn1ZI0Ycp9A9IwGA1MnJOJ/wl
qeOSetZXCR5Gg0Tz35dXuPijfRylXpd/75JtPQNGz+4/ZX5uBXKHgYriipQNH7ejbP+47Flha35p
cvmnXt4zPH6dZjbWDJk8fSq4zVXsqqFJGJxvu/laN+WNDTVnD8PRMQACi2gog0rTdKP2/JfER5vD
9o73W7yvm8Vfho4/nnHRfJtW8UQbr23kqgwnStwxR5ezaoiM6TVecVi3DjSXx3++Qqk+zVqLccOc
P6YkbBHNp4B9Yf2N6M4qnLgKAYM4HsgRgJ2wT8mTDaIPD3s2uXYFPm+74FseNZH0BPpqWagOfKtw
iwt3VyJtQGzesfjt0iQ4swe/5fJ7lPG50YIJcph9CADazOvlfwZbhrFawLz55nicCdEHZZLHSPPE
bzHTWO62fRjW0VEOxQSnv2rwtUyFnzJ7Ya6WB1OkhzX5f0sQD2KxkH2O8F8ooc8TxybjWwn5W55Z
c651yKfsdExQ1Ry1PTl9HQ9/vQmGwjdLOzAnj9l/8rCml3XxtEa1No29apWD/aMq/pCOoueTA0Bm
bxZkHMxSMi391qKmZ+jz3nZEHGjOsAnpDE5Qk+On9ivQfYbIw8zCDI/sjqa56oxhpJI7KaZ38+7/
LfxzfapXxOqoEVRKrPpthQRJeE/0PoNzKj10/PHwgLymGyHjlBRDT9scr15vgAJwJdn+zLcz8nzO
Ekf/O6HAQwZKcoRC6xBcief92Z3VjrYmw7G+juo4K0/c4hM0kujtMwCAXjvo0Jyx4xLK8w6QWRI7
f+2ZfRaLrLcVR58a8q96AO+DHsLnAGis0ZxvK1mvwLFXuWy/0TLA6G7QYdpdZUHMslmDyaFYQtDd
4rHUxQzKYASQ+C3Ff/DZodBBt03hUBW1xKVmflzrHefRIIsZM0RDfElteUAUwM37EWa5I9jbcauh
oyZkB4w0HyHuYmHYOflWjpLBPyNXZi0YWTmz4+IheJQ8zAiFtLsdDZd8bPU8PbogJznb0vMrCuDM
XPKgyGs5S1uM9U3+UPmZYToxznFjPRTkjICeBSeAoCpR9XoOzOv4R49+VwnD0nxgKOb6HLGhTh+e
BBTgy3Cl/TRoUl3Php8hyKQErEZnSC3u4ilrj/samfndvLJx99SaJHH+oYKox3ZUOI7SSvKoA3Dw
50EPtr3K/LYHGCpAlG8hmyYKs1ZonSFfhoWdcUuHM+iYmYz+UkLSGh2B9N1fTRpAVUPk79RJS8ne
qOs1BfkL6W171rhgK9eIxH300g5TZwbWVUI5GLKNHbH25FN+D7J6QwygccsnUFjGCHqQJh4uMcAy
t/UEFzARzgtQwONuPa+v98G7nhzNI1C7X5K8A4iU4JUYFV/jmV9O2eklDPp9cVQ0pNIPCBJvEyED
0cixB0X/69Aey/dnYnFJGoBqmyJP8p4Dg1zebnfg2qHg3frUbDrDFzek4r/8R5zefIIADFhScUC/
cGedO80+1+pQfr98cUjnwcnQcvq/FjnAntgdwHCHLayFWh1TzA8JXullA/myhOSD9CgNXREhiJbL
ypawTCqLHU95OjM3L9VJFAUPuZoF7IRmMqA4LJ6dMsVXohfWCKuPsDIfakAUZp0BEK8yaaXwuGgH
+gCaPSEwNSoJh6RH978t7vaLwI7exEibCmHPXQZPOcAc1s+HxaCFYZKsGZWD6x/qxOMBl7YF3w2w
105uxud2yLQfJLQYjhRsdQgvwsKJre49P7Hakg2rc5JSo6eI1V5dYDw6yyROx9TM1WkKXBoaVkL4
rWQobwbUbmPHambUim9q0x6w4lkxbcLW26ewEvBeHitf6LXvrDQRC4vNR8c5P8HJ/zNc/NioQfrZ
vEE6asm7Rq4f9vtDd4DsLAKCAyjr9kZ7j5AOL7MEnr4wY0P2EOfqZaNdzDVnDv26fKO4No0aPvcS
8IOkp/xguQ5kkMR0i/mrfwB1qFUGJSZNRDk8TutQdK7Ib4bQzlVLD5p/v3MwLyx5/ELSk7reKdow
1i/I6JlBVQHz47xigLcWzFY7vIvPhOZ9e56vUB0ZWzzwxjrFhe3c+xFjvK1B5mcUslWTRexHL3Pg
aXj2yc1EgwWG7kEgFhbM8ZOD7B2ZQ0+W7U6lnTj/jn/IUcaX7nc31be7W/5+lXNAK0tSCpOx63LY
AMeTdEthX1J2j2570f+7oAnfEoOsvYKng6pgwBclw3x4wLAh8dxDy7KYq/XnfwsCbO7d9l1OFXm7
a+ZcLzqvqa7W4lv3x5hUC3LJZ+I3k/uMaFuiYk7Eez60YdERRNxwKh7tPXZFcW+HDrR6Lu0rKFnd
i62MJqbm+89n8daJeDpM3JyUFhGxfaiw1yx0aFpUcKQKjX5xy1ykbUL/F+5ZUVTe0Ys+D+6QAeqJ
rrEo0VFEpJHADbSTrDk0YAxBdXSRmjvwPx2PuQbuUm/DoGcTmfaby67LwkcBOh0uZOIJ/L5QSw89
M303aKI0fNmOFSwUb/7A+fAR0POvBlWmONIVyjR9SSdrTiV/NVyVPnEF495V9jF4WaenPnSredXe
JMh12bt5bUMnQhNBx5tfAJ4b8iD6n7AUvWH7LJIGZZvcwLTKDhOjI86PBIqp5lPj6UffJKKKdJSO
pTJ4YNVbVjcr/kgIhOHyPjwaVaPad6KJ4mDZ2dYBrn+yyB94kadfYG+0MUZjREL4njnLFTaFPisH
KCHU404uzKRyBmLuVUFY0gx4BMetlapuwybkta9v8mwrRviERqLAvxJJ7eKc9alN4NdQr5oMuO+0
/0e+kuKzsO2IzOYnVba0SzWAtlJPqAj1w871fM6tBnDwyxsTG3dXDk/BUjvs8n+bj4fTsTtrBXFC
C0VM3ZWD93HSIkV+O9lOJe2WyZ/XIJC9TkoFQJNrzqSFF96iOUs1V0/WHwZ/1FmNCIl/gBwmg7rf
CokBpMpGiUZkYHo0w+yrLIiTBBdVS44MGqv0aa6WYw0nRj3DFESQn6EEW5l40qIL6c9Xc/XoHOqA
0ZTTKEhhtF6L5uAAqWX8ZRQ8ChftHf4qjWXBeh+hcd3JZC6BhlokT/U9SnWCOYh7sIiZVU0Xeyko
X6ces6k+yesXh0Ri8VUZrxQHPUi1VjiOpUlbedSmKPtJm/5/6kNIMb2pyAa4yN7f15pCDuIxcG4p
nR9LdTFLufa4EP3iyTyAs84MnYnxVN4C5sbbRcyeh3s0VIR+cOrzN2g4fsnA5a+XO6Xy1CtYNIYn
kHfvAm8L5hIcqeA1WHhzwbhfF3apqS4hSwHCM6gFT4PTyjN8ODko/EYaz83NNkcaCH4Ps/G/wnH9
J/Ej3efYESKAK5Ex/WT9U095VYAEaHW9i7vd9yXZyZD8JV/m4/M5/s6UFOVPVJhzCQnb4FysZR63
lXvxMO13xwEcJA/564mr2j8Nrw/egDdUFgPPLoovLDA38krGjxyx5ommsecKnjxtjf5e1DRoy3W2
E+j/9koHmAS54V6TI59fwuUDISjqs8kunWGVLnbzTfPDk38T3txBY1yKM5e9pZj/Mi5bw49iADoz
bTgAruvKon4IVrWwtHqxP3RkaJc1MLCO7MWYo2TlwjcvY41q9litFgtq44X7xwo76FzyVr/Z+Bg5
JP54R2KU4Lib92tN20yeRqryt/kGKMkMcij3gxGn55gEi5jLUUlOhTeNVZMcdUJ8JBl2M7NdQ44S
huzwLD0WlWbFsDVATzJxOI2cBGiPiYz2QQWyRH/qYbkRBxddHLQGFi86ZVm9A6sCwfLNUwECQYI9
Gss4Cg9vH2fAEWx39jq8phOEFwgpe7N7EBopTcFuDVyZu+W+FB+IS+9EITm3P84BpJdA3Z0iaGZO
+p3Fxc0dla90IHDQbNchfx5Ntg3jc65l/ASYOu/5v201YIA3hH4TqwIHaWGEz2M7Hbyo8Nfi64jy
PcI+ZNqswAOhFrXCdx9LS7cyclNLS/e82sodxbzm+wu45oP0Myi+tFSsux4yoAm+F9le2dyWeqrn
LemJNROd82Sdq9FNSEvPj9ukh4U5Mv/L3/NKwVD0Ggq16/igpJM81QENaMDzLDKf9z9qQ3wdRt+p
rSKaxRLmqKyqWwNvz0GrIEj6F/cP4B173AtQCcg/C18ZgQZ+d4UMezUPK2XFeaRUZIDvCzOOMxwU
V+wmsAJEvVq0nbnrZfthJO0nzrkzqLFHfW0MAiPRxTbIn4fHvsr2BNaDQo3hkh0yH6O3U4kRfnEQ
egGsWyNqXimDyfd9d7sq9ku7NMj0N2COtFAHrzXMUfZHwE0z8vDTva3CJ5aA8pIZz0Eayx2C0oOH
HtYTEoULB6u2S9iWfe0wSra/qKUpcPiDeMbmP1F3ujZhjp3fDh+2lvvTTX61d78lcq+FwWoi63Qj
mgUwxpdzyqFyY8smZeCC1t1geC5hnB/7lu9RR8qUYJ9kZeaDIDXIi2LK9m9f4Lnkm8hiCUFbwRSd
s5HdjAMW8DTtOCUTOBIy5T4hvaIeBRJtEKbexZ0QMhGG/3L0Gevdnjuni2ZMFEEd5rkNcbfKnvwn
+4Syjjs8Yie2HPdoV8u8HxxQ/tptOuCNPJzuUvHuIbbM/JOZBiHdUu8SzHgMK4/9P3sBoMFzzKje
ejwPc3TKrfsetk5mDUr/dBsobUhEVQ6ew8YHT1lVC2xnOvpWpRZkUip9Wzug70FWWNWbR2SUl3tS
Ih+Bugs/sEEHfhW3w4RYnarZbjrwrtx5+Ao09vPWdaQvuUycE3RPNsI8eFPGouRo1jTNqY+rsVln
D4mxrM+O7mxPc16thbEywBbxibO0i54tTGynB64KhhFM8ZbCgaOV9tBuo3xiwbNgAfGXNKfsSV6I
+g+TaXBBwwgp7xWR8P/z4KYQBVA8TRfmpDx3vd9WSdk7lYkvEuNuLnUkEvilir5tMxpQZs6EPmqa
ZA4YtZFVQ8+fnjj4IweIXtAsTaf0DJBQS1teb2oU8mKd/1p8ZfnBYnVALZ64eeJ32TH+Dah7fJhU
XZdJvnJB65M6SAB4/VpZhdcIdxt8ZJSBG53KP2ixZDP6XDONtQsB4nQnQteKWjzT83LsNtuL4j/E
uNbnB9lg/2yyggnVeiaFLAFI+C0OVnsgWI/7K0m+3tNYSquCbpIa4vnhMe3HWu+vIbdkQOmctrI2
MUiZLsOShv16ZVtdpG+uNgEOUe48GF+QWYLcuzuFsWnmBH0fbV5UUvYlVA5YgXob+3gd0bLMdDQP
c9T81RK+cme8BdAC3m5cQ6gWs96ogX1yVkF9mgfNjPASKvhFNDsvs+2PTL36RhpDqtaT7ySZF7oE
NsmL1/SmeIthB7smcQGxfrutwUQUj1dVbjpSQNW/N9qo4EVOtUaCbFnafP6tSqiOAG3JIPNf0BXt
c03aS/theT5z5bNJdhELu88Va1Y33FPhBe5RMNC+XoHikFCn9hwOqHXAA8cf38UxkOP2lxn0XkQl
2PdCJMsgSeaP2jgGVHbgQ7YSiDHLMXn0LvdSVGBuJxaBVf8JbH3hcqCl6nTR7j9Hcbscnh5SUQyN
Tb5WkIdBhBnoRQPBEyHJ4QzUkLr/+xn6gM/E//eZSiTQC7NwNfcjaiquWw2nMwLWeDbA+gW0besU
33A65TicbVIre8qxahSNV7tPNrgeHZtULNOZyS2N6CxVVZz8hfZUI96W0F8fH9xUZ1VOahfrpkdo
hRigmU32fao7LEStmKyVYiOJOKjeOkNnYo36ShYd1kAUFcdOFIfOY+xLCy8DTRbRtLvtQ4l+XmfO
C3WSrles/rSt+N5wD7L/ZxEdLhHrQZvGRRxuV/hDDjsAO+Dvp91kIXjJxfEQi8cGrbWHed/v1rpp
gAf2QpHXeGZKTsOt8Gh3LJ39tLh7edGaRiDgIEwjy9YwD8o7qTQjTOsc6w9dvcXYTprzc5lCBdsu
TUN4pv+5yMzMnMIlEVOMuHMOEZMzEejRvrgYy7GnB3yYRDLbrcym89UnpO8+QNn3RXVA7dUsyP/C
BIzg10ftM2L6W1IKm5cXwLaAwk6AfzXRFVqDFK9fXgTG8nUKhSiYqblwuGYgKxr0ny4gV3tfq+g3
4RpqMmVj7PGExJD/AnmRjSccRURnCmhbyOrUlwW0l4B5Ix4gsDvhC+wHAKNYYsBG93ynlYcB0N1S
5rac2jkRLmrZxK67e1QHUAUplGP+0ayNL3CYvWrZsxZwoorAEQy1llcxFazPPAcQV0MNdhkUa/wA
gb41kDwN0KqdG/lUJW5uis6K0u5kfd3Qj0KGalnkWOQzGbok9rrMpfbXPxTjAbeZCWUCr9aWyWzv
uCcjar/WFOrR+DdMVVPPxGdxi6P+avYlCmcMgkRb+STv8gwdcr2EomXLh/jnD8dQBqN4q+w5dlui
DBQX36Da3U0WxsvPzru2jahuWaYwgBGLTUUIvr1SF1GBywiF17BEBfhVE/SJCRdsX/urWwRLtpVp
sE9SWy6iayDT/Y31er1BYMZgwTgGAGexQCSXwVcAvUEUw7nGgCfhM3YMseD1o8JpyuJISZZLQ/5T
txqtWX8jDy4fPYtjEALKyCulxUbx1r6qYOKDDm37wz43DyDjHKH1tNzy0Arxc8w9guSMGtI8nCcf
rF5TCfYR5tXJQm0TiHe/ehFkwnpokBWyuI5F+MnhdUSIipMCV75M/kf7tV4tgSiIQ6gtZ1hykwwr
0RTqtQEPvPuGOglfUhJBbDR8fUrdaKVshh2e4rbbdN5aK3Y9Qm4hPnJqNHQJr9pe086/3WisJZ3t
Xv9icdPAynh8slPHE3CArEuZaGtvjraWyerdXO/TFQNEF24837JcIfVmJev+UKGeC6LtkSgLrmH9
852c8K8Pa4GNv4ZLfV063KzrHEBFFeEnW+GtL4mH9kVzVMfvJhoM9v+/KjikrhMbAtF0R0jvD9qR
TxHKB7URPlFTkq2AIC0R+y7qoxT6McAO5doi4Qi7bELN8cX6VfHqW4EuwscvOVAqEIwgYmeTUCjt
GS8kEcjG/vONMv0W854VWtRwfPLskUw4JjZ8vWKcXzMnx2Z4YnZmeZP/Y9XbxgmeO1e+yMlcE+ST
IxcdlrVsfYOryQhckZlkW+sSP8Fwy9lQLUQpGl/eeOTnkM6ljjosbbBzGMmvVdJFoCI2Al6e6+5R
ST8nku3cpEcDMjS12b+pxbaiFhE4AWi2oUOcXLRgbsK0MMuCBzajThjyVI2n96nH43lFwhmU1yl9
VPywji52/8cIH/hQjdeGOtAXPmdcOV5KAjaxvSO2we+KsppNFPx4Nfwjz5pr/EOno4EII9INWj2k
uAuoQt/JTie491Mp2e1uVTQ8BSDLOaAi4eaHwk55OapK2Gful0qGu63hiURpboZxa7IrPipa9kp+
xARsUhIp3rFrL2tu5RzvygWoUUwO9kiHw/HW8yZD3rQ5+WMtmt9Dqx2s4bJJV5s2jQ5TjvTnI+bi
Yq0AYKN5SuvdJVyoLirdOm65WsQNNW8hCU9bwVTtZCrd1oT6qEJdORyHnAHpI3rcl/QPs9/I934a
48XYndQXrTyulpSFnNbu51ca554bihQWwvZs2X+I0MFIJRGImnbO4tP/1sUJJvz4S5NdCrfP3xaD
DrMXANSb02m6T9MCH1DYfU0Hqn+gLGeFuQNzxtU9xjDIlsN25S+O6U00U0+/4I6zRfNm2ph1Iwol
ZgLKQ9C1PEM4ZJ7tTzI4Fv/hHMjPoHOoR9qkNQNx34bxdkbibIjIzfo9r/FGKWzJ+vQcUHJ0Kwxw
RYD+d1AyF2giIzw88OacVjAe5pdz/VIi6S5cUviKiO5zqo7mVpYU+486ixsENaXqpYObbNcZrXrj
tFjiuPMuuTLr8ecEoHBqqKxB9mT/L0J8Dn+kCCOV1cC2S1/eobzzKYmhVUUJLIgiMvfebAZJx0Em
W3xNQq4IUJH1vKr5+izITvSvdD6WtykSJp9Svbl3htK1lCIS5AQfGRsyPp0EUAIX5FFCKSO9MzaZ
imTKTkGJgfvC5jyPiSJ6lCLbv7aRkpOabK/txPDATVJOFbgu8lxjg2BYNfDOGmY/A2nyRMgF8e+S
Kndouhj7ec5VT3c0Ijt4g0325XaB34Mhkq0ofrMkJXFDQZpLhUkMVD+2+FKMGzIAfxpC2uEEikOZ
CenYR1k2KE93qnwKd1OhbB/T+4TlHR/JPHa7tNgnhImq/FtbWZuK6PrJtKKB/O6rZDCyDJ1S6QxY
41N7RuRIKU635PAnYOHKNWp6TmL7gtT4iC6mJcK3vr7aI8FSGNeVoMExeo1h5JysrNBHw8qy1TJN
YeuvVB2l8rEF3Rv5Jc9sTSa/wcYtubtfJWzJUs/5uSDYTwshSbE4pnw6sSp9r7FHLdSdCF17C2au
mBlvddeBYpdquAbNVrBf+8xGxRpa4RBdpX50pGqg0O/ywksTSArHF5a3MTHOuMCMNM1JPwaLnLv5
eBBb3X88yw3b3S4C0bai/ns7Esa4u0+EpT/Wv9DQ0lbR6D/aBeReC9pxWsXOT+11hwFGE7Gmp+gA
8+OD+NwWtLWAuj9AFB/DJ4fbTE8SIylUIyLUEf+/8r67MrIkAPItRwZ18JrrF745dmmVUc0i3udR
WH7PWE03iOR5AvfL2uM231WrqWJfb+E/00O+YFfi58dxPvHW3jBAyBpUxAPcgVFS0q39XovcunOo
9viKFucSoTJC0meKEa2gdfk8eToZU/n1dATShXHBYrojNu470hAxfea23fkZPyLzLo/pvOl/JYXp
tOeS1IE0ebAa7tpGT1jEAd5VwLGDcrI4MDcZ0XBP47nWP3lq6tI5UryAxiRd6FOHUr9KPQXyVXGI
Al07h0AfdhrXn/k5jcb+45do4G4p7FtyvkQYTPsH6AKNYm+jCXE2eZG+gJpv2z6nahRkS+jYrhov
HOJQZAWwImWdlma4Zsdu7PngGTKI1ApIfMK1JqsIAqp3ATLOJszFcnXp46/DYoDKJRxJlhC69v7K
N46hXReqCnwBy0eGZYYDx6hdiw/25gzhg9XynHC4rcxbII82Wkhjm+Rv2Aa+b1HUkFTPq8hV+JMv
bkbQnVl50MJHicquSD+SNOLm6tWuGexFORFscUL9oh0idaVzALtF7t8nEjqi4+lDA/iFOzqexL2C
UlHon76rHTkvpA3NAHOJYjnEOr6hmal6ErR2N0TogtRU+/+PYa4QgoGacQYzuf2QgqxI/frm6hhG
Wfa3Oi7olUanH65Y+DKUx1RtUFuPJp6nTt4DScWrdDhpLFiw+csK0O1ByQgRebabx/P0WsCLf4Kl
2slkfv3+bGwmKcS1miCAgqg32CwuE6B9kFxWnHXPAvf3TT+OhJ8ii3JNpFa5rCl4qXyFWyJDDki3
nMzFOR0MvxN14qilLHPTN27zIw+OpG1f79jPan1YjLQXHk/u0iLGUROZ+HMOLPZR70Fu/Iy72NJw
snXyZn4SNTbNYOKtuRZh7ImuWDCjKd5+c11IZ2HLYfTXWJ8mr+uTAzUy0G2rDOosqmdyd5370P9s
6XECTRTlsOVFgOLFqawFu5gXTNmf84cII5JRl9oKsxFfnPmadOwqwAxuz/4+ibd8Ugp9YlsKa2ZT
E6rVWHUKCdR2XrIpvyHjkDacoq7mOBIRdxYnlYsrPyI7A6KMRNmkbRUj/6h6ZGc64yz6qMr7iExk
5Fxt8dDqwsopo91I5nKmVRDzUgK8br+d6XU2vN/GXOWFGi0HnjlnWr0+sHMgN4Gzr/8S/fD1+oEm
2EyAMRoY2a08bHHcyyJZumspnrQPIhwuNLsSylaTJC6FtmarsK26oz21HJqjmSdekLcQ2BW1gjK5
QBzW5/mR8O0n1LRTtFkj5EXHVk4qPIwrjclctKJdsSydV49IIRFJpq5csJfkAl9G4XS1qKWBiTYr
Ycq+5jg2ByRVysfDF0t3U6+QG9xcqMa/Kw3P4MccWK4qyNbK6biorYYOXPgACw5EBZfT5jarJraC
WDHHevEp8zCvprcGsKsaMMFzS+V5O2dCW3Z/vrKySOZnkowvlanMUjBXIfdO4cEp5gfE4g1xocgL
k8/oDg7ovG8oCBnoqTiOf1j0VyurUBgaRIP5ExeJDhWjSACCwO/jQYcxUJ1Dw551aw+Jq+to95Bh
5v/ORq6TFh43pW1Bmx9pysvvdSlxnn0+W5fjz4P+N0A9mygZ1DK3CwqGEC7i9qrSySSb3MLf04Fv
W6sN8b5n8pNzHq8vcTMW7gl+2V/lq8itSmaJGRXcdI/hoq5t7BFIiPPcoOSfNxvqzoFMStwYva6C
Do1TIutU43/QyH5CBp+H4zAz/Sy4KBARb8aL9fQMoezkK6mj8nmZZFQQvmmb8f9SRKnGPHe+SsJQ
do8uYVA94B2zjCdkbrE+/u4paARdHkth7cq2zwPELmY1csQ2Abv5ZKtn1zHLRBt79B5cAs4ZlEsk
RApy2tAQjLYf+Xvzu2dqtLjXSIpRwVXNf8gJCcvuFdOA99ZFFZAc08EliH7Wvliai4nO1gQ9yhSq
aRH4NjajFjAK7ECAD3fnBbJXFci5993n/b4Vz1wVkH9p+/6VS8I9h067xWTQbeo6VCPORntaBBLv
eAR8qr6hrgy5Er7eJ2gbwu01lBGpKl6k8n6yTtkTPTVMN470hvN52i7ee017BGbS34i3Ufp9DVFi
6IWtMuOJoy0rcYti1s+KE5nxhq4FRcQQvH88x714JtbMbKZs3GLhi8+wWbg4uj41QAI+H09yYRTA
Gr5BvCAgraDpIfH7u5CmsY+8kJ2zSnC29QpZCrdnZmR0IoO8sOPXb+X0x+zrwkqc+lLpXhsePI8/
jWrwMto8KumJTN7AikmlaWz3v22Pa1ag2PNdpb1+/dCFds1ZcVr3/9lSAvccCTHHdytfkFfPv8tn
HWHcxIvYUyz9/KW1zPYd93MbU95GKBkWClviLLueIa68/eronc1pHveMyGjHJKcfL+Ln9BsMWTKj
qbZNo+cBm+GCvNenYfZpL/0QO7Y+fw7188++Wr5Ga3bOx5lFVBuHg0NBBN6B6ykFm9CBz96QVF7N
a4HMK8nUvgdmtKZfytu5xW8HwUAdxER06sfRd44W9UIE4VRLY3+3h7lVjWeAeDlQSU7iySxcIIYK
vUHGv9E49gRG+CnNmhSJ6UxBJPIDClgWWuDhoHphb7/aP6Zmym/t8u+HGLgBunRwWrRwkZZnOyak
EJkcZ/sZKMiVbPTjcpQcZXPb1xhIEHmvfrUtwZSq83o3L1tIsNHW/wRsvd3Hf+/Uf1+obJbBhGVv
sdyApxRReOO8onG2gY61MszaBZfduAknJFYi//VrKjzkIHfkTsJiaipJh2zd45O4LIfT+sfhJN1e
z/nIHXHoykzjo5RvdQRH8IJew988/5LaxFODz2GOm1wS58jRkJLKMlGrRNzTP88i0rSJiImHx03T
vCuB9O4hm8JzYXZwYBKa6xqAlIpMGfWIOYraAyOzdKrFjLcm9mFNAWtS8eZjHXJGcJi6ltDY/ynr
jRLhbfUZyX/wl/mu4gSCD/IekX+G2CPyySIQBtHsJOn7SC5rUtosZbja6F3Pl7Mp/9lwJvDcO/Et
b3Vk1Zs9t69SHir3fF4ETsovjC/XbekoogM/WTobTaIrLIxC3jl3wWe8L7E4yoQQIx8xdB3jN5hm
IW6LIWg0Qv7JqWqi0ncnlkslwJ2SyPBLB3z/ONRKDUJTV0Z1rRTIXxOUvroWQzHic1xb1irfRpgg
dlSA2wPWS8v9OWA0q1XHZ1dFFYaEC3gvAJ8y6YqpTGa4LSdWEl5wX7foRPvma+0SFcZaB2J+6/xX
UiH/cA+8IEkTE/aO0wY1j8d+v/JHLkf0E1eLeSWKUUmXIhCt23jJy4ELLalakdtom6hS9Y4WGz/d
Ynt2uOCFzghgvXU14dp/ZHxa8MBH4bIuWVNX7aPHIxOi9qnt+7FN1Mn5h6EeaQ8Kj1vSHlLjlBIT
VBARQwRDOF3vnUZuEPQy1QjY6OBIZh73LrOx6bSiXjiXGEltvCMsRcqA7BUlJVj+ljmpox7f3Nj1
WW8gozWDy5JeR8Vw6Y/LJ5GIBzFm/EByzDdt6DSjfFHoRiO3AU/tCCH24eIzD33U4c6QIMhamucs
fcqslxw4+hSH0FobkIOG2/kqsa38EykmbUW92EDVG4PUVI/4kDw5XFr7KJPVgCHgktxEoOCVPmvm
7Vvmh/WscwO5+FDfHN9w0M6DHGcisjwAus8OZos7THYR2gghb66WU2YDXs1o2Uy5HBbOlsmfQ6+k
L8alAMfE96suy2xm7RkFw1BH2E8hkkMZHOsFg6olJuY9xHuvjo8IfcfWPhPfY6R/DKA6go1kDSO+
KnUhXNgbMxmPte9MVEycCcarjFm8gTm5IargqlYGZFNSv3LasQrYFxilPVRuqW9+UKIRvZGCPZqx
Cw0t6H2iuHLrtl+j2/hntxFowcGc7JrYn44qCC2MFSmQ6SxdI/Sryt1Di6fdEnxoLhih5YugG9fe
bIw6TU5KF1QJrFyjyWKZsBnFgzXoi1dZ4r0GnTOxSMd1NzJiyJsxSUf2ptHB87YomigIG+nintuL
6Y7rB4RxnQbZnWfWduri2FsF/qai45smUbKjuFwgDfOvoupzTgpC1meefDatw4dPy/7C+SflshRv
ogMKGbHpp0um4irLLOEdTuCZnNe66euZ0zZMgf5c3tXSHcDmaN6Cvs7FeHS3hii12WMRcrFTt3r3
eevlUamprmaSBemgV0X78GZ0pZvetTCqAd16uOsD3H1f3mdmrC0pgcAPu3A4X4PQFYCL/KnCkJME
DlF4rqp2RRlH89DTTAs0V4U+xlTMgcdSxiLWs0ofrpkR0uYe9kNrAxkYvjiT23VHTkZaFjeg6651
mBwoN7S6EBURxJliph3BGumxuJzxFT+vhm2E7SpqebewDyyJlVeFQdq1dJM1j1RliipvgFanLzqk
azLx/srhjPkVnpo46IMCvTyQt9z8QPzP2v7hHwa6NOrJX+SlazLWhjHWpOQ2kJbi1KALnp+GxA1g
ToqprTDR7fknGcElPL2LfgxEN0vUgxMmCHkvaDrKcUNCi7vre31F1Hzb+fcIChCIZoeD+9QFG/WF
N1vUrB+BThnWfYvnVk3ShDEvGvu1AVK/nud11JFMUT5slajL5ZlYz5KQq5CkmL5t1G9e0nhUtC/j
PvGaLhMsEkajJu9BAvOpgzoUGGSaTOD3lJ8xjAJGluCI5H1zhYnzFa4rTmR90hzU8EoLtz36sz1U
GvNyhif9yYNFZe/7TKEQm311Kk8puWcRcy94c17Kyhk4aXpRvKk012kT/VLR+J1CKbM0jUkJv7VU
p3NyFJlWr5yaY9oF22snsMRj5vEJMJpZGiYrQS08jiXrTtCTNsRoMr2jLj9cg/lnjT8SCGczTMFT
zIWYxUjd4VDwhmsrkTtL2PdF+3e66X3SghEzEQFAy4C0EzHj47hpQGS2jAn8eSdfijOZjijaSWxU
gRl+iQBfXcqEVrNVWKN3zfpSgXWRX3Fwc8oBpWzWnjIm5NR7Zxza4GBwLzCW7rUN7zK7aRqPDCK7
AhkfEe85kOpZkhRTJDUzkyCjP120iTBvuCp438OFEh96hFdK1c94Bfo6UpQ4ncdYpMG/+UgJRfe0
rep+ebmfwQgbGVw5LbX5Uit7yC30MGwzl11iUMTHq8DrGoXYMIpf1q3F1UNGD5oSH26uWSlS7Zm/
3TdWMvJtYZgQLh03RcQrluDwfpVv1rwYEetU9rbzBLPYZHwQAI/RU+EIGuaufx5tetZPQNXbHG+u
fTjDFxUWUDB8BNs35qcKuT188WtYP8zmWlthaNUqJjJ3Ydl1LbJKFRftJ4pYhrpB9qUWcwa70eY4
6LLyS5o616/5N2AMxSYOS8ZdQcBuXRsIShYYmimLN4M8jBxYdpz+UfGtmU1E/ppJtHiGgXOLXyd9
EangQMsOTuCIHgBiBJ7AWSmRlKiFaaL6IWuWA/3JAD0TuRQFYGMzXPobK16QnhP/aOFfVPr/kZgO
Sf4uJbPGVm6VEcnAmWDPjxV+JSoeZW1xFUfiYemiXKWabrmhHIXf2kDBgDMYN1tO6FfJSgUSfI4P
s/H6lEJ+7I60dCqd/qtcfgsoT/wdEJhb9Km+0oz8pmc3haoDrmeza6KuP9XLdrnKWTv9e1Sdkefz
XPO7mx9dYSJRPoc57WZCnP+eAVbIniehe7QLuWSeXfE25Nr5Dv0Rc7ZkeMHd7bFqkfIg4uUAqSKT
qhFJF0gaek1cP4k1wOV2FkKNp2oyMibwmFtQT7K+mx9ghbMpQKOyrT3LAHsgNxpXDnSCYxGfGXx8
Kv7Irej33/d1MZW6OfWwJwhhRM5AZwGFE1QdiVlnn4nwTTWbz/z2NUKKkT+sbFLX19szQLXkkn+F
l03cm1d69K5VMtwhu3lR1RGK/Uu4d16g/poVfuRZCNXPrRF5cmIOiyIbVI9gn5R1lDCJ14IqCRol
r5/gKVhpwY4t0Wzm5LGrltAuTYcBkw82YMvfxP6V3sD25rIOJnZPqZM6FslpbV1fhFBsS2daeMVL
INy1fCM+1HyjANcqgKT4kqJc9W2WHsSqguypnCpv/szSG334cNN0eTiyufteflCJWDkO07doKPv1
LyESxDMfKtHaiC9bhcsAW+hroTYPNqeRIl5dUd3IycRi8Djbbj5JcR8ZQY5+75tDtLcRLXaEbr9k
+td1DnfjK1ONWkL3zdxfnwbMIcUNFhIMFpSbuW6qhdo7Z+qyLGJWAhrBoUxDcR76PRTCVfMa76CI
Ho8aDOo2Upglhqh0R53APn9+WUODfEJwXerj+VpcH9B7m8dFjx06twFlzvaFyCh3893z9tK4Xdxn
oTB7MkE8tVDTUXeq2kRcizHGLYQ0CPY3EJ1b9/E8wM1h1zOjniVTIyKp3EY93b4035FKKtmbNO51
AIcAOVlJBGVJOeX+q2j90aP1/Qxx/3CiAlZQfeFtkaL3QOEB1ZNCU6JuLp4IpBhn2TUqr0eKBJsc
ydM81qdefBxvtBGoQlvoCg97sNfOiVVke+Efs2iKp+DMmSnLVtratc6aKghMgs6VvHj+RUSL1VP/
8wTl+bqf5+k5Dp0XUemWLNpPCVyEJBSARQ+5IrDXaMjDQzJWXb0rq1Ba13Fof1J8b9C+cX37ZxCV
7QzZ5NGVwfWenrJiD/ixNsTZNjYO4FMnXqwiE94+K5j7ZhtLQRd1xF75UviiqC8X8p7c/17FXJfg
L2ohDI3/8cO45GcCz+U69HqHN6AHYQdDOdxaVJ4zcXmfwI1ToUR0BhjTsfQbUI4mlksLpIixxnG5
NErg38DG9RmKdX4vhXrtcjwvogq02dJrDqYNUTm/c4LZUe1/zZnK+RRg0i3ty/OBtBevDwbRN8gr
i/cCxOi/k3H/lgJUhp5c8o7o+CQuK+sRGhKDVlTLObaDOHhDTLRqnFmAe5PCJoUOVcvcEDKwXncz
qD0k8uOPnd8MLCrbGQFV3//1rwAYmQjkaTi7n4L5RIyIogxH3l6OPGFAgMzkCeilRcBwPdZ8At03
IT/h4JZQKd369gnl+BrFf73myz39NmVLp3AVsZbsEL2W9GuDnsu2fyIGXJiN1RqfwOnHeiJcM0B/
RHbGpNGqdkWCA27sIlewhcrpq6SNQ4ssRGfu5ZqTjmflbehxGyMi9Vb7f9BRAUflwDGBog4P4JBh
GWo+Cj8e6DB/t54pJdIh2YSXotkMBHPueFbQXv1RB7qpSq1bVUb7KBYfWnKi4KJoxbraEiN8BOxk
i5xRoPp2fcibUR6wYwi1jFGppiq35PeQqntqRJjjfvVZyiN8SceshAOq7uWlzXGdBW8/pVZgN182
LyiiByFpeDHO/zj5WDZ3msfCYaTtv/QTY2WWFyIEseA67KvJUuG+ZbzRAFaiHB1apd3bU8Cf8Qzi
3chSFfCwhMuSiu9fDUJYGOVvJecdrGV6sJU6alSYXVjd0nMx69XMj/Hl5w/lhpyKUYAIbaDfaQHL
kK0tWLi9AKm36Sg2cAO4Q8SjGz7Prh81QiDYndzWEkvcgi2g27vRa//jrcwl7YkJAHr5m4+7UcMV
y//D1KOsLT8ZjmUQHNIsTYkY+u/+x8gFZELjRQeybgyIXzUimun//ClPz1m8CCoS1xPMP+g2JrmZ
9AS8wV4MjoEAzdLfvFTEEXKfhcelAv9TLE3mkfA1JLDVB3+NYxhRwfzC6N+MuAQto/ZdITPqyJP6
QqBLUvBB51WI3OeZO5pu0a/rFFx5z/+eMiBEkW0xh0bRPRN7soHu5dqJqZSirYWg2tvzf8r/3LTl
LTIiA+8GGR43nVMcpwrTc7hM6wVq1wIpUp9LlpJvtcpGzZDzrtDVX3JQvGoUMmXYq9YteMzQKjYl
WYLUQQCquL5nAhw0sVkoWTu/IROf9z2o9IKVzW1FKf9rQV/hwppFlw6k8XeOalZeklYghQRiXzDD
URhl/JsueC25meGFbzHEmvgmKwWWgWNOee4pHlkpQx+uDv25duRIE807mQrnp/EmrCFqljKmAjt3
+ZjnnpbOfep0AhqzVC/GTdn5N7GO7GHsKhEtLfF+eo1BzeqwCcsPJ7NNymtRXmO5nDzS7L1cyiJn
bqIvRatM65MfeiHQ7VdinmV3YSnohZSn+DKR36MbYYkbnC5/tlBnDuhD+iiJ9tKpudECYkBgFil8
YQNhygekDX4PpElhxb8f7TIjRI+nndilqn9Coc+m10PnUQ1Jr27h7c+ind8MEm+Rl7pkl8z5DQvX
YkQMMTMQdHXtPRADGCFk8RfeXQsMNKRH9ODlMZXzJKMleJ/kJA3yjY+ribdh10DD+IHZZKnL05DQ
5+YPN8NeaXEX7+LsDKBqQpyAret+Eimodk8zXa3WwDiWRX+a9ldwRr4BCmXSJ6LUqqYPPHTzpq7j
IlwbBqDN8XkJzqe6eCyUK4ycwPvkCpWTQsyviARZziApHiGUKh+Fe9AMfwz1v/BGY+GluHELSn7a
4gNYMA0OHaVABIJcYWtsBhVvZUCq56J5uQdKmk/Pl41TJ/Yv72/ker8UBQpw2/MTS5gvBGXu10Je
1sucHhuKkpasIarJbXgC/OCOya7sHduq2JrrdC5R+tefGYa2W++4ZEs22j+jP5Mcuyy2kXyfc0qd
2rl3DGa29XOOmmmkWYuDvo8db1ydSTe8guxUvwpf4BJ9/nHBO+172gzwL4iockbB2j1FacgDtHdq
xKHqyhwrfHo3PUrTwdWkc1yFpqWn/aI8myraWpbKjVj2SsTPK3FADPT2rNGmPXdVbCmzp4VJeaTK
ZnXmtV/ok7uRJ1whem/c3XXt1LvXHSVVgVqXU1fM7HNF6Rez6nHsd2QNZ6JWy8N6RxIq3/iANkDq
7iTDmrVYWek+4dvOQNdgK96peVx0tOwjOoqvaC88OfzaiHm0wd3oAd21ULhFLVDfsB0WfUcR3yYz
VA3XrA2uhCDOxIkcihL8vx2bnuVdGpYpZglv1e7qbCxvtRN0if8GjIdicETskcxlkRYtZ0+wBXCs
2CAMB+Bdl6wdyto1Ysdi3WC+CxQnLsWHvJhJHTVePib23h/iucPnBBVRNySa3a21B/R4gIejzNFl
JMN2VfW+v5cWLGCFfFLbS0BSbiCQVEIBDyKYk//ibUu7QDaQrOwfWOyAGVutOKkJV8XTY4ujnvzM
CGIGCWRlNXxEmvKqxc8eJN7YDvu2dpswgCQqqsVg53w6Cp68Zgu4AszWEO+EjGNFZgK1+qmmIgqA
VzVUjZUaZoLr4l2FA7WiQ5UHl+GhLp1xkmI4xnIqN2B24JDgKeQbeExk5RRbQPdvgqbPG9qBtJnP
O5z0fPao68Wrm6u7wuM4QpYwDzglXrcwjGDWGJWE064RzZaYsIBoFwu5B8jhpwcXTrlVnicFlLv5
cleysp7lBl8/BcHnxFeb6FbRk2y0CMh6Lymii2oSCUcIy72q9Vy8HUgqD86HICphj6Iu6QrZrh1F
JZKWY+TMvdlds4HypfXEYNwY8utUlfWPpM1Jt3NcfA4Yf1f4OS621VWY6Xzm8SBJhHgoLWfhl/Q9
EMDqCY4xRuq8EIbu2QyGt75mvNGj4pZVcwtNS58vOoNqJ7jS1dpIHbB5+3MDJgLDuz8zDkKisG9d
0gqkWMyd5Xx9iwXPEFg1wSs+w8EopwdKmBCqKGH96vBBmEOm3rjl6Que89Z4FRveXGCUgRTWl8e8
4EavwafFhnUJeXCnmIXarU3ly//mQrpA7RKd1RNiMvKWJH84YxaGgVjgWEZxA2grYVpiOASCv0ND
Dz+YDn3vz1FnrPmjnoxfqEn9rZH/THBPmM78QAHm3XgfdDsBlHGkAK1PC8Q9J6WuF3DUXhWbeVy9
DhMUokq9XKtS2zWGMM17iVV6t7ArjeWU5A5PqXtozgu6rvh7I0IaWva7Fbh308DAG13cyWwI7RVg
EU+ZhIEVNvWe82j7dAkgosMZ+3m9T385u+n/F8FCUOa4Mj5XRwVTTBN/ZeiRsdElPktYBS7QlfIT
zgUtN9EmVVb/AyrJAZnQFo9bktRc+aHZs5itOwcHYn3ZvuqjuiCLiA12xbcSVTara9KDHWWRPSSv
nhi/xdDS8bm2Gpll13q8IAmgYky7nPx4Z26WsyUmrUsmna2JX1qPfOh1ePN8XQ1erncKEg4nzvTa
eU4IRwculWMXjeZel5bEjpOQUfIHOpyH/fWh3pYOG5nPLEZY5VyMvM58l72x9i1Dzjaj3e+Nm4aa
zaYjE4pYY12baP0/4QtZde6fE4YTj+Bf+G/jgVwKKm3YIOoYGnRyhYn/CvnxXamXUtqYVSyw2rHM
EInzvhJzyv7FVfarH66jk9zRgzLU9V1EsHYXzZtJczjrT+8fobXqAlxGBOoYyXJmZ9I/V8fQ25jR
XHioGxXQmk1rLePPsq0RQMZzem748nHuC9s+8O7eETfncTRQTob8fHQLRoDH+UzJRuvBk/OogZL6
unoh9lTif3YARzqsrL4CuZo833HTWZy5TJTecFbjyfUhQhlREPPYCwOSajRO9I+zGyHsBlwzTfnT
YGerwHas4EUvJAfEyah6JpD33aEhJi0n0zWv8mjS6BlyI7PJgouQbAkTXh8Ok+oWtj2zB/lp2+oX
gYtjwr9JmcCZiC1dQd62lIVthVcsqQmWWnf1G7bfVTRbn24vCHUZoRlJjX+y8a7rdnzury4b5pGm
CPsxpk7/wCCsK9Ehj6e99nGmye634CVpt3JUmmtMVGQ37ueuIkJ9AbdahI01O8TwF8A4OVxMeH+9
Kp/lR59mTzGX5hzOziEZ1MZAaenGE+S6tx50V0fnPECLavqDFyZYMEdr6qIDLyFRwbfPgk0lMOjK
p6ND31JMUueJJUdpr21L0FDWJB+wGdQmjhH1dpoGqQxew+hVIWOXPbqTKqFXizxeZEuuXeUh7SOP
Ndos4W1u/zqiqRxLyz60z/UMkPeuW/ZnmDVlKjkLX+yRe8wasmsx1VYXeUIaCrhIaOePmP2HwhoK
p0rwJvU/i+ZA1YvWppGfO3cZew6XBB9khkN63HdfCwpujdK1idFOJg/FLSMNuKxg9C4a0Kz1rJtj
EUIdZ1go8Ke4Awrf+uqqJ2vRj/hMjBsJz0L96vNCFo5UpHC8XBd3OBl7tXKsSby1rWxmLjGNGHSw
p5EDPZUomyh/AI2T+JBSoqIysw37Wer6bBHFgrh9Av1Nc5O3fjIU5CBsgBMGny9crf7Q9jxA8MvC
dACKj/wJQ8yf9oiRsD+PZDUI9wTaSFY7wIB8k16/cKzQd3SfJz1Mvt0CEwyvxsIaf+NbaoGA7lvn
a29CZSgV4b/OsePdY6O0qCrJ63IfiY1a9I2X9VXkzqFMqrusLNrMjuJ2qP26xPIJPJ/xbHcLv+97
W+AmnbJ0fc5qMaM7bKPFdJJLQdqF4cmwTaSaNQQ74hqEAdHoqF4IgG+u9QFc1pnffr+bNv1JMD8N
X7tFd1aQl0rguQH7DgK0S3MIZou3hHc+8l1CXAZVGs61ekpO2TuSYHEYlfLdy2m5zZdjrswDIPPc
V1krp4MeNU6A57fE8ufJ0nyw/SO9x7T461xhN2T8kyt0kNXTjllUR1JFH6BWZybhK1aHtLwtYGOD
hUyx+TJyCjyvlWQWHbidZrlcWC78WQvj4k1ngZ/ALmqh4A2x6NcRhNHy9wcI7QBsQhdqFBQalUSH
wByU3NtD2ZRvW6VWFeBiD1yTZ7RzuvUP7b3RXGuhckyd90c3FlQO+dGlTIfLZv4HWlZYDsAGpC6T
iWDtwTNnf/4kv4BiYr/iCH/RM2XlOxB39a+HINiKymx07GkXBwka0sm2GguByQHlUjmp9v7D2kyO
7r39gCyDUMl+cpt3CrjulTZ+Eu5/n6NsoBz2cgQ8jGwuGlGXQP97gjh7rHTF/jLSQifkjcf2ekw4
ePv6ZSNIM9An5OUktkecIEy2Arkv0ud1BtX+EQJy9W+HC2/w0IYFHyrZrRpY7h12CWsCqvue8Bpz
SZZoLwU2wnx8epgaIc7YdHGt6btLddWGf5YYcLjqW/btmK9QgVDUnv4DkVqUXdj6h/aIXTpioz1R
HSt6ZRowuv11VFV0NfRoJkQDJNKq5V6JjhQF+5Trq3Q9MklervmNkMQLk9pk8r4lcKcw7L/ef6/j
Jt6WlQyXT1tFeaG8HK0270IXqJIlvXLU/gkJmkzZPWKGRd9zDLZkWlQKkSoWv/aYZu4y2TRIC1pA
kJo16lh3gJAYIg4RYUER3zzi5NzUUg8BCeG0cGLN/CsJu+doj2WIPZmIkBHwf3nWnSqqI/xsu9Uw
FxrH9jWhP+EqJzJoZdUcbDZzXCwAz+5B4M9si9KPHO6KSURvcHXvjgvkdhvMRyi7BrtUyC82q17d
0DT7BWGV910jnEq2YfGbV7V4qowRyE74RzPE9S8l1FD6T6TKaxrjhg9rNu53acGk27OTn3fq6rdi
VBITyha1bwaEQM9jJP0+X0ipnzlVv8zCj8jCB/jgyZxUa2G+etFwCjei8BMYq+wCZvifg949j0Pj
uUosILGY8xef/m6XDFHM0Z0zwWDfbK3QDg3VpCeU+mM14+DuFBngvGmvudYTiEKFqCML33z2D78M
+gFqAiY4sw5Ocpz02fELCf7Gv36q4cZdgHpqivflWvejsFp1zOh2nWxR66ugq+/1fXs77slN97Pi
49tQ/5+qHbz7vS2zU2HekElT4AefoWTNYJjfVGZuPzAFjx/u1h4/vN9+iMl1qoFU+yjjgGKRZbgw
qTKA1ddBMPxpesLw2D+OeLyGcxzAgP4+EwtmXmrstbcoD/+cWIwibwNN3lzTaElCHwCSFMnEab2n
Lg+3oIrdslvERnI41zzv8yvrh7l7+CHnIrQ8Rek8KuP4j2ssul4vdJPSFWVy+S430FirrmA5/xnV
vtYSlV94LCIEXu3LOA/7IuOn5k2WKUCV9zjZ+FJWAVppedzSvooQshiC2+sTo9QvVF3SvOmlpBlB
rc5+dZwlOLloEgyBMaC7hBxiVgecl2z/oF/Q5lM1ihHm9MccstrsZREIdGLcAV0iOPeOqV7qJV/V
m/t1w0fEnN1e6+GYYEb6Ig1to58gmoz+smLTeI3BEmF4XsW/KNdL7ZDWvWFxI3Q7MzM61ZZN/gcz
39UusmNAyyu3eHyf959Qdd5LMxeGa3Aj2FUL9o8G3qFcTxrXcjOATWeZOSuf4Co8WEO8eS1fQl0N
Apoe3zsv3qfnC/rZrkojbXG25Gxs/I3eUQS4gGv2gvx8Csg2TDvZvVR8KAxPJL4EroUBy3uKLwtz
MzsLtQp81QJGhiaWg0uEmhQrIfQv+P5BnFp4LCncQnE+lDGu8GBtZLbH5Bx1RGXSOaibLHLyb4Ec
p7diOaMTXMsgjsWB3rw0U3cSQfbDRv83xZtDFoEBECw2OBNwcbDl9lcDxlDrO7oYdCttfG0Y6xnD
TLGUO9Q0toi/NF8aV/76nM9egtp7VGaFBxaBe0Aw/kqrpCm1W8yYoGrrRVMsfKjI9soqrnLwvTcj
Xj+E1GPifDzqforVzm3/+LhSMDpyIJmaKYnRv9QpvefT+aqddpgPg/Z5kZggA/KLeNy99XD34fAh
07eF87DrMVLGPt8TkjedwM59axz32Gg+qUetbpuc0J7TLTqMzwugjmX0zpw9YtxF/Plvmz7dj9Hc
HB8h6sQfmlc07mqBgwBKaQgh2pQ8hPUuOhf1D6PielsedttMCUTjGTX23kDQNkqeuaGP220GTxTy
0qJDWcvvjyyQibsIOd4vehpLL0mPMfTX0mGsXHV49R0Qj7sqqHmh7oYRVrTahreCywlMEITiB8Sc
JSLgrE1/3okI84gRuTYckLC09oIi79wLSt146NcZiUeehIbv8yhZGSO7lc+CJLM4yi86TR71021+
rBNIAWf5ImKLaaOZNtbo5hUBpp0AdFVW0NLtgO1FAeNGbc3mos9jU1IvQqdrfGAOCNMzcsw3asXD
uuFTAjb6h5jkZ6CoycQO/PLI3LerF3fLgMhq0YYDPLgnz2yumLob3eQ9LIyelJqdHGqQm6lNfOE0
NOlYQnAqlvD+J0Kncy7tsFNslD/cG2QSWF9MoAyf3ZEhRlFwVPDd70zrwtc9UEktKLsqOVdvXGCo
y6JgCskwpcCK1lfY6IMFTegH3lfswCuSAsVbTtY4/hrJt4v+w5gtUxm3yD5ldYqRV8qcy6MKMDht
lu1uCwrjNywh5IczM5epTfMPN7AgXEJ1twRZpkYBr6A7BrCEwcPTh9mTFftEvY2hs+K1fyjrlSQi
pvE6NDwyrtcCtaOfr0aET0rwoNfRqMVoISk1ee43UYiiNW3qq6IaoN/U1KqZoLsJalo9NCO+WzAk
UL7ozBoTiIUBmW0wVUUqQ21yiCRWitlfpmpjXI/z4SEK+L/l+OBHSdAVa8mO5U49l2qgf76xMqGr
u6z9Q7yGka/UhwK9rrwea6qe3FCPt9syW+gyPU7kUDTptriQtR+jPIRqUa/AJ8zzVIA3zyyjwRnQ
2FC2Foz2bgOtupPjPfPcLSyVSWETPpxLHioNNzKrK6cT7kPQFIr6OmZ8Uo22srU2D1e2o743g0Oh
tpzLBzLp7pViTn7vQpZVxoEV0NYdzSop3wQjHeTj9My8+G/gMQumcNOJV6s6wDzBp0sbv6QjT9yf
Jf8CRKfqXU/r+qFb3FZq0wXXPsR8Ak7RDt0aGEruoSthrdnPb/EjcwaqdpU5uTVCEmfHdMfx3M4/
ylyev0nJ+VoCkpw1MR/d3jmDBsqHhZuixfcwJ/GUqTIiTeWForwdR5KEnOb2UrW65SKdoPEseobE
DiHnv7LBcRnTvdGEb+mZMBgfzoVztwuP/LWt7Id0Wa57ZRcpD0ykwFJ2JWzRYw7vS4FmZD4nsyaJ
xDV9TQPc3ZuWAu1uwpnZTqGJqNfLIXh86rKuTBlj6czuN08EcX6945FWF+RPuZ8vlYlbv9YWz6Em
rFkha6cmkXiKlYRcghldOMFEGw0/sE85vj0wtXlFLa3HCxl+M+1AIhdaGsxpD8WaQYKAxNGYKMAl
UdGcAWUrx0ykIeJ6K8CRJx5tLLR8fwkHNBcmNPOEOVRwIJeAyBLu75CC/ljX400z3A7uk7JIaGsw
mU0k1ANe1H0UC6zmxmr/2siWRpljGnBKbv/jZn9hSUCB0lzOE+/4ozLh6dXDnZDZwPFjzthpx7Xn
YB/W7wtkIzpXwXVUPO7BR3y6FG8QckoyXZvXR4Tfe6dZ/wtErfiytozkFA1dLev2Ds8i6qSYrsPE
y9ZrqAEaM2HyQWH7OXiiDR7WBjeFgbzROQg2lIPdHtxFQ80ecCJ3hcLJMRa4q1MRacisWNWuuJ3r
ik9SGwSd0FE3C18Jl7VPDgzOoxARF8qFw3eJOAchiW8rj4gq3Vm2F0W7pBgMdJd42lv9CLsjKOAC
I1Cb+5Ja9an0Gw9xd+EePaIFahsbwHNXdxnEEzjsUwpBIshTzEv/eR32l4kOdjiF8X1H1SkdnhsU
ayBH0bYb9ssqPgPtdVBJVo2GbMMFMSiSOMUCTEe+IN2l1+7Se5l+Z6zTKs2DL+eWZlJ3exHoBk20
38pqdcwaw+6CeKnwJzubIE5fsN3tIFWMr7gmzmI6p+Ix5PoVxfxc78gvprUB7WxWmGVzlmyOt+4D
NTG3ntdycKyvMhWKlBAWfXwlPEP6yga22+T6WxPCwC8ptFzRazSwvHJF5jPWJ+8Po+doqvriwa7x
Hh3KbKZ1BPfAY/ftk8R0hUJAMIE4ns94GGCoC8gbmw0hDMmkOOnBuY6pV6X7+sbR+rCvOnU0p1e7
AscxuzZSTsLTyejdL8nqPyABUhvcGGO1PvlJrXH+YLcCfx2fILnKVecypPvXnUA+Tp47u7idFpkq
HGLQpJqpHwl7IW84MroYimJ41apHVBpT2Y+sVTSYrVkFJ/qNkVujdrbaASWVIJj8h/O4aXntjLYx
E5DT/ENNWOdwx9FXrVPeVi1yfDAIfW3/x3lIlYeQWSILVnVYvApbDKMswsotTS/728IIk/4riQxX
qhMZNNQRYBNNsybvyGUHDOQAHOBCrWb3neY7yJ6y5ghKAhbe/1oziWTcUlsyVOVC7tl4eXeqqpqi
Db/XdEg4Lk8V/8KRC3nkTLoZy1uAbFmXTvSj7LiJfGmArydRsRGzIhPdVqCHGSO/CFiKQ2cOgNbk
uqnxYbG0qHd2L6KhtfS8ak1/LlzvF7z7XkVqDCoaUg2Y3vxKacTQwI7AFhxU7pfvf47r3Y0xjhsA
UJfNy5Qty19aRQD9GtMPluYeFO0zXLSXKKbGy1HqSoR9D/DWGdV/EerlbEX7CFraq/BDyj7DsADQ
ye219mY52t37xk5vXrmTWr4XYssfQDFclg0MQhQ8v6WLbqNyZvjxwTRuqVraiKGN+N+m0tR6FjuV
8Ln9hUlbo28hpC9KtSsarVaWOSWaf0jQDsGw7Io7orkVImizMi4tFkhd33C2myZby108ZxZgtkka
TOERNU6eSVp8Gk5jKUMqqAHuU+m4V6aq8Lh4gKn2sQiFrcMPM+fvvQRLur0AaAMPxLEmSg4rTPYP
8jG6w8sWsC7Evoa3Hjlej8mqkd054SIPUhNxXBxHJ92r9NYiDkEL0tv5oXNXU70EAbHmBTtNeOZM
6qUFBrgwIZk9wXj9WAIN/Z4PkxwLIemU4P9S6NH3gMn9mHsfcqPYHIwwm9cE1VZjyw7blO7v92L9
xdqrdATxAqCsNf9XLZJj2/hGdbaMCgmcOtEwjlofUcci5kiY2DEYUsFqiovWmufj5y0K33n8Q467
SPbKHAsrRJDQub+OVRH26IyCN9NaTeW1h40NG7wB7780bYPErtX3KmXKndb3LGqGddXCPNaEtLp2
6rg4vrPAgRsy9M9pVuItdF9sl8jo082KvxLix07nW6BAjmg2Ha74ZYQ4oZxJ/BtPU1d8QNFJR48Z
pJxyvyrdPUbFxJSQOHoKfR5DyNoB0PIlpYHnuoPocX932VuTbiK6cgvO4CP57LmblgK3LHNUD/do
h5eDhYcAxAiVcemtTQEykkr+fub1rygy9GkRQbfJbSa3uZp08miBdIwlvk4pGMkdvLz869zFz507
EEXajVkUnAFUU4gQEHewOngll3IaukuLOWTUONQ23mVvPcQfgs8M15ebU9pvpArwLkTMSzNjT/SS
Kyu1aWMMW5ie6HauwjDrIrrIkYiZlF/BbPFPTl8rIQd18W+MDygUtOC+ZRzkZCI17xP4D/32Tf9T
Jb59d9i3L7GREES56mhLUSFWi+3KaSMwQK4jVMi0yUSe9oeDMeds6QCwE7LKdPymFkAjOUwOtVY/
1i4rkHLwSo0k2g8JgCEuZq749iajCnJh6SXy9bsBvLWE8vTD+JK5T6AHLlDQsRuYcyc4V6skKVLC
AucdWRbVMx0rI9DYY5vAkT7zDdHFEsK89Ep8vI2AaQ5yThEBTJXfYaswAN2qp7cbB3GWQZYCVarb
VMpL2DOWtgefmhYzOlsAMdVVLwg2LavbddOCsj/eXuTZB3xX8El+5E683i90RiGFsi91KXKJ3v0X
cV+S8gnzSujeUsShREFN5tHhUsq7itdUPn6czKG11mINTfAEblkd8+y7uAiM74CBVbgMoF25uqx5
O/MXabvKMJZagtAB9Hjy135iOO+HxAvZ929JbBK+7yjETvMaAQmvtQssMG30MQp7zs6kFVerAzqO
HpiqjIdaoYJn3OL5wU+NTJi5ggXkmD9Wq52Wdp4TrQ8vlgzGeJpZJH7O+JUS3rgUf3ghMfcJ/O18
lavvxzCrnyLtoIjByM11FV9N/aeohWvvtMM2P6WGHYcmKkcjlkjE+Sec+Q37qJN00H8RP+lBRubz
RNg3c6Vp5wJSq4Af9+V4YTw+6wPblJm145YkTP+h+d96+uodDrfz9v4BiWP8ZDtQc6tmeUUkB/mc
/LaWMOiVwxTHpfavUXbsGFNormNicNBwU5ulVM3iZAky2UAQlUUBZbZkGVH2XtN/MQYfG3p8OKUG
fRWAOZ/ylJpfQ8xFMIYV7v2vXdmxW/izzrkqGfBp1HQ+kCtvwrLjX/gln2ixhRbn+Vh30hRLsBAl
neYs0uC2wB4BZ1YggiiGsViuhmREtfrOiZCzJyoIKqAHsNLamfMHs8z2gWy/MCKWVoD0ZVP4EvtK
WfBe643wnFgotLl24YciDLfYPM4HTmiYlnsm1ApePoqjwfkv6i35JRWfyaiajRLxJHyhvp2atFiJ
Lax30f5fH/C5amsmVczbHAVLdzgSmCltnUax3xpQbVD4yy80ef+7kb619El2v47q312ozsTsRpqB
80ExQtGz7iD5TaVeJyA/Xy7/U+10srO1Zsn/o2rSlNoI0xTYm79i582R3O9AzT+EGX1Hwk3y0UHv
l6JzX3XMrkw/+ZDwB9NTTTRsywUyrjlGrG5JVQKtnpWtJKCUUeSny67s4tws/ySwWUpkJX/VrIEB
31EvyZt41IBvZ4WsMxVkcMS042P8HHcZqfFFn8H/Sj8JZNST/+7QGOTJZiVlamw5ZBk9/gB5Qyo0
j3ypaWiIt1x5GwBcvl58ntHcJXXCO7eMU1HN/80G03uaVOiwJ+GXcQ/YYVeAScALQ9FxOCxR6if3
PFTCfvLW8F/lizlVKC42CPFCwJ96Gcwt7U+lnshEjr1oaFWlUuOBpqpoyNM7TwXDtjyvSF5Zy3jl
o6ikZPf58VX14lF8w/WiX7FRS95AObBjmmM5WLpaG1MeVeWEkc5qmJe1FbtEuh9TJk9RSJhpq4hL
DZOyifp/JrS48qYhyPX9xxtDUzc/7MJxs8X99RJTo1yaHMyZrATlSKBkYC6sS9ycBZQRgzQGCR9u
G+mj/nlJcCd0m7/TjfkZZfn+RNlw0z8AMkOtQXq0crGw0aCEZx5ULDK7Efxs7s/rP2ZG1tfj3DmJ
SmhCuf/aHD/FHZTnIRl4XTi8al/Q2B0sD8aJtkINu91JP+ksEIWNCZlE1hyaNllcvxVmQTwgTu5d
xlgnWDf3zv9+Q3uZ39iFFmFrgYO3kwXBV8SWPna+jX2TOYheo6EENeTRUJB/ZSenq+bRqJk+fLpP
D9ZifFxxuDy5N3csWqSriiPFgJ+UhTVo0wNeMOOauKQWw99AYVBsCklZj0Iv/Qzti0ENxZ1m7W1f
zHtkwrap2g/lKyVgdfRsMdXqF4FLdRtFkt1TNBJ7xSyoSvuTjMZ6aGcbaNoNAFmOyzWx1yIikPsB
HPRtcqRNZmgZ/6BXpzH0P84pfIQxJBXew+Y30IPTHA2d36cYpPQF6W94DSiHfM4PQP7aiauLSRmE
ld+84veVz0K1EYkn4Kst6L6+q5k8VJ3vBjjGiu25av8zNbCo1Byw7qGrFDnuO3l5Z4Fagaew6u8x
YdUTUOKVoFhFs5XGLPeSby96MD2CUEC4Wakc1KueGAM6NenYP5mDvX3fBJvSZ2nHv9PZ1ZNOeV0G
PehHfvRC4B6hPHyZgWUKlr+FhzTvz+oPXEjiLZrMGm4G4Oxl8C+a8wBKPvPqDHWRjSqAKJZQhqf9
5Y260Dz/1tUwL2sxn4LneS5H/rz6Lc/WfY6RgSPU1B8zP4mXerrsaKz7vKx4QQmxdrbACX14ntGm
BmDfYiqRXp9rtkbVl2FrCTuJwJhpBNbV4QAto1VlT4ABYeeFa3QRgtb0ud4LcidD0syX7sYmalki
icsZYRrQ0TAV0ILa9uV/UAylC3UB2tQ2Q/ZldZW601ITbRU2evo6Bh8zvo5IZWlFCxfHlhLzeD8D
zE8awCAoDZddF6EGhbphIvfAbkOarLs4QhYmShHxnkYcT12xqNTCCAchcvd/4G6oHfabIVIw9qv7
9K3p1OlF978VJIL1OvyrROg6wCGR9+MZRiN91VV0TjdEUJ0BIyRzzSS/tC6GbT/8elK55OeU7sV1
f2UhPSw0LTNBSLBbdv4MT6V4Mmt0oMHyXlLV/k2akNvDzLDvWXEq+dyTMKL15jdqlZVbynWOil/V
sRNz4YfmN5XJ44KnGrSrmt0EATPuXCOxmib9CU12R9dhkVen2s1lJI8BZErv50vAKRm8cN3jhCD7
fa8XyX8qtIQTSdrQzjHl+Lm3QAvp32kSm+uYpeQALv+8g3Qbrib62d3FRZbh0Er9qSPIdZy2vPfg
fwS2qAoANt+H2WirARH8KGWbt1VtNlj1RbBgMscJgjXnEB8ayr8wMgAqb7iEr3sewUJUqL9YuRhG
GbvMUk5ylLkZd5GZZpuIsh1EYsLq/iOmT1P6JuMzvaTY6z1jcltwO8IbRFyuEU2qFLflfSv0voqj
Fqoa1bG0Sy5QLPoBvfU57hnM3075FSa9PC6RNtuFRUQMxonta5dEIWADlY0sb5/6B/VN0uriDvBf
vcm1VZDKZT4aIFDjH0wfwTgy9xME1fnqUxAR6uieza9r/MYsP/WAjweWr8D1r9M0x16oO1GdM0rp
5RPAtvtmb+grniNH6AMXKAWba/jmWNO2H8eOSrsBOfXwvsK9DzXnveXTRKupclPte1+8BUCErJzn
rRV6aSG9HK557D95IwbkYG/UB143yxTQ1auqHjoNxKWpNxS6++QQ0SvajpAQ1rl0ajz7j/rE893N
EDmB0HBPJnMVrBw2Hw7e+Xds32SzzeN4Qvd6iqQW0foL2pOZGwdmDk8+gvPp/wBNOA+usTmooIsC
hcQp77Af+lHz+CmA10eIb6nHI3vq1Nuya8P1JyyO9cqj+hmy/0+R6yao81XNNgRIFOeKuIXf420O
35wQwU4kpQT345v7i9Fl7yql+ldbbxEa3O+PBoTXl+5/HrJHTYXNiJ9AkVPKtO4D9u5d+S/UramI
+t3RVhreV+d3rMAqjbrD8z3+P1XSqWRbWcbFzexln4yykVXPCGrAbxQNgTsTiuL2EnEpos0JjHI1
dvncO6YLhNtquJAZtWzMTMVWwZ/RPDXS4kP9nP0SpFflU9IR5NWS7Yafr+Unkm5EQUwymhaBi1ff
rUJuN0V85EovHFG7pEofrgsc1WBQWAtLZK2AkALDvTIlAbloYvzK+awNmOl1VUnrNfDJDROpGqUT
4ugY+dAOJsxJY+osROPNkjO/Ngp/sxSncCceCHbSbbiWHt1/viDgUz/uc9by780GYeFOiIapAwvd
prEKywcFcCIeBlzPitybJGSAxZmpWHbuawNfoT8z6b0r70vM9Uw5ae7wA31TWI3VpacK92Y8xvVb
2v41tCkSOvNW1ze+eklSkYP/oWSx1DRU+GxsKy7CEZuexCUY/+GEEXJ2pSO1ZXi6vpvX2e5gDKqf
xbdfTvGwLf9K3eYuahnf+kGTcIooTqoOqqKWiSe2XxCI0xkhResgsrwalhZyurYSv+tFXs5o7wIP
p12QLP4rWepr0O2oaEguT0/VHTl1SB/tyjtLSCD5adpi0SEPnRsPfGDEUJQtaXMxzF+Vpdby2MRr
StJ6pExwNAr0tEoZX2bQ5oxUh89OKYAl/E2hI3RoF8NqjY+Q27qc51k9mP17erJfJOnUfZF4/yXi
ZMoBxAkai28aS90jAbuwtLInP14cKBs3b/ZcOI06DOf6WSNev1SpQOgAEITfswXjjHvgKe71kJyK
Ce7qJ0yOTGU8YbWUCnu6gxO3NJ9wecCw7IDXskh6YvWfC3NNb3vrdBvRnCcJke7bhcJ4whKkVLyx
7CWe9yeSlKMd88Vjifz7idVZ0dSFUgNykPaX9vEFykrCPQXxMFL+p4FAwmqb4BO5mm44jg+sSf+7
F+AOMO3AliiWhquOyJR4ed7j6cMQTw/4511VkeYNr74V/5jDRV8UgipEc5BTns0B+xDU4608SSXr
I//kGKEY9+nmx0OQ/gE+UP1XosjCbkwRBE08mdSVMfcGEOvM8kfY4oROiJHyeWn5IFW01q4ixbUj
VcPrRF0MCnq18F6BAgi1Eqq3xhBmYLFYNhX0P52noGakpWbWPk8Y/Eq2MwrA6OQAqMZgntKhAF9c
ZBmjRzOA1H8X1w5lYyvQxrQPPiDWKx32jqNhNJScotNsbLzIoMb6fDxmZTBhEgmFi51caRbV0Fuo
6uJLE4Dw8JsSEYDts3BZRDyZqWR3xTar9jzL09A67S0e+eZHqcX9yJp1xQt1lS9nYZ0EWKS51mf6
q/siMzNn1clNB8Xu+Z+Uol9g3Hh4Jp9cVNFsTVe8qmWKbNaBMcxGQte4FXZphEFd112jU6GBDOjH
N0CpqS9Tz4svm73GZ91wdxzqY+q6itejLLVbFtr4KrWuFQkRUW0etO3h7zJ3zuCH8gp+Dn+9KHBn
GjqKKGnuIBSPVNwrPoAetu9iuT3tISkR3gOuRMOlrk3kXM9HKrmL1ydjYDO9EEm8n839rt5J4FkK
Ltxcgd1zj4YgysNLiKKKv3gi89siWxbD+1WxTgPcaPMWdUAZuI4fnyzxSSwEDuCBr4SfMLEoHgqv
EQt3RXCU6aiyooIgdNEJ5oA47Dwk8Xr5G87QIUDQe+Uadwb3ub2GQQ123JJHZet9JCIRiFDgZevM
muFp6X2icXI7qsqBmnmeH7MfGdXjltVdIpwgZ2KEVwfcOhcMG+wuAlcyRLJbAGtwNvFxDcRe1zZB
V0WUDLHYlN/ruZJDFjiU1Vkm6oeey17RDJD/oGufASZXP8K63BsxK+LR+nfG8YNB4MgdQE7nbycm
DRnjtqsTrLcOaRAET1OcvlaeVEjkiVi7LAtzZKAeQdIUdsp060dWvmoY18OPJj8pWbFbQ+9bVVFn
JeOnQkPbrezSXGomFDxBfMIAxKbTS25z+asWwoMUdP1iR7yp1lvw88+qlDrqPDC90jOSqLSNE1gS
sWR4PVAKm52SfrNTIVCB+az3sw/7b2D7+FdexDF36EZ0H5bAkN6jf/wVuFl1znOtjblc8H/K3AZg
Y1e8YgDfwxUz62rZ/LaGs6we4jzIRl/375fBGo3DruqptW8jvg0tSveBlwQ4/Y1GpaH8aMVjik1P
bZIQLq1wM77qp5ZBf+B62DoOQe2PB0TFODSZomeLmZOzpH/JyvdzNUFwg7IJCYo5LX7Fhe2GptB3
/3YIEnl1eC7yZXo3uOeXpNP1C3sFqqN32IHmWiiJ/+hdJ4B8DS43SoAUCkxEFWBveVNkAE9Kpwsm
icoI0+ln7nGVTvIryts31D2MQplpR+NmR3BAteOfMaG00YJMYwUqiPQbVQM2NjcOLOV9x7yFVvJW
vcVtuqY+wTf7adTuQNrr1C6yDrYAOxXlAerhPqJ/YZK5I8eYYSRyqAuzq+DWqEYhxdRBxX67NuHV
pRcq1pmfnRALSAo1L2nl1juvZCNNMuLMrNITmq6eFcKz5mwA3PueSUyFA5YKQg0SYHfcSIeglMt5
hNtFnho1my4WHWNLs7CPnWI43cQMXwmMqw4o6i8UetRyCKMHO0lKkKBlGFtqf4M5DTxBW1kM/ohR
fdN/rYIyBzYk2aGdJRkKHA9mksq6rQzXxZuDI0agCx5VMyuOAm4NvJBvVqJGCM5YJMr2vM9YDXcc
Nlxjh3yEWKXujMsJT6kgH9IWsZZr606gNzSF4dn1UlocsTuJabcAqylIqdkg+TVezhcZezJx0kdp
yzdGmaTgJwiHSjFtfhfQ//NDahwS5Jh9Jpx7wqqoKU82tnLN7kvkEjELtYRBQirfWGEoKAEM0O8q
OOK3HzVsI2sx/AME9Zyv9uFhon1tuBNN28cierSG2Fu3I1hXYxsq3+XQeMNCLWsLGUPoYbg6txb8
5EkTYi/t3qtL1fn71t/1u011rzpXhTg+aM9hfEYH9PtF/wfRSnbSZz0ci5MfZXOOW4zdCYaFHW7v
V+LpaFqnxjzx99Y01dT9wLLzS2rbn7I6X42fX8CMHhLYtHAInYMNYFwrw2qb4q7uXOErUvmrcSLV
O/c8/8QsL40NHmH8pNj//r1ScvDoDn/P0S7w1IlxfzqGl3xy46HPqh0LNeOS7nyOYxhJhQ3UAILd
D385SWkaHVEE3pOCP8avl5wsitx57WaUNS4DxJerwhrmg10nBO2KzkMIy6ZiqQlE95jWEA4oA46x
a+MieNWgqfK6bX7lxkUveocrsD7ZlMuztkft2VkNRI6DpdL9wYZQnpRBz8lc/4UQPnKUaJpwAs51
X7gj1Gwa/GtIImQHoVkYKK1aWhu1ikfj5b4SPFN52Uli+A2yBtJd9NCV7J/G+/omUWJkD41UtyDn
dhINBgxUU8/X3h8odITMR2r2n4aqT5PcGNItvIkjPdhOYNVI2my6cEAsRQ4ETv1AGkQvhMCFvKvZ
oqSZ1DHHcLMGa1MRNbAPAKXzxGuF3zsOzCObBBoPIGw1rTUL7AtJSLj6Ox+7g2naH2x+D4lzAcQl
fUzT44+pCIeozowPsUI77CrLK75TfT/Vm5yw2xVA+4reOFe1SoIDX9uXIFoL23PwJKMBM6GKgTGe
SeE56SQZSTPodofsaL2lXr3qCmACNkXiTmGMuypEqoWBkn9Qq+FIEBWSLZUk0VEJFbDwo565WkJs
KDExoAMEZTDw990vpXUYPalBGG0L1cWvPOhGR2fUQ4pGqYx0ptgw4Dlb0CuJls4plbmSK1rlCqXX
QokOTM41Hh8cSJYqIcXvdoSUfkU2pJuNctl32gvqIDqX7reRXGhDZ15aWb1UX7Fb8+lY6njZZG01
mEUkoqRXd3VHXr8m8jxcgiF+04ji5DknPS/o/WAqZR1jNA2o7uMFYycq65eNQMVsPSiHKo6Owfe/
leILzpLvRCUY1JGC4y6ZNd6ChO4nuKTFFqmBe0+IXMiEBWnxN9nIf9Og6CBOhJQvT0Ru8tG5Pkuq
WEcSP8fOjE4gRqyaGjof/rXmba246tWCNkqxKAVB17PVWb8gXG4lUYw6GARJ/r+pn/7x3Y6bkb78
afGLtrDYobK8aXxhUIXVbKfQz65EhVZdZq9lYWOIHhrAmxqJlGU4xyWBjPtWyIgpFJQ2hyNdnTJT
60Yw4ZRNrGh5WgF1BSuKRa+5dV9bZ2Gk8wH5uemdsm36fbaK+8mWAcnIqejQEbN+FiRdMQ+7I3kH
bnT49TUqxfWZQHPicEJk3/j9RcRDKRHxjQYF/uXtcbAuoUKiYgy2qhvc5VlCE/0OZhlu7pshxx7H
ZwCoqejfDdBqPBXB1/erlPL5tIfD5JaM7N5BNJUcAHkT5bOVRhzwWxp5MGWW5wQJWUxEYZJ8vFpD
FJBZC3334t6FzQ5DhIdwhdfN5suX8XANS6XmaA+sCFMuz8YX/iO3k2gRqj99Q4YivFKe3+5QQiQI
05KWhNdUtchkH7hhQ3k5N2/0s5tyLpHxcC8af8xSUQ98ujiz/Ntj+AJo83RW3ikOGPc7PSTUX1RT
0zlkoYEdpx4Rwv2YreE+uBs51xX9H6j70Tcb0Gccqzvv8bhyne491Ue+IqzPJSoALSFRGg+DWNY3
1NzOveUTeGrop5K5xOSdI61hhpjAibk6nfml2Y4nI08Css33q10eS48sxNX3xtu5ZbvHx5w7P8oh
HwBaaPwV3vbnb8Gk8QWJmeOC9pVl5yCYgqpv0k2FuWJoTHQKOq5y7pMtC+YATs3Br9l70+AHLOyW
V5X4HHaQ+U+QmCz4et+aYw9kIR88fuAl/txi/bwlB83MKhDnoO2znySOggZO5nhOmZsLNplaIIOY
A49TkpZWXEyQC4i3SFqMQT27yr2A3aFGYjEpPoboHl9CiBFS30+9inRvriEvh5gUUpRy96DneTE7
bv9Pc3FiNllfM5MTCMfvw0N6Yn4OY7cU4UFHmF+3S+mOmSedIrIDjVLHPu/XZNpBKiNT3S79v+X6
qykUNIomUqLeYRGhu00ckq1/gvuWVCtT6kMvYqdRyKXccSj2CKmC8K5Cd1BHcDjB2Cr82Y3NAV6I
sP4f26hgg1RnYNUQXcnhHokV8mqKcptEsodBNO0hCEg/4gX2ql+MzZQAM1+tA180VlLPkLcH2/ZZ
A8W/gi1tqZk2VBxFttfn6yF8huxlmTrGe1KrNOZ1awXttVqxyp0+Y5+7vFGYZ/sdNeGS8ihhQV7M
Nf3f+6Bh48He8h34nbvquL5umJ2OWenPYg0HbT7Bu7ial6M21+dFD5GYJ2xA4Qxa2NopS9dAfQPR
/weU2hQ+ogYih6zBhpL1YO+9PnS6DNS3q2eniYV/7ih4UNEdZOTgudBa4ChaRg/jt94FWSWiFDll
96HJ46SqUR4T7CUh0iXcBm+3bZoeBn4Y4hCL29frPyY8fMmlQsnx3S7QVoCGqmOu6PuGqQoq/fqS
Dh7e+CgOVFfIaJe840BvJnx6Aj9ChYjF5g0CUejhYvHBRPX/74OmrtSjeqXEMxWXqitl962wTdWZ
0K9gSq+aMfmRTO03w+DY3YPmJ6eRtDAt1rOxuzkaBkbQ6sF0njGXqxC9INig9WGC4wa/s+YjVrIZ
wxye/2oXK/1xIY3XHGFlVLHVyNQrDhzGipr62CiACEY8OsDshXvmiPirZ/Pvsr9z3IGWtT4sMp00
4v+x8ksjYSYtD8IfPfoO5v25FjS4E5Lvbo25N+E/IVnvR5u1gi1PS4tn6W0e46dsDua9pXz5BByL
sMzCL/0j8ux8sVuBxn4S1Vfclzj5pmxdqX033ZCcldrFJCPcWVd1FiyRIx9shoKc7op3P067GA+E
pbDfGFGnEHN9NXH2v4NeCklT1WpTR7oXcTg5T4gNXoFT2lXumadTwOP0kyRPpmuWWa6Osbo0CFw3
kS2rO6He5eTUf3nEocOJ2uEXk2Vhhvl7IVWOPfVjGHHq21TQAmHVvzD2kH0fsCc81ulYuTycgnHA
Ua/Gf7j0+Jr6/Y2nqW9BX47Of0vdsPL9AWL3Imi76HrDqCUe06i1+za8KCN8p2BVbRp7dgGrkwjn
pJqEM9NNwrPIcI90E2dl7an/7gCg0JJl8RUYtsG6sKx1wtrl4LmYfxwnDS1RVG3YW/4SD3vEdu22
Ds5nkE5c3wLmbZkzZFSM3ug46VJYAh2rLia/XlglhHhbNigo0MtBJKYO0B3VCVO0MC1Y8vVBTba5
uJng8d9eZc9hr5VVYE54EVJbLOcLyS57CS/FWANSPeSZDN1XN3k98q6w0Uy1f8iE1tGK/6wU+UVU
ABGOT95Ygsw+VqRqT6LQlQsmhllyadWESWoWBoxqGJZ6Rz8ucfy/I18DpYTlWWLF4auVWSjNtQT0
XHXd9y2Q2VWVMaj82IJv0xxgercaWWCREPSQ53YSw/MqBmSJqyFC+IR6rDnuZwfMebdWlj3zzLrg
u9CLg1UIqAZ1dKtHubAQkyq2YnNrHQ4a2SBQCTHSGq23k2ivvZSoc1epLbuoXajmxtSx0udV9o63
mb5M013d7ff4Z2VNL+5H4JL8fwqr7KHC4PJgAYsnXdSunX7iIQmizJVJXiQtTfP0P1RXkTfz5geE
cbJDkweidq8N6zHFqHVKWMqZjuGcUuDhdeE07lKxpo6huwZW1HjXAVsoRpngnS5HssyJis0FCEGw
SRayK8obI4DD3eGWwXF/zruQbUSXJD+JOMdI8HVyYVviveMULH1k1JHIKBAp01DYeOpn9sZKROu7
3eUe8lGhEB2KIChjBWJRD6Z9Jxn1f7jhvVAG84Cee9xYONTjFQ6LZgKXPnNb+bBwaI8TonHgZ6Od
Qd9AgYeQ9FyUcLfMU8puJl65rosMuMzS8Ju2mO6yqK7Gg5YjSr+Ihzc3+frh4i/ozscPthnICfmk
yq8kylzw+3GADTXfnuQRcIIMkpXYdC9aGPQpqjalTQc1y8QpLTWk0nml36aofEZSfzULqTZhizyy
ifzwCxwGESCFptcHSJ7P34RkKwlDJ9ht8DYgF9nxlT3RZiXpxW00XdOSVbYiABvSOb5bRPErJJec
ebPhcr6U17LjuRQ6zVaejujjvFeYqK5/tD7aTUVDEQOo59g0DodPhXHU9iVYMtsFXjhV9VQhq7Py
t1Uj1F8r7TqH5T2YQLhp80GopnDEmzwbAUuVn86M7Lsu7oNafZ9xopwA33W4NBdVm8+aEAW5Myv+
rYLOa/ZO9AtD9M8neXjDE5QNTrtZ051MrHApjhSlK7KoImT0mVqwlMQ+KeAVPjE3HC/7NLj4y5fS
gjhf3EllEuOOXi9GyuM1Oy5uw+lNmRhShCdeXgWx/v4m37z2Osu6nSC71KhLXT6laPyTgyUYFJam
o83w+4hTN/Yzx1uOypt3oPwBu7hCBFCCa5Y4XxkimsTLdTzYqQvSv7UhlA9Puzg2geoRJSXuGW6q
fsVnNVdGYeySymzBz24pJ2yUTSjh1LgeuICbHkF/MX5WjbwPTJUkilheTsAjUTn8SvRBg7nX9tl9
hvMKUPfZtL+aji5QpoqqCHy6/9EQe7G5YDpJKKHnxxvLxdE1052oj0CJE6ahH8Ai5wrrHf+sd7JT
Rs3vCno9Eh3LM9DK8YueAOrkjVmewGMZvNLfL8EWwp9mi3setZFS/CFxHCZVDHbjlZ8iZrp4BzIX
yGHoaMVms+Sc76RtXlsPOfRIRLMvKKcg6XbG13SiJyfvKiyiU7mig5uBKG4h0xbScvge1MVx/izG
byBCqfUgnUEo+GA0yrsRC1A9HeQ1dWIP+YrM0ABYV6GP1ad8FRI7duq6SZEB45Pny0OjDqDZh4ZI
ax+P0CCGldtsy7G+reWX4WCvlXI2tb/CEozY7UzfiiYlW26fVmwBFPJSCdQfsqvzjBi7DgL3kl8+
LmfQWl155eKBu2d4Fe+RmONZp62x2RmMg6P3YPUJxfpIzxdZyNWBjsLB8B6Lxbi8NSBm8LWl1wO4
qkwTSAd/KqZydxO2a5XBdSamp9XAJJ3TQdyiAtPjlrMmuS4Cnf6A6C1fVjaxFAP6TBFS2I484viz
m+QTFjviWqB5fAX2MoB6vD98grGTEibiyv6ADpbW8+TqEUPr+o9T7hoMrobazpzNxRkH1DTdfqMn
nnd2OnnHrQhld30tZ22F1D0lsU5jDADTGXEErZrpVaR7nAewiWQYIqYOoEcIS+2KdKElY7oeWZNq
g0PXXUrhtgJQeWlJ2rMYgcmAwFEeBXhaDIkU7biIGtpKIUVYf8G4eCtFHGCEcIAkT6YpS/0FCzR3
NB+1eZmp48EIdjC1GoMdzY0yxsCpMoCPGjxTUe5uqeI+f8Gil1bGoV8HsFJSfYGPMDBiH0bvljjR
zyWwMqb1fbOxjSNVA6J1MSLI5zlLvU2ZuaXTJZryfiKDS7NkJpRmC+f5xu3ANm3k+SHG7yfMeH39
CtchQ7XvkHpi4zp1SoFM9IYdJar3MNR/fxQ1Fs3JXQMYm2NwDeYwWiC0YEJQGF8ZYm+ZDD32Xve3
LPiuIcIZYkh9daTbMCopY3Y/0cwRtrhQBPpFSOMh2sy2X3F1v0E+l2sRMb9EXpTPjAAKtmkhCnNc
vol+COr4SVR7rrT4AAhTZQR+mRIG1ce39bXxS53GgQZw0pBe4egFW2420fqp6EYD6jB7VA9Hcx4+
Ku1H3lD0I74J13JAOxvFy5d2Mx+/iBvm5ivKUQLKQk7xt1hi+UayB8PS9+Qp6UKPAIuP8mNBjfvU
X770a0CT8G66GAX7iXivr5lrmm1wvI6FSoh09JdnL0EYVcUtF02BQI6MRxA+2zUpKPn4PbKSsQvs
BnIyNBDKo9ehZWYdBUJ0S2y/9X/wKFXkS0UXmuVY+7Plc9rheI3FHlQUF3TeO19HkKxLxj5zAluB
WMpgN+gFVbWnu7SHxHfFaY8Kse4PxhpMi4GGQuvwRZ6O8BSZJJLBGLt5mZevbg7aa+/W9XjhpyXM
wJafir/uQ+9ii3LEQs2fNO/GGPOD/AZSGUdIXAEFUZZMvbvUwvXLl1DuiyxIsI7mZUINqEiQERkJ
o8Lym/pZOum1pOT+sJIi8ITMqTg6HftavrmJ2KiUslkb2qJ1CYVPU4oaqVdxb8P6UBlmXj3FQpZJ
5IdM6I6UuwGAMn57eipaVC8Dl+RDCL9s2PhpQe4+a7gg+edEld9slC+XkQiqA9Lafq8OxlXxzps4
BNtYhlMYZiWEunYS6TtUVMuVG6wvr3DPhmZHE6sF8idtmUXZM0lIOiEWSYCNJPgSdNZx6ozMJdsb
NiD1c1rrHR26619cZ4uEmbgwZUPvglhBixBtOynv9sWeiksv45cZf86dvIMjjiRROo1bxYjWYzS8
4GuaqrejeDW7MFDu5M9M2C8fn4Ii1mjO29/q50MiJgQAcoWRFgWZZ4rkuntjP13HN6FD2YazWyZL
/OjOCy89SpoTZmaRZnV61EkFifRiGSNjnViAaVQBOHbfblmeCe8eRL88SWfbV8ldkEMU/ouhiPVz
cnqqvVv9fHXNnB1Sb+nF+nrJl6nNa4IvaHRG4rb7Js4xqjB7jM8XRFujR6ftKfdrUx0ABsMmbQkH
RC9aLyBkNw76gqXbO1wArdQtcQ7T6KE+heeAag5XLymd3EiGcZWEn1zcmKP6T52VEFA9Z76rJKus
fKzQNCQQfsbZYnPvNzFu9aRmTKqggFwfV4g+ph36Ts3q/6Nee1TFO/B938OscJEdrYfHPkc2BZv8
G0lvDcer/U9Qz03yxz9itPipS2Bb1EyHUGW74VXSvOQV5TfreiajzJHHmuAvTRD4wdfGto06XD/7
2w7Oqdmbh2P6SW+O8OCBdUqF3tcO9HyB0nZo2cpEWnoVrSRkWPQkAxmUFic7B8NgjQsleUwP3iD4
jXYyXJAVYrL+e5ne13as5EGXSZ5h2D0oGyOJ3efFuWfRs4LNbe1wXUUUuDrVKkFJNN5jAtWfH4pf
b9c4PsF3kC7z7dCKxFDdIqXOu0d1r2g9D17Po1F1NoetH5YNIXIFR9dmq4ux5PVtDYjD48/c2yz8
4wIxPy+pvSMAIuWSV89uMIUxXQBbPYw4422rfwrjXRl9wjjS+N8IBbSKS5K8vLPRyVuJpYHSYTjg
kKx+RDSs0FDwuDOBl8mqXxFTANqQzxjIB2105gvLvCRh/CQQnYPzHzDjmsfhirTHhVQIY8vcZ8Cy
4lqcj5d1GiJ12nbXt4Vsk9S0YbysJk2vQMcv9wSYgFlUzyBXOZsJvsY4Ra+BojbD6vqrO/sRdGIq
KYQlzEjrmjHl0U9jL25FcsT1EFgpXU91gmFttCnji3ZPYpolOdqjhJKE202X+U+NGmBEIToepCaA
UzuJLwZi/S8IX79ys/V1QeDVuvyqF2JMhYSj3tr070Vq5BqG2Iz9sF7gj/52g/ozbIYyOZXgWOJf
t3riSUcFT1jtiwMRe9XT8xtvFGIGSbEX7iZ2tnZ7I6EYZlatpM7d+q0SWTQTrN3F+qjPZghOqYrS
VzDqiYK9shJzI0jbudOWyPf95adPAeORoCyWSpYy3OJIY2kQzcPdnuaSN0HUpv01et75q5UGhSeD
UrYnmfSB3e33f9K9dbF34f4x7DDPpJHCjhteBFv5WaOTTIqm9gRBfhk4/yRtRBkBdsqmuRcMfifO
xCLShbboqYqJyW7lYBnvjcCPQQY7zj06akBbMennWi+p8sKdNfrG0HnaMaaqHcMVVyDouiUxXmIV
+TpKrAGKnuE0ZrtptqehRy6CTJYJZhjdx86/H+JmChaGFaLz2rcCSz1qQZePPbJr345Q1TygVM/W
cuLwqr85EFehMrF0onsojym/yvZOXgUlEiVu6eETpLoWlyY9wl5VEXVBvoGsshOikNbrw9b2rg6U
oEuQ030d0f7MxoL4RigOY4ff0ghM2YZDF1xgcfZOQnQ8EcvIz2+ZmgEDzhkLN7H9uk6dBN18LRns
kQ0ZyAVH6BbBS24bODi8FmSxT6y8GHU+ZMn2Uor1MYAoPbCPWMHK4Sg5BGuu9uHrntEvfb1PfD2f
7WtCPHsTNaU/K9LCAad51HtHD4J+Ngd1iHjNWgMIAyERZMQKQSG1xT6NUsDOZoxSCW3Y2WxNI6oK
mZGzxdp8oV22kzHj5GDpzDitSPsh1TV+ELKt3IJribu06gEkwxztiNhrLx/367mlXgdxzKQyR1c0
oHS0CtScsGSDimGPmHcMzQ8wRSPpNw0bgncKWiQd+58eRiImXJWwZ6nehHElMzL9yQJ2a/2i/LPV
MDrFrUtlyU+28z/1V8Memotodt4m34fPto4os35Z15mBrRSKmCLul/DVwYUrJXtydvTAXqdqtkBs
iYlMQls9X8reqYoVlqa1Ky6oAPHLEnWHhREeBFwkJryzxIDG11mVxuRCvC9lGSd+nWz5q6kSp6Rh
MLFWrInN2Qy7sfRSNNV5/7U+9N/TF1KlEfmo9Ad0pZN6zYUDNQKKeitl0lyGrbwGCrqXoUZwvLQZ
8sj1adGAGYmAFV1MP4oRGxFJbbdegMNW3hXYPa0vU0lNM/Zlcw5lGzaHV8DaHzexKiCD4MW5wqP5
Q6PGfh4p7ptinH3rMO3CLBRb6eFVEXHEt2KGwjdT47XGfvWfz2aXhPhTmsBhKV6Svi7GKRRVUKaa
1DCy5hK+UI0BOHSSp6+Vb4gt5oe2g/Yfoz5Hhjcz84tvv3aiHWu8tmOD5V3pHa3r7J5Ied8c1wvJ
Zxiybxru/eEhQcPrZtYLbeNYsOfoV9uOtodSV+R511luYlXuAi16v93d30Vr3UqUfKfpDx5vwWrn
6OQAdytJYms17QzdswOWaqpmCVcondPr+mrfjaKuQoFcdTNyXaYdvamiIg/Ce8oPi8YJBKCXo26L
xn3ZpDaPvUl7z+sj305x6LDIvs+5yEDNqI3dCiAaUXkJ/3qF+YipXrrk38FZgsM79b/5KdKr5J/U
KKspqhe0NtOK/RDrFnOj766bJq1Du26+E42mEqFXrZhuQajDYjRV2OnYZEkw8q9dGQMZLpmvMhIT
07tvnhnVh/oS8wXpR30jAWKBhAXCirri5IyEM2PHXGLzlDQjfmujG7Vx+grp9IuhrrsaTVwhHMCx
E4A6fiu8E3EjH9Fs16YicOkACUEgTdAw3J8H+NIQ0r0u87lx9J4oKPLVjZMIvelI3Szi53UkWjFl
FOi3juCyslT7AVn4fWQILqzK0L0FgxaE2yaKa5u3hbLUwIZcSaJfx16w7VyyZbdiPTBv9xWCM9da
RgmSf5UiwlGU5yHepEUOhlmVe3CmhTzZ9rsJCEY492DIj8OdLoCC9vBSwDz2rWRnRnHfagtF6Aes
DvSp+I3Mc5GfzpFs+Z4pNqrZ3MBLL/gpCKVU02KtKGdJDDiTMcbLcXiHHG+ucYSor2hoSbWFU7Mj
w65TV8ajJv8g/2/SSlVUoPkv7/UP1HdSNu1o9Yn7x2R92sM0IcAxxCa+pRuHMqc+9ZSdrk+mZE3R
1dFNXPKJbEbltX9BFqgBl1S2humHrG7UsUdMRVnNTpy3NqhTGIVbeDi0CVQSrpGuV8gCY2PWKUoz
cZFWiMCxIc4j6eHCwIFkeBqluR12oDrIsGHUNDfoUMITcFUdb4fBKTJKNKwH01bFWXpflRSOaFyi
Iv2dR/ZyHwX+AgsjpuVoHsUPD7m2G89luKPyyxf/QKYCeeTp5xw0UUWmnrLzJYzgVWcDQ5cnpWb1
F4zAbcnnApxaDtphuYovgeBYqkOo1Cn9ZkRr5hmImCeg3NqQhAvRg768dfTztzdazXhob5xIm0pi
0Si3/Jb35ugNCZH5zJMcvN3zJQ5zlyCn2hJGHE7Bg09ZQNDLbQECRc+Ffpdlo8DWEL94Y1TlZCEA
eDYh5YfY31+m7hNPcNEXT0jcow8ctITZAWX8HbcDUFPwbGXaCm57aXlzMUjV41qqAQd4kpKGYBD3
C5e5EjbITcOVPW3rbNlmKG47TkKf6zSXrm1mk9gH+2wdorpypcGcFqz/JWR1dWESR2FkBVaMtqbN
455bC3tvkv36NJ9kje+cXLsdIRpfFG9Q7PiYuTEfDU7gLWrf7ZoF6i9qXLsRsJfhtTlqZwIDBx12
hrFylUKFuU1zPKNWi41/UsfZ06KX4yFMY8OMVeWlKKE/4iK0U+aPpuYy7SXaPsu84WMbHt89bVML
KoqCqR1wn/Nk3dt11U6FUdkWPp+whkN4j9rExJNLpKdto5oDyt2jSzfvFx18IPeJPph8Tdn0XtX0
ozh8Aw2KldoYZwsHNzQCbPSQGw6WUq4NXgRtmG7GceWoZ40kRyvwISDZnHhLrbyEWIXkQNlCcuIB
Ng/k+l+qzTrHdYyPA9aAKHkKIRP9TfQDOXC/vVN61z6sF56qDWBffRKMyXdogRH0QzQrXfWZu9Pn
2CBKFmayTAoOOhXznEowV+u1cYvlHEnjvZVcRACZo+ixITKp8HRb5MrwCiYVNSADq1BUD5qvimNS
UPos7wdnqH42WlXxrmjPTe5AX3mAyF0REgxzsESWdUVf7GUf0oUPPl6gnAnjm3TMPDVX9tjpF22g
M1rXfdMXQjWMfKDAcIi5sO62wiq7Yxr+nh4VwxdVhrofTxYgyHTIe2U1vzjRhX447hAto7CtSl/X
/RgsZSsoM+KuIAe6Y0BRf0GnG3hOoJSIjNMoOEg/g/gcLtVr8DlovBBU0pGRx/pKFCFVF06oPZEN
T+PYxlDlTKN7m8RAmvOIO5EsOLfjYcu79oMz5a5msYt1vD6Z6o7uQREx4bNmIbGo1MtUYeqa1buv
R6yNipJzb03Sx+xFkaa+maqtHmlV5cGHc1kpae8RLQuvmF4oMYK5TcGBvxQM8ihCdmnTxM1npurS
NGuFBx/Bm6MeSBa4gQcno0rZxECNuEmwzKTX0PCUVvrguaECJQBNvw83G6gOvOZSsMXqgqHjmrsh
mDbTsMgr8nc40dqFzTMyErUlaDoANJjoL887WMpjwwflNWgY/bkdf2uvKTWTWx2LDXoH/sUhvjoa
cRarUNSb1wTfQVNHUdYrf+EovnaEr+ib90AAT2iwFJpPCIs4hWbjq3fj8dLspYy1W0HvhfaqOQbm
e4pyrpVIuKKZc1MF18w9ZbkiFd+zVAAD/cKqtllpwO6WlmeRvjI2LZEXZHF59ANrfhZfPyX0pRoz
X6lWBZ3sYUJrneCxtfmdJ924FiiUqWMLGvFvtF/JfhzSZclvthMkeazipaCF8hkAoWUT66a/D51B
MHz4lfd9TauJZyTDffoCKjipeSLOBMxrcl19RbPAYC7mHjnQ5ffblX2AC1LcP7NMIliQwWqliGNb
5Gy1RJ1PCYtfLKoJlO99QzRhMVlwsTEKosWt1HgBDo3Br0MA27fYDfvB/d8IJVQa8oov2GH76vxk
A4aPHfqQmQsBa3DB3aEx7vLXyBpQbtoTQwc4bhYPviEYU5xnQQTHTkbIw48nkhXmg1I/nvS8ABog
BY9ZiBA1NRSheWn/LhZr/aXcX1fmeLxIAw5MhDMOW5+IJJhuKYbVoQlddJ2x/pxbXwM79hGvi2oH
ZsfgFu0vn5jMU33C6aH0dEuJsBK97EXZF+9GBsVlckbS216sZJjMIT5D4SMdknpKiG+rwX3ca6We
zXUccNmUFcIyA516otCJKLxxzoXyIxU4MreYLNRxeP2XkHCKJeL64GEN4Ay4aqQctvC9SmfKafU1
N1aplWv9mYuP23S6Z+F5Ygp/XR857e0fe2+YKqv2/8Es1b4W3vyGzCVyf2ShBGE/5FXcUPQJrVTQ
SGzdQmlj9yk+M2sxs6z3mTcpa7MffGdZA2FQDQYc4qQL3Y/zq9A2E17vxgu7UvdWjbORHFNiSpLo
muU+fuzndWUe6iTkytW+w5OjJyixXwM/8jLhNPcQD7ufFIqQ6V2dQfr2YRsweewxsaQxICIsZk0N
ETA2PChIWUXPIUznfUY6489PM2ydq9el3pO8Gzb7WgjxsZUgxGMANqizbV4rDfKZPn34QggnOKg/
2KhmFKM3KoBVO2HWw8cebrjttZovB+ofm7+nbUJrkR5+Di5UxYYVQDDBo0hu7BBeE7G/ijy74H0I
HtO9WKA9+69JO4NqhkJiTuPubYaBLEyXJquBKvl8K/5/Q/bCElCfI3TZmE5NSlFkvzqiE1+sCLFj
kfbXqvZfHurzSr9ZTttVyUldcCtleZ3tSnNaZa8FKJ+jHc+4AslerxIi92bZYxcgNvjQwnYut1nK
bczjULgVTyVRJJjbKKbujQtKy1zGiDfmZjnoVRq4Yedg5fU2/WQfiOFBqJpm7S1Kxoov14zEsuF3
vBYjdS+1Zc2HQ1xslSZ6DVkevyWKgtyrzQV0DZuBUeKM3LAMhzZp6tTRhsDYtceZdQTFxNH9Xq9w
IUZnoW89hVIC1YtY5O+8Xmjvt5s8iT4wxta8p1iXf+xTVoEDUie3mrdmsUjxvLGNiCTg7RIcye7d
8h47+eczfheNSHhrgNf+l1UdIRhXj+beoraCaDqr80dERFD1meGYQIM7wYch+IWLTm4+SaG72H3I
JrJRCjd+3/rmJo/11K5Q78zdrux+rUBxG+HKNXiHzAZNTsG4JkYvUYdCIb+M9Aq72nTm4EVJCRbD
UN50sMB/i62lCGwoXoB8dWd2bxbRBKZ88SgQEE6SyRe0rzxCBF4ZA+dlGXvk0qcAkLYx/CUWmFhZ
Q+S9AVMm0g4E6znNNMKASajTsrJw6ODAYf9SEfmbHgu9KKYRwsBWIFfOBqkWIana+XTolwAZ7xOO
0nknRY6paTJeyWMezam+W4ohjJj6H6h+lHbFjqx2qTANPzAvZJal5DINiRUh7Yhm6/lJKEof86Bt
LG/yjOulL2coAJBMddveAYL+Hrqs1b6tHxyadzy7yvqUHXgd1T87fmJOmvGkgbPIzuSgrpj84o/x
nCCrMXxA3wseoFKcKvgRW96L1qN2Bot1q2Bf6VrWb4mbwBanHU+NckleOWjkIAXPruExW5J4HjM3
9YY2aG68aaZ+dpPpzcEJBsBCzAmJI6cBQZC0vlSAtmmqoaf2UtWMTd1NLswwgjB4aCFykFDLC4Tu
AmERSLSe/AonUGoyybaZZElJKKn+tOQFR4LhtZP7SkzrDdpJzTOmqTKQGGW1jKGegGkXSWWhHWS+
8W2THmH7DWmclnX2aDNaUpVU3ym/XZClO7FiDPw4QOQQAH4h6djfpiOGiGPD5Ue+uQJDTFbNe2cq
fInzkr6xrBOUNCYinUcq1eJ/ql9UmIG+ZYSRO2quy3PMgE7Ab6B4r//V4iqMmQgaExYFVqQeUfvz
9c19gdrSktFYjXj1t2iPAVwE3w0SPkV3nUEDPui7eveoE5RMBnVAMrP51d8p9G3sXXE72d0tIuFi
E+2axAL7wKO3urogFDNEBsg1Wk+vHC59UbDDpzKJlqaDSIlRmgaSD7+JAtxtqlBDmfgJbRucAexZ
gjMPkKOt5zKFevwFUDU99hWSxn+Dz5bUbckrMvoCyfdD/BO+oVT8kxgFtYHHdTF0TeT8rtBc0/NG
n2YHrxcpqjfaaWq4xTSbxbv0crz3Ye818PALviIe5iQ3hrj8mDrzz8eafcSccd80r+uEwKYULt9I
QTmSTbpc5ztunp8PmaJlrTPQiO+46uYdSZKSdhTQ/uCff296NH/doRFo/y5UiTqBNvaZUb6yiRnS
MMwU0daUlrrYnOXp2acfEeQXZ9GYmILf1hhbFxDwMtLzW9KDDopy/VUgFeIkBsmG9lLnfTCgrpEG
NX0Z7fs6HB7dPITLRNwXAdZC80vTW3tAUFIwTXYdTnCh8WKG/oRISIfxegLj6HnWgYl7Bm5GiIGo
Mut9AghuJtnjc6Inxh+G8iDyUkoW9qDDqOUp0+qmOJhrx0tdtVymMWOLLrCJsdwX+vpRP7FQvHaS
SfZm+UVW2R1EjNlul4D2iHnHQmwp1WZINyF87700EcSE/3RwNTBUQPYUEEkbJDeyImN8opFLPgri
hVuQ47AiQ6JGts6TJk6u/6y95Iy/y7nMhzXH4aEbel/ZGMHvaJSZH1hsX7qh/ALY8Rr8c6csKlEy
3oYb5+bsSR5/AVCPl2N5paDgrWpRxKq0s5Wt+hDoRSLyWjbLFYjEF9kbePulNmkbxcT7T0GMPou0
LSfUJaKyYeN7sFIdOMYIvN5n4p0clrh8H20duU9LN7V/wDnQIqvKE9PUtFvyu0gJli/RgHyIxyup
avJgHhlI9hMKtcDHFEZCfJtUT8ipw7kre5gB2zD1KSKC6JYHieYiyit7WzuK5aoEUtjpsArnomAK
AT3d/dpyMGz2j/dYpgdtTpsPwiwLS7fk2AKo+K8AS5+7Xrmcs5XCVyenMRBQBs4bujZdQdy0ar8H
+nPf/q5rrK9xXH4lz6WpskPASyZmm98mpWnNOHuRI0DExULCVDI/giZtSH68PtDL/PNHNZ6tS2wY
fHFSkEgo5tCncdEumOjvXGWMqAVL/Qtkf+4Q/R2U0SSvFbM9/tSA3pZ79QonE/gh9S1MMK6I8psZ
zGiGCXkRZRqt86CCR04jsCSU/xA0IOqUkj7Bfmiqsv/AnsLA6FEVO6/8OzwY+0N/y38+9OU9+LmQ
bPcHh5qRcdZ89EqfZGByxxa4sDa9j2SeOtZO88g0tyLUp1sG+UBR371qd74d7N8FUW2zI0LdzgX7
Ljih2X8HGVdfiwphb+3a/vBWmd5Kj0A0phHbcdee3f5BDEQmHc+Arvfwijx8TKeJdp0A/pRo+lC0
7Oy1Upn3q1VorXvvU//8Hk1uzfuq+yNrrsUytX0S2kjRy72hOMCZtMUVtOzn3ZLs0rmxsFr5Grh8
ICOK/anxfYeDKZxpQ3PJsanOreMlmRdrbpKEGEhbKFUAwtLaLDQGzosFREtfLAoSp4Qi6K+8e7h9
IcB9Iiaqgriyy/hBT1AMVE1BCm+zdYZmlFOsAURp09PSors016bGGKY0Ulch/CyusB8KzqjfxS0U
C0b9G/1kFQIli/flJUkqVLbkrIVuwJy5gR56NyfJ8ccNzFHvkBvInRsHCNMz/c2mCB1s5VBAH3h2
K969FPHX37bbr66NGXYjrqOiFfVXNg2u+QFBpkHVAmg/+U40JoagopfkqVOoKcdBRFwOfdWrhcDS
F+GGvtJF6ODbRl95AVh/MgV1UKFbuC4WEQAEjj6g309WYmPaEKP/7bAN9TGFRp1GJJGX0bGCi6kZ
34tTemgNmOXdu6no7DAmZs26HzqFvBqPlgujbkWNpFgeQA7iIABXDRDvut8xIpncPrJeHgzJ4f5V
5rw5ZKDs4Z8qBULIwzeuQPDdy3QECCe+crGs8LtQnKC9wbnZS5Om3LtYEaBlruIlci6xQpCEDTad
m/npXXS2N39zAhk4DNaPoA3jfPnWjgDoSgALdfiApvLCEW72R9dTmg3GUhPR+C3ighdkNQU7Ia2d
LNx7ww/OJU4iQZX/8Db6xniCWiMaN8vuYy9bR8ts7JOp/r+QBLF+RkUXXlQBVCKEtwGxYR77qzh6
scrqlahCaypbVL/x9sKMjkPOeLvrLuf1YJeU3yztelRoMW1HDPggM/g9e/6eMRHya5gjEDTA7Xso
kdth/ocXMdIEyrilk9/yAx5Y1wtZpL5KnccExG8K4Bco+wqqd8nWJ51ZR3QTD4yfXgZiWMym3Qdc
m8sZdnZQGsB9eG3GAS6/XsvoBfQ5FDZX0kcLGRCykCud/BvX4xUE18il0/QWzz7hynQiEcv+w9hJ
s9FpkoiVqWAPKUlEyX9kg9EgmReFRNuc64bxdszezJ7jFN0gz64Vtly4IOdmN3FErDDBuOGa/1fS
0RqqQLBCiBOHZUizBh+07226qOgsvO0+xXHiiy7mkUZgaualygYq40h91oh9JufP/Vx6y0wbYrCW
Xin6w4qybE3IFayeFl416UMlgCmQhH2vspfBUL/1vxC7ea0Kbj0Nw2Ol2AlgTuctu+Crk/NE/mLJ
KglIUbTKaJqFmxmlI2XCxa2cmbpHkvuOdvvaZB4gsLfEJFNJma4Kj0+VaN7G3yDPEy35D+INfeaZ
yN9tRVsWqP4I2MO9I6Kr4954q8ZYTGfVenkl7torJ3P67CwzAOA4sYayNrbs8WMR7zbYdIUkHLCF
kMTdv2bJrFaD8OQZwHTvFPkbWI0+yhAP+rJd4+mjPfyaRMmTbq/tKz4P9PQWC8FEnupvIUBonhks
4HtL3xD+9bbcgwyyn+U5t4W6p2aErzhcofdB0/qMiN6niQMt1cDM0tBCGKYPrRnTIseY6nqf24RA
K+GozdtFKiMa/ADUgQYP2DT1AT5W0P/G7bUsJzA11buPZohzVDalAWU0F6JarreNPxyYq1y4IWZ3
M//WcL2OVC1263Ifuiv6ADHUHK832mCMSGpRlB+7kzbZKpMoa3D4T87kar3nrXf2RWluRqLr9PXt
TMNI0+K9sX5qEE6O3vRguGVeOadrk2zewZeQRlEXsA1lCvTv/pa1l2ln2vz70jNg0Ps+y5jRvcUI
EhREdud/1Pm1ijszV9vU14QUKKglbqySX3bQjeXgbkG0q1YYmXQrLSmgq3THa2fSy5joK7IBH38q
hehmJsXqhKnjcR4U/b6YzpHcrkXpUE/p6wvSRqREVCkmmu+q50BYD5EvjuuE37GPFYIY+ZsT0LWx
FmvCfH3MxAk7mpPz3/3IUZZVHc9zxB1nfraufbma5grtUhN+q4j7KYr4e4ehvd1kAjJl6kFjeUIq
eIXqHsGjDo37c229AkyKQRY5IF51labNh/Rck8YyjlQ2rnTsze9WvLxNfmLVV+qU/oe5N/ozo5Rg
Fco0SINYFbQeXwX5XC02wH5hgFLovYSvR/mX2NmumxPm3IxoEYWRVu+GE1ElLr8J/eA8aEXieIrb
hAtf4pl7EpIEu3ZDzumOfdujsG1uuOfkuF4BVwLZHE4c4+bBY61KninX7XGOV0d06VGZ/wU/qdqX
gQekFozCeqC428NDSu66aaXFdGfPIgsdZBUv+PD9k73jrSmjs+liPLQHqzDHOGKA9S/h63ptKv+V
Zr/JZxo/X9HtSWyitm2BkjbSXcWS/TAsqwAmZdPyLTiTaiwI6wJWNytgBP1plqWIr9MH1kmqTo9a
tc1iPCiQ/GWFmNjK+HUw1ey2cP5joUhzPI90EIrB91zZFlyGBIm1Qp6vKQHQ6wNFYvOMRzUx8ALz
R/RRhUC6AGyXGlAIxjH9eyLlH8HvrTeDVlU2W+I6QUuOmPbnv2Ef1Z6/8mSIbl5Uxs3CQW99/NkN
dSI8SRx/t62SIpwpqe8KDxgtFUVLM2yPXZwADtZFdJ+gmTLERLzYmmfuojWH6q8HDiXCHoYQSJXI
MqFV1o0vTJTFb1/rAwMEL4fHRHPTp3L68FJJxG61TaJVD5uk3TiXC3vLldf6lyONuoC2fFWHZ1eG
2zt+01pnd2NASehblUAiW+pmZa1qEtX+i/mFbzacccFgqHl3xPCQ7RyFYaIV6ls1T5B+HzT4BKcy
KSoVDIONGNykTQCayeFEEX/UVG372p1CX+hxxL7rr5KnNr/S//+KtoT8SsAEwqaFq46z5g2eStiC
E7C+lQCMikOooAJe33hPrgl3Q3sj2YGnMerEbKx8J2dEnCzEdxperpXyNJfe1WvyCu468kYgO3IM
Ydrahc/02IioGtg+K5d6vjcDFVb/fXMIQF0JGvEVVOOht/XpieKvV45dwLohK/JYywMdbMccOZXi
EZ08HrlH9IqYBpkCKjUpCM9h+kuOiRS8PHN+abW2lvLlosrklX7+jQQBKdRrnUrG5fTv5jB5E2xu
QrLcH4H3aGw86ahDBBSnUBOtzUMQPwKiTyeywo9LqBBGKRcTSqCqvu1wt6zBPKPsISLtMgH6OI0C
7qLpe3SdxEnjq95YT+FzVxqyGWIaKOcpb7Zo4XtCnyecccRMan5m9jtMM9c6xmqJikarz5g+Quvr
TWY6sXxiwCVfG8TitmS289aAMvfUaOmQh4sh/7AwaLvdv0Anp4q6c4Fg9vUCtoczC+xQLqyPUoCn
JlZMt9vtdK6RGpL7odbq+j9bk2RGwBkF0X7GNYGweGJf7nAKoWqzrcX5WxXmags8LykwsNfqW50J
/7WUzdOu6RV7oNp2g/To/o+Rwv24eR5r8/3gSyeM6sNRSEspAAp+EJaS1fdPkN7m+UNbwvHvmYjy
AZ2jXQF/BktBmjhNmf539QO/yAI4hpaO94HLWIyWugHf3z5acT9dztqlc33vO/eu4yeHMZi0OCcu
IkJk1smSaYA11bhG7XMlnR7uISo/Fliiqk/iOBs3RPFHUzlDNE7asbevQ5/Zcd8kTNVKV5npCPzG
S1kwV1ubwQY7h+GzTbexYCDPiz9k6DQASD081hadh1tCgunpYzmErJhyA70kdjYF8B4McPYTiGfJ
oh0x1R1ws1kF4yo41UsJdCzruf2sjjHGlrzwag0G0rn5Z1/g7IDuBkPj1IIzOWIsu3Rua7UI1pzI
t3MToFtdybtmhbbqH53FvK6vm2kYF9EQK9jLF8OqUw9SeEAaLwpAxyopD+AWLkv0LKCAgTMSY0Qj
UIe/rZGVUGPsZSarNeQPGzDSjGjUB0rwaj6jM/xMnyKD1ZU5lFJzqoaiFQLppGPV5JkclF0t5/vt
WXXPUz7XXIEx6cKAh3WeKkl8kmw9dHEjKMr8xJ/ViSti8kRpGsZ70R/fq6ntmhNaXaXLDC6CmTXL
mTyHg/fClFq0wl4SQZ+NmbZdnACtixlYIFLQ/gA1cWXsP1JxrehxEPP5K3SaVSV83XAqviwVLBeF
VRvtlPLXaBiHhkudYa302EK7zzfdAC0fI2LnI4UF1e/NMSu8Rxd8TzgeIHWoDknz18bArmoQ+uIP
VQPJ8/dkTpYlluT48VjwGTi/rsWwvrhLRsEbVCDN6TgtZUuXfl+KsD9A/zLAP5SrFYCh+JwnEm4h
XdeuSv7Qb2KMl4iXZqnLYlED2diZQGC1Axcg8WEuCK4oxeLpSUrSe1mJBkW7DU1/j2a5lU+VDy/R
l/63na/R7/o3DVffF2Ti6uHhvaH+vcoPQcGBlmtxiDiteMPoQOamFh4iipupSoi0Non+TeOaep7V
TLCc+/azTy/swaPXbmyWORNdicz4GnJ4iuSZ7qg3STp0d2gB52upDpX2Mi0rcTkWZOenymKEzmxV
Uamt5vgge0tbfehORPLA485uWrqvaswsx5Y+C1pfjiCI9jtxr6HMg2x17+jG6wmg2aXGpEuE7lVD
eh/O12fSkL0GT4HXHsEHi783mpdamGEDZ3rbUW/ZwbQBPEGhgjjQNpPyIl7ZDk9RdqBQkKzhn4JD
HMtKNP4zRffAxbveq8+dFXBOfePjLEMmjADY8q7jakSOMaZu51etRp8k17f2cfBuFEq8twfEliKu
P/HaJeDmgbk3YGxnYemkGiIWykw0o6J3dH8QQzM/DaBQOmnZb02/mcEHVSXws5S7QZ1twu1uqFYc
P/XPHabfmz90ZWcpvEFFJq2rWMCPDCNfYGmRKpxXujwM91oMEmqRJc/X8mfK+TGc8sFKNbM3PqKD
vUxr1sxeinP1Nu4cn39NRzBDEM4bMy7oupQ+p84gAfX5/o4L0xVzTF4eGZpnqnk5ZopUhOa6KIq/
Gghh00xBSbvZUieT2kt+NWRNZukpqNsLWMKgTLJnqxG5BKyn0Wa9oXy7kUD5SYb5yZdUKSDyBi8k
DG1rL6i6xd7NKZAca3nJcEXacHKDx0zVBMZe/v6zru8QKNTQGjJW02dtWePkU3GT9tdM1TuLr8Ho
9hF+aKgh0jPKJpfhfzt6xqqsfp1G/tNVVtP1gmGmGaEkjudwNmuN3ILfaAArhaOYaQqtbAP2G2ze
mah7xxDJv2BEfPupoxluBDSG6dTUatrNhG5IdYisxt8fR2WH/YV2y0QtE7VaFY1nzJqtb+ZpeJN6
RfLyIKuF+m4CQ93H21hBwSx4ZAgsJhQDlbGV6jFPvNYd+N5KuhddNYBVKZDe61iUC8GC48eWT71s
7wBx3PKIVlrYwEL+kwtWpOYr39Siqu/jcqB5Jhg2w75KKAXmmwTAXjAdRnCf1AQCIvgTHRuwsM0F
m0elQhkvJPoNkL1bEBC+DRno/K9y/zrSZ1jawISfSAD32OfdmtJvgBSt45YfQnBX02KmQTPbZUXo
ffX1RKlWTujziCwHIh1b6DStHkM4COoiG3ccdf4wdL1eBpDC8GfzXcs8lwO4ubiKfSC2s/Xd9vo3
mf7JIZoonowEPTYEjvjMWCxcJIcE/qZlaxFAVpz0yDycbsrqKezGGZvqct8THxcrwQMYyI5fQGmk
Z4Iabhqk7Y2aMANM2FuFq71WlGhLIQJFVuXctagdYQ4A/pg6deRgQGdXDkxcdjqV5A9J2JHWrj02
ID9Ap5bSfX/TgNTITuoljUmz1RWmu+tRGRNxFjh09cLYWJ+jizNDolp8oVc9bhnx+fGExqrlFrnU
nB87jCXBOZCgu7aMg7Tu6e1TkXOZK2beUEU8DbVQ9DbEvFFXqEJp6l24/vlmA25LNK2Xu07KivAq
P3J6DH1oSoI4/dtQ7QHaAaqvSyaY2tJfEjmOlejz6oq95rIpxA8GPx1kMtz1bgUhnxQjpnOfRzWT
sYdu5qqaN4N9STDqbqrPpZgfGjSCjy+IzjTy0KXv2/Pr1isAWw8CGBFs7fmq9tWGN19HhuIyOLEr
Q10V7QfdQrs37Q24/Rts2huGC5ux1HdN5rLn8amNCXBjjJ0tGTYkEPI2jimj21r5gmfm5/mREQmb
TGpv2FRKZyq/m756WGDY50gDqJhT3fJMLt0D8hYVyta8DmppHdwtsB6jl/dFsapN6iWnp4NtGWPp
6j6GxFTGLSYtyf8DxAe5uzKtN/xeNBQZ1w0fxam0gJMk2SCSRMWBMcXIMkIe0KtQzYp0g6E/LByU
iVbbGAPyZYKiqmIhkcHFxpLuY+ec9vcy/9qNcUZriPkkywgeMCSmxMbo+mkAPn+buuG/7ooSSDR6
ne0RxBMD6BsbRWeEsucCz29N6FFBc1sTnpeAx1nGEXkKUouTcTA+VfC8thA1kYk6WdpV08cPt4mI
QKT28UHUiAyJbJUOW0NmEE0FEUebG2cLwEYxxScZHxWOjzDB4HyCMEbfsHpwJ4E7APsghuaz1h5k
8f9xo5pASDLBMjoxAYdmelCtASCDfn0zzCkQEsHkUfbZooQTrYb0Z6zvQYlv7sRgCfYEnAa5H2db
ELjb6tVBx5rT415mhYUUuruaI6PbxjHlUWlkEt5jIQh9PgjqXaaznlAwa8Ga7LEtDYK6L82QPovj
r1EWm0U40ciy9FufoU06a7ymTAnwyl9ml9dn/HzH2kl5CV0/e4ihEzE5cUpoV0kbSXsFTPSARLJA
Ydgd20BgUPR/fq47WVq5WIPaLB6Lsip6d0po0lIbVPzcdk3VG4BxMT3NxNzJxb27hFue3pd9g8Rz
Bl7Lt3YwJoGZVMzd4JLy9STpFQeMrFTWaWMysN3Omr14/X6SPl9fHrqlDFVNvV7CEWl3XMSnf89g
sja0/ruHDUO9NCqJrePeF0auN6V+kAA8powRe+zi47eVAygtCXKOqt8BpEpw59sMlBrcKYIWFwQr
Sr6EYWTlYN8UmvmZd8r+YjWzqZtskNWtXxYiXZTtJUzLryXOpIJJV74k5kBqozTdtNUqSZRgL2Zg
Cwdfj+Bd9wbD0K5RrTVM8N6FdyYw7hwqgcEVKawW2a2wYZouFd76B+v+q+xfo7hlYf0/zxhyGIHM
YjCFLR/IkjJGEuI+U7nDumAesTPfmjlclupIpEWmx2R9hXBL4WNAyduii7dxJI27tkEdoFGLpsoA
aysFnLh100nlnNlstmRcCtY8sSW4gJx5rd/MBpLN8KJvjqQl8aErcvPphL7ezcM4SbMmSwtE21nK
OvKFuy9cyBqgiOS/rHDMywcKsA7BUeSaB2TDPvl0EqfEGcz7JNStTL6hZNMXHdg0FATk+j+y0XgD
2MP/LObxlyjYTb17xmNIrKuJYQSXyQCId+bOPSL0IZBlaf/3yM3RftWUj98LhuJ3w8TbUfwF18gP
3FI9PeZlPUKxEW7FvpMsOst5rVauTgmDwf/FcMeeYlacmWI7O56nWdWIaRp/lEVTOLF7ypcHRd85
mbjQHMV8/LWDw88deRCXWcJ1Bzw4gTbx3OTDjhZVFH+oySVivpATznvcLpHJDnFXc9B/S3+nJ/YM
anOUWznVgS9NKKOOLchknOEB/NDHLWnxIJ/ayxYGBfG5a/Or1SCvhElEvpeRoI3HB04tSvAzqmIu
kPypNpnD2kJtisA9BxqHLv6PInkXipCQC091yiCDhTpFuCMRe4smZiMwozi2H4BStXPzAiBs2vX5
GwNoR6Pi2ILArCTL6C9fs08+ma2Beyo7LXB9CyTTkisbLTGsCPbGxm06kTMvKseLrwN1/3kL+My9
fJiw6GnHWgn8ndF9CyjqtqcQm06TzRfZ6mcUhPR001hmnsVrCv7R3OuBpwLB7NLkVVdIcZeNuSls
k9WmZUOFv+onTSc85PlY7UNn2A0ZCibiVbAr53cU7B3YeOXHjf+W+zkZWJ1PSbcMSZLLnKcnIs5d
kkVXE5ayWVOevtsq98/OHstQ5oKuyHQjtpUiKJyh5AaPfNTgHNIMC3DwFUhVg3OUvqMZ2eW2XuJr
CvjaKrqGoovIou2o/0etZgyiNRqCOS7acudQ12CsGcDhevnzV0YDiJEwnPzYiyYfC42OJP+VHd02
1v8l5obd/ocJZHCr72HLpGbS3F1Kq4F17Og+L+WBdKQcpub34+uH7eXZUH6j+sD4Bxd6BBnR2DAE
QeGdHwZ9QGpxEpXbqzn/T8R3yS5dchpVMx2N+pY9dYj6Xl/nEvfK4Kp9xorEJa6fSXzhHu5X/UFB
I8eG65dNTboaRTbAm18G5M2pkQfiQka/Zkldam+CjlsNG+HtipESqnjXIU0LtpjDnj2rf9HaevWr
t/pCllLtgLIZ5h/s4xyJaegNl7HsmOD4um2QmWOwGOAj+pESOGiHR6JR+Q4NEnrbc/O1RcvJUbWA
m/qc8kNTmufG6G7mfNELClOwRWMke8Ce51t6HXg1YUXkMungSEo3Ap5s0PiREFlpxOq1szVDE7Kq
ofK5dxB5vRazn4r2EoePfiQTaWUqS8SLlDxadL4xQT1bsLO4CHNkg2aFLOHPBNnWYbEsHvqa5mii
EGgOlNOw03ICrJLJI5zBYB2RH04EInehsjMpx/FlBFB3HhfMw9/3vAfEQ32Oxi9KERupO6+e5Ycm
WkatKQ1JoetNGmg7aSBffru+KjkJACVggBJpfXP2XgAQt2NLdtYiQj6curdaJuBl5hHMC0h8dhAB
OTfsyUMK8mszAoNYCvoT87g5eTYdoI2+Qo9toMO0gvGNHy2c7Gn2X8YV3hPp0sBxVGsLflBsnQC3
2kJWbeHdr7XFe/jAGUe8xKSORblX8w3vIIGTrkxzGmVTNtMqV3UDeINy/37GZ/a+C2tFrLIxDnyA
P23Ck6yVb5Xxmb1w+Hr1XY5/owRpoAqmScuD9/54twXKd0FsS56mxcIw8GxMjE3BpN5QS66jptFc
DzoyHe/XLTC5Iu2KjqFw6HvmP5Mt3kFlxH4X7spnyvQmQk8oCsLvRu8Jb9TLzNnpJZsJFGB2Ujhg
39LL02hgdPQ+QRe6nhN3HZqTMOwxNKjwHqsdWaJLN8y0PKCF35Na5Cfcb5V+6qZX4OqgaAVziFBF
4TqJOzb5o0eg4gGQXsfjGidp9YHsGStTSu6m12HcevDirVNMpaltSAjpJ6VRDH2sAAXLpfMB88Or
zKyJpUhQk1ynjuyWEjv5jmN/u3aLluCr00HShQ/KeDWeakF3WMJvt7Tr9rUoJK3ud/5WqZ4d5V8T
cd4dKfKJ2hl0bIIdHyXTb8xtJyewRDcdwKQ95aktCrLb1lrAvT9363sYM3wAVKxQLCSsUXGMbgnw
Yqdmi2oueNnH/tVnq2Mm6Y6iKfXtyHjtx9DULwdirNvzqEzoQ/1FKW0xytSj+V/s+QcFjYvPXfab
8DU4P/+aKYUx7WeZNP4gsn/8DCCyLlgoDlP9/RJahDBvCs61EmBtkgNj30Y2q0B3KLvoUGjb36Fr
TC0auIaF8z44JMEP6gDm4/nBbJEU9oPZOf1nGy0okOIPAVe8YCt31eGZVBUlDHv+dSW+ULo4M71h
9l1oxq2tYqO66dFzgJfPhjIhbgYUPT6NahAQyDZIiYUFPCvMpegr72l5diCyQwOPMx6aIFL2GsOi
FBpNI6TCDWuG+6CH3BkP3wicAS60WgHkVhqqJDYhIbga0/n2I0RV6sUrMy87+zFGrKInlj1DQimK
l0EG+pehIrDZcmg2wx3C1mKOXNPX05lXdJpYpRJGD3CeMjqaz6O5Htcz2oeWVnUl9zGGjMNETRi8
Rcs07fJcyciF0aHwfzFVUGN7shQZWkLw9ZGMKvHe+Fod4M1yjBmjULMC9s0hRq7d9A4/9U3uJR7K
5c4O0Pm/AXE6pCmDWth0E09PtqizCwVee+bZoZc32arJq1+lJSimA/ERvs5BycE1ztqMsW345alO
hniCK0Qz8ka2yYSzCbw8RlVmZBY1jxO3IbmoHAY2msN+/SS3dGh1F4PHeEiwSxO4bFNPBJ/sYdBb
Aj2wDU2aLalru97L++npFsnoYUHnucfZj+CXuMQ2WsNnjmRMRRPATHahT4Ht6sKbCEQlPvXinDor
NCrOqxvAzfJXngZSinIXE+IFBfRELxnHXw1sZOho2fQK7tlg7r/zcF6vOjqdinAaa4KDBaP4jpXF
Mc4u8eZKcZmFX2D8HQ0M/CooHaDURvo+EcD1zPlja0KWxY4UalsAH+ZCYmuqAHDoA6P+M5WQlfZD
UL6GkiuVD7/ijfXNl1hy7w1dvk/FJIB4iZM0ddRA0S++/TqszSF0pW4lbIQ3/277E3+Or7fMX8yp
vg1bBXAem4kz03DYSlC9xufIbIJ1QuWipAx0CsiUVTHedMjZlo84dCd/vIzf40NyFg1nHVYkhd50
AvVRVHZOLqdTghl0MPhaNzD4bIWwipRgaJWU8H0TayzDDyPEWBsS+IQhAMB69K9WY9SK9C1JGbRT
uohNNa2Titnr3wGh5gx836lN9amZmrZhY+pI+xg1raGr1070MH62bcXZDiW6p9WNB9YBDb+ONo1g
5YgAHNouzGevA5IB66igysEyWq4KAKeo9/tgA0iVzxmog2ucgl12vdwYKHY5J5Rfcd51xkGyc48D
IIPiTZ2LIJzbTC2FcedRZ13BA+rf935oGDGNnw98dtcY2YRnHOhjbLfLYTnxVnTSHV0Mp30DNJaW
+tuyi0+H+XlzBLvDxt535B7FqmgWJ+/TbbjNr7L60eN1CQwuQGRApHtiADoXZ5erLL53VP4y1eJh
+dTgDtNxrto31Vb1uP1LRtFgq5I2OFc0DaH+qaTgWERCRH8mEbp5mzPmo8y6r6WD7LXGef3eAacG
vu1vCNWO3S0Q5HZiN+qpylYV8dksXi9VWEQ1BWV5dRK435Bclu5HsMK91B4vxreTwKCiVcoZRmQu
ixLU0k3b4do6c/9ZlWPFtUtcNRv3oQtOWqXEG+FaGwQbOdFGsxYXHI40GlYsMlNdfHuVbZ6WKHgo
cgz0iYnEZIagkY9QRMexryjo+d4VkaYuZuYh20nYw4qO79sqr9avBJCM/8dZMdVXKJsunqI/3G4z
U/wV00yE/PzIvR0yTnCYKKX9bjfXGDm4oedGXg3A0CFHiuM1wrZPwQUfIL8wiYuk0Xvq788GsWQz
eC7xVJDaShgUbY7GaSFl7nfxiWyOmgYfEUGs4KqhvsC9KMVoTwyIGho4u8ZCi8u/BApZtmMUppeb
n29+Y9gX3+2maBIwmRrfioZmFz5BC507vlBtvPG+ESrcF0exg77k/ggvHvNB7iVxqm4y0Gpinqsc
zM82ZKPSmHq99oBDJuP08xwPDUY8Oh6E7Oe/FfUiDzy8+Pth4k7jXfgPqh8IWF0MHuPE3+qIuj93
idm9aAhkM1GYSMbHtFt9cZ1HrVNVVJWtzmWCv74gsh1fT2xLfwBYAxfuF/T9j3AxSqZ+rhAFXzT4
i0HfZPfJkv/Gdk6lkL/ttpkiT+nGNjHTtCJ7F0n1p06sgnWez1Axkz4SlX1St5U2VKpIpww+ezD/
lHHraiAHvSkUsFlngmnKqGmwkOdoTYSWKSs3CAl8pBRQSAq2q3ClGdwb/PXnqQcnw6h5PCkjhLVY
tpQVpwSm8bDC1ziuYRwS6QO8uOuCovvDlTYzJSEuEpFm973twByJzIAR64tmTXHpWX0JQuLp9Cfi
xa4BUkyrjNFXx/rPAKL1lcCuDTLLuqT2zDedU97jjshmK6H2pCnYGjs+D8qVuJSTYk1OI4mEoLv8
uvzurixX4Vw8HrB3E3A7bru6zpkc7n2kmtXNGnFBYPOv7p01nVVTpfB3rNIeh4lF4/5L6NSuVY0l
UM8dwfKbyjBO0dsZZxc12i+TDhlTr49Fqe/HeLucgdhKJF6X53dQZIo+KT6+FGqnWHJragXMTEjb
heGz1cjCcvZAI2UufCwt89beddxIEEikBXceRby/CY1nK/8e8lkQ0KIXzPJqeMeXO5XM1gmCdDDT
4Ipa/e68ORJxk6rej505nZjYNJNQAZUOcCkyH2HFife5JPW6MGVzLVxFizFxNlmn+Zk9zA8YBbWi
07c+bij670/vrjw7ZwJkYWiaPiRSD7aJRwV9ra/WsgX//N3XTaB7dxMK86mK/xhcXcYBuLFsPPL3
EuA/o6EkRc0uXZIsfLhfidjjq1p90S9SLSZg1Gl9FPF7LSGX/0ziYL3nobn/2QGONIIM4eQ1sXWI
UCRNWja9U4BqOF1Xh5WoFe8BvT7hDgUrItdGwXY2miXzjHlNFz/o6Zdbw7vA9Bjd4FavP4jwt+90
Qky2dvmyqVMFueOaEnBVdcOQCDU0eqMIzi/a8o0KCck25ehfp1YaEdKQbEGwotXbXj28RpGiE7sE
NjHjG3ZtzkWznDbDxhVN6n12Ey/qZggktDrSk2lycaRgNkRQmqFX70NqGvkREK0+5abnpQpx67cz
etwUlfinvf0MBbM1Dps0kYOkI52epa2BlKRYRSmqvFDtLttgDeoSov6kOdgRh+vbgB6kAJka2Uea
cjL9ZIk3MDz/RkinteXXz7uZnwQsnaEE1pfNX1MDuzhRJ688DR3GPIv939azhfO6PIGk0Mt3e33B
+T7rTAneHughJkNBEGaL0DJyfRxjnWOYEu1mEVC7ddMm6QQvwnMoexClfY7y3/qbBUEET6BGnXUI
VfoDYxYPSPEkriLjh1rjvI3XklIN4DUvkwNkivKKyLoVWZ1eiZizUzWvCyivn3yuaJeHz/tmrWLF
f6PuG4oS/MrLJKW5zmMWjEMqaSvkdVc85aTEK9PQHl3epD/+ThLSh6JhEbtilmd89sY0XrtnJxEA
tQ0rF5tX6y/rfDZcA+GNEaZMVvclcVrzToyqYJUZlFCiO5tv2VtnvIvJQKsI/NI/UTjVIAqS8kr9
ZRUG+w63Z/yvPkBAPZKj9pP+V69WNUQ+CSbMOJ/eNAfJBCrQ7MhD+EPDPHCdN6EtZrGAJAlZi9yf
7O1cTZ9unQeoK9J4GPaJPlvrRsAf8ptaA4628p/7Wiq4uJWL5+FSBRnFJ4R+NEoj22z3zjYz84wd
izOh1hWiIgqiRw38XQqQ/nAUR1wYRQTLsA44/G0rmnq0QA97jlyhyrd1HPeEW3WRGeLPj8QrschL
w5s36aKDH4iWPxDLod00aI9JtGMlF7APXpRAJ0Ctz8ywHPuK6IQURHcS/kvK7ngoSO6Hw650AGlF
sO5Ijymj2RCR4X+Va4eE4CdVWzSJllnGiQcbjLXhR5TbCcQzFUU7VRVuBQCjTD9G3ZLZf+R/Eqj+
aIAjDF/h95t3CV0fSaOwKbsu+G0ox04gasYtV95XnJg++qDYahiZXQD13ewmyNNZ/uA2tssu/QY9
g1w2pqHpsSIEN6nl4Stiwll+0X2K1tt96spVXe3UrsFX9mfhfnfYMJ+zLGVV2b6iijSs0SEEQfS5
L0uis265Exd3zUzavyyvlckaJK1YmF8kYiSHwEiJxdz31hHXZClqlzNFRDZjc26mBz4sezs5ksca
wGDc5hAxMhdmbDOsWO1qQiYs3oo8zjTdEqaAsPXCoRcSWEmlSNcxijX5WPLLZ8lhGQcuiQH6kvaf
XIOJ/AkwRaE2ppIZkejw2Z+NUGhc4urNJqLFuuseYOBzWQe2MLtL97XLbe1mMcHdYdsr8lCFu0jA
303p1t96hHgHrkutb/GhdI6yT9QHlxnSRi2ShVRDkHUO76r1H8F5Bv+5b5CLOPYRGLp0mPT/qEZa
NRYe0yLTtoaqhE4OWhfO0rT66dd1uO4lM/R+dwHjjp2X1MSNrcfPJLLFuPMpQAcBUfvGUQaMT6Gt
XfMemqrJwsiJwP3hHrb6kglALftOopdGjJ4YrIyOBwk+VNFvhzufsILJsQlgqcEshOZNqcqVrUAj
O3x77FQI6TaiX6TSrpWHpUu4Xioe/AuMpp14XZGURD7dZGrtrP5beTZQYU1qyDd1u9QteAzawNen
FpGHcq7r5Bhe8yc9n752aRZgMwR1Sw2F6huXmOyI3ttHphM8agcVB2ieEcB0I9r9rn6/SuisqWWf
bN6Vl8zHYXJz1oTN08avhoS/IMQIsTGxKz7Ga5L3WHM9R/xke7ilPbNdl7NNizm0HUH8geLz31Tx
WBP0MwWRy2yEZWSSO8F2K4nN69R/6QVNf3nXEGswbmYq0VtVboOE/VFcJRXVqEfcYG4xnWyMHcND
zIGil98kyG2owMdvlU/qvq08euKsh/qaveVybz0CMzrSfj9ueqAVCj5bm27jhE69ILthZtmJndi+
E6ORmE6jGz9M0OGVMQ5kyzUIRJe9TuGHrWuM1gt5wdGiCv3AoHvi2QhQ+ynTyfGX4jylEsePxuBB
pOFgTeEVCWoFdNCx9R4N3/mqwkB+kxolujOvsCb5fwkDq+IXi+nCqCnQDO+mc6eAy2aETc1XIxgF
DzIwoOZSQIZe4zFtPd0F2+keKImPZxjAY3sZo2V8OmL7YgcNOMEMCylEA5brG0UnHjHbGcrFJDoV
9rDKUPiM65ViTHqLReEtSO9//aDiysiXlF8VgdJEQ/Oq8AsZ0g3Yp1DXNLKf8hdyO21m+Wf1vneE
IP1tJ/Hr/Hjclq2MggDbBoeQBIoK6WuHwPtq4jFTA6r434n+Ga4Vwr05lhBk+uBG1gc9i2W16zNX
XPQ7et8jtVvhvkJdxHgKJUD/u8ICTGvebQ+NjNXi4gq2RH42+OhtfjjkP5L4PalGXQid+xhabviu
XI3lOUuPXxumxWMYp1qNs9CwTD+ztDddblpfahnopYEGDeV3KroKT4pXV0RMDlQQX9AkWuF2RLfy
ZM8XVMWiVreEC2xdQHsoWwt7JUeD1CZ0pZ4sI1ZSytOPCfoRRRTOPUdWIbYljw4I+EY/1KKQDGHP
XKp3c5PuPAR8k5hRyuohA7IGWeGmV7XOJRVYIEV+o8Hyds/IXANNKDY6QzOyfSwYpSnZAtmeHg3Z
LVab8GPcIAOh0XJzM83kYlQXtIzgLA9pVClmu4SA6lghEJeHZ9strKLiozmsbfh2wq+5YYgQj8bN
BPeBRHyKk5vS59UL6654Hw5GSJtowWDblBBvqr2qb1w3tWgk3kf4QTEPoVTYVpDC0fwyB24SCPt8
hDtdd0LsLywMGmn3t5BZHG2avIIqWSmXcdcjWn/yvjN/2p/NsJIFZ7+naSElAO8QwIWFuv+0Fauu
un3xanZBd7gd3x3XSiQqb/p++mMM/F7AfExzYbIIKzVI+6ZVwjg14WiSN1geY6KXUZPwTfjm37G5
jUkR3Mbx/ZfLfzDQwUZ3KsQBVxkD3LE5/Us7rFLGjc4KBkNFKe9waTLZDVFnv+Hqt1W59eLIWNgZ
CYewt2XLKPe0Ad7dE4qrhOPJSi2PvDQmOMHGGE5GxIHpH9I1Ee5zf5yNPq8eKLhfxCDmWmnDSDJM
Xv99YuMadJsqdNMcpboLho/BAhIwhVtefyR70YylcePm5d1dbBkhg9cdz4Tcnf/GX9gYvkKLRMTb
kRR/Ja4psySwTZsWVyIecwF1ovmQ4HKLkGj5+XGeCUOUrIQUfDUBK3HomwipYRsWVi2eN6qVDalS
6XkDplMCCjcZOyqn0MAEE91NsWeF5Y2rMZA6IkEV+PpK7hhuDBmr8NxsILzT2DSfERLDOGhhHvKv
ChoBPh+PiWABibHb/UczqwWoKhCDbKvHqcBolA0l6SuCcybG/OautlWAuybSS47FP2tcOHLsdKYs
jAxHybE9QSqS6ParKGgwnW8jgn6XcMSCHkr/6ImsdJT3B+oxyOJiL723DbhvsCqR8/0yrSjAdrA7
MzaIBZExEDcVGryG1IPtY86D/ZCCrgNUh01W56pQ3ygjenYrXid62ThA0CuUckoM4ZQmJubZj0Cq
vyFS+CyX0Eii09fuN5s8KOx0A4hWo/z9B0A9l9g8vUvOHHtjVMLsGpGxYO7cZ+MQFIUR05Bf6MPw
sxFlo6fCMZuOAEDuwIIVZ5M/+rpnLFOll2XPVZX8bDfGMDBmVzUxJcNvFoOIp7eUDXxml8EsdHvC
yxc1nBWr9ecCJO2mtBMmCS4nY5Wx49cDsqK3LaU0zfqX90XELqbSn3ed5hVgUoBs1Bkv0CW3V8WE
/4O9ECpA5iUsuqku2cQDDD+dienEwe024SY2U4YeexDnZpkXhQlv6PiS/kI55GXdVDSst4jHfQHM
ULqlT1Z7QuInEFsVFGvrgUsJwjhBgSedc7+7RhatWBwsJti8mxWIBnBVSyna7xgD4d5ln72SWusv
DRozqetFuqnZPCqmggyfmJhBkUC9AZxQCvRj398unBNXzfkv4ILf1voq4UoHTLpJwvgsljlNaxXY
YkUDtPmaX6ufcvqp/kQFtRbbJjriFJ5CV1bDy171mJniJ0HXZ41vGzgKXfDL+KTnispCdNfSyOof
AGIKTEcjCKpHh8wN8sCq+OV7ZazwedIjUoEebDbvv3XfxxsuRaP2bKp0p3G7Tp8umOYAo7+rr4Kk
K0RgVYmSgMeL/GgNtlJ04Cib0wvR1QzqNhWI4xyjPQIlwN3+5olOUlQyvkLeQQ3Uq4l1SI+X/N2A
MAkhlTDbJ5qHluOG/2v4jFqu7u6oe2xymvcQ96VQjfJlgZgrt9ZjhvU4ge2lRixTFNsm5h8De8qN
qxEA750GIHa8pjFyA2uXxWx2RM+XMEedKkbzgaFUYNTgPC8ehzpuLne+FuGo69mq0SUe9Ob4SFj5
gfh4AUzyXC/UJ1uYr9Ir/5xgFbKaF6gy08tjPSNQ9YQqq6t0k/XGlbO6eiipPqq+TcDx/ny0FfX3
0CukVAwirdQlwTz7+fuS/4ULL2cx6HNASTK1KxsMDn14p5+naA4L9TMMo/wPDQemXQ8NVBoC/OEG
V14abiY0oeHSVLkZiEMvbFDqKSZK5Z//Omhs4Nou3A2PGW/zBbgflIfQnuwtQwP6nqw2yqJdi4aM
myNJlIl+wBrX0LBkrDlZQRrC9QQcptkLkac+LqhlJimWrdWNSYfYSV5TfV5RHHDj7mpc5+8hLk5m
vWySwBbBo55KnAzQ4FdY3ZUvQObw7+B/BEsCuXqkRQjN/ySayVzI395eShU8kEiqN3szvfIOdYOe
G0ylXhfsOsyD7AwCs8mlUuo6b9Y+qtouAO73wJgMciKazNhBsz7N9wGRX8Q/WIoN+HyO3SCQStuB
3rixMZyiQGA1zQmtQUmjPxu/N91MO5MiHGwVBSmHU2hn55rLulkQ/Ek4UE8xT0mZHOaSPnERbXhZ
avWtGtcbpGfGZRFGX5sNzH3iWXzwvI33uCFo9022c6+4Qrk97FoZ/g8js80pUEDiAvQIgB4Xps5p
vgbjGNFnAky+1Qly6jHxROPFNnTO15WohP2jEGLXCue9+r91CPWwfI+1kYXvgzhQPtGF4V43Xd93
1wxbeIrV4w4IvdwFXnCEwRs+heLuHzPusRQu9Oipe3guWGFGDBNG0A/Z9FhDi2wxbHnaZkVDZbbq
l1kz5lPRb1grf3iSQMF5+IoIt9Y+uTyll3ZVNUPpp1EmQ3U5cX8PzYLfzyYRx5xuFPEWjrINoNys
c1iMmK8E6Ev2M6GJe7XlPQoW9Uc8NnJjEtCF1h/m3IPVsEnQe7l/lxfmayiC2ud5IvDt4vdZ/wE1
IWqUb279muPbF1bgC7pjGU7qeED4IYTz9uW/v4VdDU4pujBvpRl8N5QcktcyPPNiPLKVuhQWY2lg
T/qZRuo4ljS1tVNNpQ35K4T+ry9BBdvpnsX4nAaTDkzFQBznhAW5v/Ed+4jM2B3AjaKrQuh78Wbf
6oF9PnSh0v7C43qCHg6Z9X8aa16eh5GM2LGUmAa8HctfrU8vDUQNGfVdBUqXFTjukDu6z79DqXFM
OwA4845yjpOm9PEY81OSjLuLHWThdtcVtePUaDqxJRPS8tXpCSyhdnSmcmMpOjRwjT33zTy2px4g
oNBvpgN34JFnVhBRo10kyyKIlFLO+EAUf2ZP4MpDqnhR/ugiQCBwpmUuFM4rtWSeHZA8EWwKvWtK
4RxNQg3Z1qow6PhmiH0kZLHrMpmgzXiSj29o5e0PNEOP+qRYNSo2BrmHu6HITy7PSpLJrbagFgln
DFLygYF1o1VpidksBd5zcKDh9Ojkk8TnVicVeuPZIzuWYBOJmvDCTDII/cWQtv+1tlemC55HN7Nc
y4ysQUXPNSpLAoaIfPIfxC2XCSpB2btO1XuH7DhCskedsCGv7nDSJkM4gMJVYExSqmE9hIDKufWf
Wg2XpTyD6X+OY1478Hb2LiLsqMqLU4oex6WgRMrn9SsRe0UmNEye18aekZUseBORDZe0DNnjdavq
b9eeqONpOqaXOUfqEmD+2N+5t7gWpzBO6DVnHdIeA88hnUAMd8O7bQidOI8DyBVddRji5Wu0ddbS
O+4LEFIq3EmRLm4Pz5RuFaHeX683tzvA2+9vpzvJPqIqvq5zNZsynOADKFiOrdhdX4zda3aq8KNn
q3o0/yt6AjVmEkcfSW7pSM0NANFCaEXAPzWD3t+O3W6lcR3EZrRqr4dyWfOhsDaRRil5wJK96X9A
543g9sYvcOzTHPlOWQ7YYRT0c0+EG2eM/08zzyXVmx64jUdw/GPbMGSpCyQ5uuRzuzG6+fCPB2vi
Wy7IQiCYEhSceNpg1lL94+W8rVc/pCLPwpmwqAwC+VDM+zUbZgrOO3UbN4sDRUwjPr5lpqv59PpI
r0RgWxTZs00rIjTi7uM64oZQhIEy0trwhTMj8kccD3AYxoN3B5202XM+gUv3BYlRutzylhCmqD6c
j4VZrYB208RBKYwF6wWulVivoXeZdKxJ6us6YVn/UhWxuk9O0h6xjK9AFx7Xuw+i6pEDpGOb/xUx
ON16uh8a1QT3I0tQZhQ0Bryi6nzl2Fg/JdyMvAOc1c8WgkOaHJIHswqxxbowNPi2FOuW6ct/Ncba
oSTvZnHfGStlXG/ryrjRE5BMPWDl5HlqubcZ7QR0iL8yuhGGcwufvOzRzK0hXU3QaDRIQSC3ljfx
FQZYMOTxHDC1GVDj6jYEUNpHfLEfmtjqBr9aIL08hmwfnqEZBleSckgL8h/cKtDBW9Lcfc48XN2D
TqAMmhKuxv8Pt4OsIKHku3sHbAgZPd2O5vaBsOCdlzd66RUko9LYohs9wMYF6eEr/D7J0NDOFpHF
PIWI3KcAGb/EzKUgn2mlEUe/ifuVUVfSZMr58l+/Vlb2nQ4dccE7LNLcTPy8A9Z/OnOEoVDRKJvr
jaQL71FqXMtBGLr+XDSCbAiTWcOUCkMhpOIeC4R1z8O12GQHFUetcHcNlQsRdTygNg2gc4E3cgEy
VhBmkV40q2XQZB0lmHW4gfs++HdKHMxBwQACdgvC7jzIr2v9QB5RsUgEXLV2qhnPAWQKpXioTB5v
/BZg2ySvPgu+1e4sgsiXW4cAEBoCAVMP0aWYiQSUKlc0KOZQtBc3PBVMegnXeH8/BFChQsoTre6H
vXCSQqVE5GsZg6xjajDvVHQYHWk1F/oIxj0yK6wFWE82NprcRfgpJZntCikyWG8IchWMTeVn2ijq
UjLUyAaHJGWqN9X9xHnq3qBayksy89EG+u42Chnf8V474jjnTd1PllBJwZga8u4Wbe9BVYtz2tD6
z2KTPEwHJCxV9C0SdQz8aQuVVrN6Aovz7a2Qqn0CPlnAlPefCprA2VXfBJS0CeXCWhknF/ItDVuE
BrZS+bypSWa77TJi4CbcJGHQuLELqtV59inYVbf4Dtf1JGPSEzgty+0nI1rEvZArG+h4NhJtMYea
SQeZmVR9KSo2wbuPxSwtvpXCLVvqnUIi4nldk5h4QENR97xr9d01BpeOofZCIvsPAAFASg56cNLu
a8VSMLafi9PcthEAEkXjGv5a8I7RPVaaBekxcaMMkPQJBWaWAWtgvry2PqGL7zVqxQztequV4zgo
2uzPIehJ1VQwYVrg4AlevoKR+qKo0aZ9DJg1slaxCAwtDrUxVlI2yinUYveVRPvCQLzAchVGIH6I
9bDQqmwXScRZJ4RJPnnuVIjtAD2f/ejkQnk5o1uWS+H2zP+Lj9ea9axEpR2YQ3YMlHQgEd0GxZjB
kq1l7SAMTDMhA8BOas2nU8OQm5iXdasEYAniioaxXauG31AN/3YTJHd8j2iqLsk0cljgKcMpaXGv
J9QaAw4ZvgCjg1mCVfChm3BMHfWHs2UqL3yerbs4DrxwNFrP7TaahlB84F54+nMMibCOrWqCSABr
Ip7tCFi3ii87ZXStakSNnDNAJW5Uc6Y4FcRAqaviYQFZPRep3yBAJbb4Bz6H0TVyaEOz/pANex7F
QH1/b8Depu2i45f2lVyDiEaOTXw8juoHWZIL2z1IwDWm7H2JiJ65Po26pDhNwqVe/TRquLd6JyjQ
HIYAwGoY3QkYz12JnwQvVHl7Rqs6TDA1Fsk5NuJT5GZbPTZZxAyKSH8yB5XHyyly1kXI0NQa2sqe
DlHVDPpiaVNR+DgLnC/hQUbqQg9h+eDybpLeUAR7gXFV8jTnZknJYgb13B/v8kF6MGJwRsGiA7PJ
6MqaPVzRzKgZTTkGoRIhDBnMrYvb3hA2diVTCU82+XASEfV5s+NrTUEO2zJOouhc0jmbf05sqX2l
BjJMi/9TDb49g5yO2GRciCAjHwoedh/1G5Q7O/KeQCXSdcTez1DfLH0yaG0pvhArbGtSSQfFqo8e
lIqfnkE1n3TJ7K365ne7bvdAwXiNjQf0CDtOVSeQt3dmjVVmcLvFtFTazrpG3Nv4unRL8vSXqmM2
WEZSRapxzaTCl7jsniCwG+HoJlJ7+XnlSnet+4XBlevNQSmR+B6GkXhzLX9i+wAo3uvkCMcDehnn
iQLU4w5mFTjDdwE9q1qhMEt68GQnS+Ledyphhs1CAca91hrNOxNEuyvTOSS3e6iv+wbVu/FgAfpY
l6R70R1/TYYQe+rLiw2lp63tfA0TXY9EccyydfnEkheYRr8nfURobNVu3Q11MLpw/NSddqDmQGo2
n1CEsW05HTbpdHThHlb+TkifZWEjRiL7ZN9If3PtYzseVSigzfy6FuElJAJhKKlSJ1bSeg0e149E
x1NryS2QJsC12Flko1jCgrkoi6rTCSVNAzMzGMgivJufyxpqkjqTHL9oxyjrMgp/hVKCAffXJMIF
4rCCZBw+Ln6w7ZSFdlJVqtX2sAs/F4ZG+pVYarHkYjL4mJXvnvIP01HvwLg+tlVdP5ICzz9B/4rT
YTh+uYBsBEtJbTW7rz2I60SR3DbNCv4CP3hav8Cb0tC8tH6B7NNNFy2Xuxc4j44hrpadYQ4J1WHf
X4P4STp8R95nS0kudrPvWtNdGkjlUS0K2jsGLvCfPhBuRU65IKsyaFc/cxav2wwEcwrjkhwqhMpJ
+DrXtTJ/mHIeaBJbh1l8uo6GgexUloN0ygEu94Mo4NHd8AtclyzONoNt8JD50pnbTpLLTORqVZU+
S4TUUYZakTPuMnmsVOAHly0zyu73bjG5PmV22Hr8AblKVy2IdzEroblAR9odFVBgifj+Ri05jXeO
dpWBP7u4YUfxOTKeEqN1a/CrPgMB5P+zw4s3LJyWtpXXE+endOvdzY5VUaEIE2eYMhhSQnKISKKh
Gbk2JGRiIsQ3VgtxZ3tCCkyA3sP+p+lyTv3zBB8uZfCxVPmfzg5c6QkoMCf2lmeuJ6GvaP7z2kIF
RSSYCbuQl3xZVUl3HfmHHit8LPNRBCkXdVqadS3znahQQRyX3BG8UHysmH/p6m+RCGdgaMduWtXh
dMndxIXHasB6C/W4SV8CzcF2HhCi372EFRopYS6VXPGtn8j+K3+8Tf4IhN3procNTMg97pzSOBNr
YzXUm4yj18XVKpwrtniaNsN1a+20sQCrppN8pSfXSf9i9mjn5eV+zVEjpudYLFt5LIJeIbyBs01a
iFmJ35E5JrKNrulzrZ/i3jBIlEBx9oGKHB8+9BQ0sxU9AMiOr2fb1Ez/RniNAGgh/FRVf1egRMMB
Xt1gkdBwEWR4yMMCYGdNE9OmFlxDTvOEU+Tu3gGFrZ8w52LrhTCkqBKDfSkvgC0jCmaa9Ge3aU6A
VoaeoQppHgi7yhsS0jyysahZEjAbWRAKvXPm3Lw5otDVE8kwchAHjRbXSrbPGF/363oaiHqhRq5W
NMzLoCyuvFLL6/14ljtIIIR9a83rbZwZ9DZFrGZVgL4REFjLjWI6iv468gMlut/oBEt0ybeXSeaF
3G23ZpSoixzqNaF7cYQUmaywgSthbk83wNvRn5Q3Kl2RWHw6LbBTL6WE1YWfxyDZvmYJYYZEAWcC
kEPu0YtUH61a6YKGhjUz67A2admJYbPbRB4j6W0ZgvXpLDELsrSS3IR1NCxLxNSs5r4yMv4Sw5Qq
WOpAScenknvw2HjO4Bjhk25S4Fe7NVyGQoY7TaAImKD3t6n+Pbbg1E+nubUev1wG290V0LFgm14g
i4SnGnOLb6AMxvdsqUXMbDOKR/cP31J0NfD0JUiyJrm1KQoTjjicBsn9KanmDhFlJeHJ6ROdkGeV
DbZFquVvk0t0N9BCOGTA4OhOwt7WZ4/hKcN7mNaA49QhQ5SrcS12716+usRlcoN3oT0NJDS/GlJG
BFbJVgs1I01gwD4hYx69B2piNeJ/OpicDtaCCF8mlxagwfc91uAVnldmrsu/ZniMQSr+xAjjpe3N
5THYPBbXGF/wbp40JCDdLLv0YPBsREpGoD42s70tYo0nlcaqQeI7Sd3/NgJJQ094LNCVLn05Mzi4
2WhuMFIN+wKvsvsNzt4cFEJ8Upp0Z06HgIrAxltiZBlhRR17N360Iv+pNaK0fIMtVYCa8ofI83mw
7shh7F+U68LCHxk9ZaTUUjdUNFD9cz1z4JZOZ5lO3+t3h6tsPfDIvnTPCPofbzzKKe/JJek+GcvQ
JGQFmXX+oHExxJ8dgb7T5oWPn7jYDop1DnCEBh/u7EOhNqXKQ/YaSYiCckngv4PB5rm8aK9AYvyQ
5MljHdHBf2QdZqCGVPNcdBhvwkPomeUD13aEN1vQ4Rep0QwID8+PPGY5PXYNTvHMAPHs214AE5ZQ
CQXFDGwfB06xGFzPKWxOnm8wVt+9bpgDLSmEhnTS073D5KTIDVQje89kQTxRaMfvltqw7D5rGW3j
zoo56RoxSV5CjupPqL6r+LnYtbnUIrnCujgI8ywl+SPEq29ljNmJz7Ib7SbRNR+Tl4rw+z7/4Yja
7AGmW1v0yuPYQoLX39/DNmELma67E4eTuxYCF+g8vlNrpdG3Ua1kI4Z62tCK6aYWDIvfL/3+II3T
ndFBXZEg0ZRHUYmluMPuo1elQowEtrWvX/4MamRzDk7bDQln6QTnAD7XTgATDWr7sWHXOhPUIMah
FSFBHRx9xX3szlDRZn3wf7pEgd2F/uctFelaYyroPid7hWd7ruMke8qnrJHbA0I8sYoqutEvIDhI
P5+o/wWXpnZLF8W+paqThQ+JcqCquofT1hx3rZQS+NDgkUA4JzdDa01iq6Ih+fXLiECgyiTCNSZL
GZO2n0Fi8fqUex8I2Ba6LODba8hPsCY1Si52UWLLTs3xT6LPsRe7zg/0IoTWRszA2jAt3ohP/iTa
oJ4jzLZgDHSMDTEJsA57yQW3CcR2QHGjSO4UXtJsNkj7rU+EheFPXjIWiShvNEtMEpdXSsD5qsVy
vHizRYh+zaAhrh9hMY13bXC8hkmTPv4SyYLt6yota47VawtVjxMlPv4AHoo+0pauqPbIuWvsCKZ2
hhpn8BZYu6ElWaVRbp8kFRiBgQPAjkCca5/PBh1Eni1WZTFWiedkEVVy8QLGYhR6cAJ5x1Jan3SN
619KABZi9wI917ORh+gIJFtoyxxPPbnGfFXQraCHzXNQh63WOlRewy/Lr/wO7fzT/OaYS8O0fx+q
bNQTCdnDXjIdfnEgu0VmAYhFnTNiAKoMajrgx3j4r3Rul6tG9/cURySYpcoCyuc9pI6af+5GFESI
SUgCENBtNvfjzKvMi6+J+t/UtMjlD1BWoPx6frodpS8Meu/f3cyrsY1nBj4xmCHkZtTMFYdWYp5n
7eLGrd9R8Q/5/91+0EeqWYJd+CL0TTwwF64uViYeDGucYiwdj+qQUMthhR8bFS8nfW36PJ0N747r
HvINBp6yff2+dvsPgrvfXfP8zy1Xj67UYjvL+oC4B3OdErOGZvgF1cgIILVWsrXPbFhFCACVZ2L1
kORwWCeo+Yr1Ya2QHYIia4UT8pLFiINZ2xmKQwDKt7m1xDSD9xHDpeK+YKbxhscWc7W6u79zxDsY
THPYTZ6TN0XYg3HmAvPkgGpj98pLrgAzpF0MsoKx7nj5LReEB5jxYciOCBKgw2cUaylWv2oE53n1
pQviqGytNEGIPO/N4KTQmk1cV66vrbN6I3ro4GxFJAuz6z6gJIWvvCnuikL8GeLFfesF0+mO5Mfb
uZz92zscJ/IS7gQvL+Ukvh47PZEQKiKuoLWwibWEDBeywUp4j8mFoSmYj3/MfjK3H6+EXfUTqL8y
/eQDU0y9pj/v1KR8JQX2bFxwQTEHzoaSt/T1g5ulkzbxuAORCUeoze4XZmjL8cGYEvV0nbP7CA/U
AVOgfZQ++g3woW16R2WorGKPa0uyBi+NDX/goIfuarS2r/ZaiWj1ENAtozF+yZD1CjiBs8C7jTFw
YkYCFXdLow4ik+gmmbur2vMg/oZN6k3UTqEY5ugsIqTls5ZiV7N7lTtYtRlkqeF8Pe2jBFJHNb1F
KVSm6sacQBlgQjl2g/iA9R4GXG2I1Sv7Fgbj6ItjJ2+KArY2QwFhVk8BsoNrcNAUNBqFXMXZopay
NB6+QKL9CC/AgDx0aBciwu2m3AU83kbEkXy4Xv96ua0EuVV+VUSzd2JsS2+0k/SaYp8a5bQ9Ufpz
8fKchYGDWj/0QytLnC/2RpvEUMseqeTRnOPq1h189VFIjhQDe9zCIPtGmggzIu2FBCgxqQPD1VoD
AXR6hppSfOtsJoXyD8y63IfOn62cbsjQULZgZlmUNHqi95ZHqKSA+ioEmAgRFDQTeDm22CkLHkm+
ju4mw4jKTD58qAKFrjMC6/U4iknXNNNamkLkXLtGlb9zQoAgwynXw2RtV1wmzkYYwdyUqL2ZRDdK
Da+q3mX0c0TgW/Ge2vVduizzWk4iGjskr6Kg96bX6FRHq+ga73eoPXTGR0CR3VVl+8SOjSflrXX2
Ky+5Tz7p4xiNuTPAyv7UeryMEr852efd/YC6N+Y6fInVbCSSpYo1SJjSW7kUSOwYHsGtHrrHb1ne
tMYRC5BUhduZA2ERBI3+tDvM2jwTdxoOeB6XvFYOgnzXLUaYKf4tfp2eYdrkYEauh76vOBuXPkVD
mzEn5hkej8cuJcLn1y1lAnc7gBhYrbUb+VJsE3l3RseuzyE6zR7jF5eiKq4xh03AHQ5AlK7pRIR1
/I6tocM74xRIinUlD7c9/iCX8VqWKkkps+ng0BkH4ekDMSPXgNmiut/uM8bVVI5gl45Nsj0mZqM6
xMwCWAGS9MsP7W5DYXzPN1/Xtuv+14AYd2C2RaQWFbVRTtC1YqLCtLiwVs+PLq+d+tCo2A8V+WaM
t2rPEcsjDsqBYjuYcVuQB0s5IvTZH1L0YuUXv0ragvZuTFb2BjTwy3OD2MVJaXiCe33B3QrTcng1
3Kyp2L/90lVjBXKlwELgae4DQ4NZEqehQH+aUjo/Z9UZIZEo3f5NUg3nHsb7jGR7pnKtF0gTZxbS
rqFV1SEcYtRarSnKHNKYvBNRzWpBkdWt00ZI3Gal79yae7j2kfY2F14r2I4UyHr080bVNCgvtbS4
9/xgJIYLwUTYdkP1FX85/AS5vvmrudacn6EFT8vzPzVfAHu9dNk2T4v25l4OWtr1vMKHjD9wXIuU
F6zdX7v+/nHTLAx9N2NTfRQHTfI5TLMyhuTRC/iYmzR84bmDZgYM7/CP1pUBL+zbBOJGtpVjD0vt
ZmhE8UypxjFl9cjbJ1xLk4G7PV1khmCfyDRf0fXvMbux/EQaHnIAt/6EDO8GMAs7vKldOsYhPx4k
VSUksAAN75hKk5LhxkicX4G775795cg0y4wG2WoAzgVc6JgOra6AxvB2uDAdmeP+YPs4k0aPMyPv
c7f2HlfEfAIzRVFc5eQ82ORjHSt+ZnGkgLQnauv0NK8A8Tg2JC/4+RK0lrjHvO0xjsntLPLxu0qu
Vi5F5zZtH1QSyKbBi2gPq3jRMuyCc1KTe20tBONwVFPB+2vNjf0Zdo4zEvFHwRoyTTPaMiMQ4Y75
k7N/G1pLKfluxozJjR4iw+xTrAi/fEkhooic7ukIGlETUXyvuCDoNwcqmKLckLHWLyAh2IgFRqxI
b6TD0vHcn8b25q8gZk6mrkuYsHXzZ4P2nB8BOG+uBVTBmniIlYSjnRWp8+xujD08QSO09rMoE4l+
bwVC8HZrJbZBGCs5LznxSR9meejuqpe0CF86CaQuK+YduzQh5Sy18nfZhSuYkPvOqs2R2SBrkqju
1ZnHGFIjpy73qiI/pPho0FCufcHzA2anbV/6ejS/QSU4fqb5bnJmymimTk8F/wree6i5exYAMEQp
qSDCGfSnnVUMwAkho9iUoI3AcEXJjm1c7vUcd/wjj/8826o95Jq8DU0RsebIokMPcGOw4+H2TwJL
6arMj1AXJGXng7sRRdYFZ4jkMLyVHPJamfa47zhUlkITvkgrmHdrMYCTYX1LD0Z/nv3d/SjsmUit
jNRyvJz2QUftA1dCHYmAPJs4dp4YpNAjaJnXWtiXplmkRptDjc9jy40YvG4hd0axsTO7y3MnmXBT
TtDFLXGEmzaHpMM/pWKbR2FTtP5lWOmTdP/OjyGuM0jBUyhWFa5DN/1uc6ZGz7G/un6ncoZUCow5
o6K48Bt2sF2pzBIsoMLI6VcqplqDF4ceJ/4JT8k9udWltpz7o/kzglCzK+3gCMN6OEZh7PBvWKoc
Omgx+oN6d1zlGBFLvZWKjF1yG+/2lUB9lAoWxSLYNhh5ZM85Z+ktiYRu7MDQ+hMMEdA0dSEh49CS
JZ5bHBY1y59PsuU1UCsqX53L/GpTxqX1z2xdXG0HuiShlgSAFH5rFYZs3rYLxKz1G02Z5w3LJkEf
VWiiHstImUtXhulqxJrg9NM8DLnoOyr/TpfJ7A3z5cXZoKNqeSH42lC1cs9jJHRuTP861kh7UlFM
y3YfrTTRrBoNGizxaSWu387HBLz01TJ+sQv1oTEN7MUJddD2CTD/4n+ivAPmzxc0eEwUjn2xo/XZ
IMWz/lY22+cQlkT41Wd8zSQZlp8l+LTRjaOxLZ3PiqsUe8eBuPvYl/Xd0gxvLRJ+VRVahVrwzcEK
aoIyNXHoXk8euMbWSudErX94WojpUH775a6ALDPXS/Tp8HQmSlvQ2UzD2NAZthTAUL5lPbB7ybUA
g7+zRnnp740YyzW7r+25Xvfis6ihpI6lJWfwVYCXrMzMGRU+Uq1SbKDeh6x0+cK7Q78RSSoXlJ0L
oZZQW/g1AYJbimp4BTejuBqIQD/a1LD676tpNAkhn1Ccu70xbn2a959vyeeNoYdwX1UK2GjH1iTX
SVmHuRivQGOUepOh8c/iqtNicWEaPG9mSmItonl7xanQ3j9s7wdDE946UggUaYe1npwAm8GDacUK
QRKHP3hiAdXQSe0eXPz3Fgg0jEJaOIg9hcDHGGF46drnI/ZPe+pFHUhlJOFW+YeIqgyCPdMmZa/7
SAirId8YjuRBL5u1dv83ms522Wes0jubeYMHnfRUddfkx/zBOR3Nx7td2liurC82wOpIBvHRlp9B
X9L7AsX5/vapOXrS3n/z/D0SlJSlrQiH7p5CXW+D/hBT7LNX/M+TsAdIv6UiU8q3DSEU4pSTq/Cp
g/Pl16ohDr3ekjfpdH0irkkShhiRSiuR3PRvxI77cUdWlY0WGFk3OefAtkHd0xxQDJHD7TzhTDo7
edwen5gzJPXBo3UkENAu9/GAYxTIv3ZSgqDE7tHIXBROJNZ4PBQgq+wfTI3Q28eF2TJiq+SEjo/l
8otPUlj3W7qTCbLd+lAMHrwwyM8gM4zDKILabh9eClA/f5+6TFiTYJBzLyrC66lq0nQPNR0V3iHP
g3VaDFlWSIMZYpqnREoPMOi59SmPFtwcxI1z3Cf26Ze7mozwm516q9e3bfPSxslKcUOxSA5BC+R8
7vBKz78O7EcqHhXiGCeXBec+AqfGqght0qMIHKCNNgr9jMegDR/GQ2w/CyEbMAXHDE9qPnDgWbsH
UVp+cjWBz38P+Y4zVVM26pIZtNCbvq+bPPg9Ad3gWMC0YIaXlKTtzPM4LsVhV+9ix8w7wFRYzW1K
VcscjYZdK0JF9pjckR0vu+MArHFdk6kz3zxZ6bHgENSjTldusXFvrrg6O5/BEwntSRZxL4j04NBQ
4fKX0yHDs1Ub+R8gqfE/XDlul1QC+Y3q9pYuw6ZzW+moRV9+tN8lZ7Rw4ch/1GvEy+6cMUJ9Z/HF
cMZyeKOz15m8xLWBSv0ZqiB2BFRKc9DJ9fSRa+a0//ssFceLEDNGIYXQ3FLh2GA58+c1lPMLeTkm
6enhlVU44Vo+8uPpCOc0gvTeszm2am6xYgu29SEVO+5n9L+mPA+aPZpFImYRolUaDr4pbqzaZd3O
cCqgbGk/jCplLjwG0D3DxgkbDrofl4JBIKtp0oxJDNFhf2yqmChFyHAtadL1gXFa9qR8tDZcJ2Nd
c+LVLd2W2T1BAuoGbSSzbMywlVPNplY4ZNsk06sGzX+7E/8uv6TW+KhmjDkHmY4+CBscoKi5Z4ID
REmyCqFftHoDLq7eRNaLcjuTWn1rJ7uVpI6GOSWJk4PAXBDVMz8igg3IoU1n73PJpYCxnh9t7FW5
ntBXhephEnisHjq1bSm0HoIRUHCbKS4pS1p9+v30E2a6J7FmZ3JPwwcEGjcme2m38ENu0/cmJWG7
VABiQyEe//E70EN8aVdMN3ET0Mq7hm1iwXs2labPFERPLohUrfomcts59rKt8klAPp8WNJDEY+cG
6B/QpePuo2F3t23k1eLLkCbXDGnTsqgwrGE/gwvLBcN0cAw5TKlpQSRGbHHtz9VdGd43bc3ATa7K
59O7NqxDI8ed2i8kI0v5h4vvBVqelK32SJDNS4El/oXOunk3GRM/i4eG2ZJGtBxI1zHFj0NClrxh
cL2Zg/+ZpkQ5fx427ceZ7OnN4AuP8VtY8weOLDLydNAmgqtG/G3tECUl4zZdxJuPyIIwxgyTustt
vb3t7AEpFe9CV/AC+wwe1aCMm4QeFyEY+O6Gn9K5xBUX2sibMdevF5Cd1gJZPSgJ3NIPg0CJ91v8
kn/C5GqCXzW88+pEzMGF361C17n+540YZW+0D0CLpvq4wAulENEJTgwbCQKtgNhj9uZJJ56uZWzt
xNsDV3T0+OcRSO/jv2e6P0zHBuovkUsfxbjSoEkiNDhLAKbL8VDsflvgspH385uO7uYSuf4wRLVF
tn2w6q67hrmuNwM0HnV9HjmpF7ZeMn9J3KtzfabZZp+zNkQtfDMfzoPe5qPU4RmLy6BmbJFz5FHa
6ueGwdZ5wEt6f7LvX7WX7U7Zv5mj0Msi2pu95oW/WwUppxDfojBMT1G60UtB4TsIYzFc1q3GyEom
QKcLwhpNdGavsDMThUNhxhiVfrD4aC/YeI/ScITDjTQS7RsAMsS6owo6APpOy10nDMh2Yb+a8ZXc
N+tkHS/ikfc3JX5tuMO9zwf5nK0meB5QKYBeWy/GdDyBPCmnSMdgy1/auZzu71nYROwQiLCCPPdC
fj5fWFMOa7KXOR2XZVxLkPJOIt8+lG5B/ILiqTwo8IIyvuXri4BCy7WKnQE6EDDX8fhP5RUk2wzu
kVLKpIX9QBkomMjcHCsn4YkImWZkjKvqB8ZhVv9cKmizRntDK7D3bfaGywz0XM4f3haOQQ/NQj06
zhkN8SyCr9QcOwYt3LAW+3Rjlga2aJ0B9wZB5wgCnkgOYQbEu65Ji0TgBJx7Oxd4xnNODNR8biau
FO9pN8/OQ7ZkXMMngV5Ah2RzO+vvdCmGonx3mWkBKdqtH+pxmtT6e2vdn90Nt9hvGzdPMWnUz86A
bh5OlYOj0cLaFKYZv27SlI+jjTJUW7rq357B3XX31GjLvqvTxTjrqe9/3SCdqrTWq4wGpIH91zv2
rDElIumOU4E56kBHwkhZYXSc3Dg2spg/Yi01VI6SaiZUPwTDmTk1g+hec5NomzIvR13RIOqsupuV
4JcTmHaeotVdtIQP+iT7rud1F78PzpkLpCBJNHL85IcJT3iT2l2ENAehTMUe3O6IQL8tHovO4itn
UQe+wh2vYDGlVXkWq9d/AcJGxOoAUCnrIaw9bRKZi35kLlhl8nYu8jqaI+FiEylC04wvLJft5Cci
aMb0smBiRKpZGBh0B6FIku9NateH+/8v7PpFr5pehEryJfAkC22Tm0uxkvS6BLlYnEcoxTCUUj1H
A6JZ2/gKg9vpMLOFfp4zfCo8fMtgZBe5dBnI2LmxJRn4StsbuhlVeM2ZQgTFVgApuDenfe2etQ3Z
4qpKSwCHIe0Pb//84uSqoBddQ5Z0K1I6MBFMiefr80sH5pOO5dzR3KPymLAOProtOF4ZO/laUyVN
VToGOBW8faMgXc60o8JdkQR6XK3OTirAYTScXnk0Df62G5ssU2N0DI4XMZThW+cSM9VHI4lHmyMO
NMGZOlt2peFw8VNvTBPu0AgC2go8ge4FvDLnpO4g3E6nDHeW8zsjRXXxEeZ8jBg1is66OlAFHNt3
xbv0jFO+zc4/5j8XWKUfx3YDpltio61sEXaTIGN+EBUcoAM77xcgCN0Yf8R4Yw/sSp85VM9pSCC2
iX9ciilotSdVQtOSgl70Rob/nAj8bNNv/yb6J7bU6W0PLvqf/QmB5VCqqP0klG+lut7wGrDIYYPd
zIGIm2Oow0Vc5k040sIzCmjPkwDuP7kBoOUjML0JOHLtqJWTQ+Kc0zalYjlOrgEKsOEkussMJDMl
Dg44p9iJ/XmYmcCFKPrV7iPnGuUqnxq1BcY1LcTf911tsWYfsKs1+bsG2q8pNYF7rbIik3YwVGq6
ggZ7WyTUZNwQFs3aBxhta3U5kD/6EDd+/hE2YhdzsoWQAceC4Y8JboFikDvhSa7LJGaydvCBKka2
HGd4oVjjckiXmAHJty5iBs2/DSw+ztZmsUhvjm8Wp5E3bgS2pTyXViT8tI8ywHEL0Kv8wE+c9PNu
u8tCZhM3N3Kt/tPvbOSc1nWdvKJybNQe5DvQU9+nYO8owPvbJROVTzLoUf5QJ85I8ULBlMM0wF+F
Sj2sg2e5I6Glhn31F7LCjJ3pzagqW09CTm95a6284f2JJliFZbxssiODb+VEt6hqKAfOxl+C9Ae8
YSPu1Rb8PBn8CxNqi5UbNAvQQbH7pL+gIkGP+e1a8vkpZeswKg7KDcvtQ6uBxDYb2ar7zdJl0Vja
txD9dSGOBD/xIUipWfGp4fhoKvvaSVhqwpUIwpBe0wY6gKwm4wu8cvo5w/Pt6PxDDOAAjwoplGhV
qmmlgcvWtAZ7sqshR1W8t2N310hHbQDnD2tHJJJRtVAVJ2sO6bsA90NTVpK1dlczaQreUip0KR1S
ysgwWhEoXINx0E89z2xqXZj0pCR1/I0e2Dz1/e8poizsprVUUjlkPkVOmCL7BH0SV1o1wYj0PJm8
PatJQ4pvpxatL1jZFT9wBn2sQBuskJUc3zTeWc7VN0qnGVXpy5qlIgwl/PvhXpmRLRDQmOOGhr2u
pqXE2CroX3COMWLJ6itpgcPraQjl9Wpk53/bAb38eeDD9N5g/ts9sAGJ59FZ5qprtBtFHi/ggWLd
SyFEWOzVesYAyiyu2+zrHN0Pdn965rNNrDA8IXE2E39x1Op0Lk4anbsZPDw46mJYEYV4j56SMLqq
+Ysrn6hfHOLwV3VZY5DRRa/rI2YIWTJZQ+Zny+xDhpZQOIkKUyJONajHM5KA7PmBvXrJTs0XvCXZ
Jz022DiwNbkg1MqtjZWx22OIWRwucrjqBdwZ4dkJLhkjcfkDe3UuGvo31oyXvIhwIlrChL/i5k00
Gop5lA8Kqft+0Jya4lQ8YpaUkyKukUZ8vlb5fP3ywytdkNjsIXxB5IhWRbnrhdoJ9XoS67Tca3rE
t8mW6z5i6LPTBBm08jcZtCPFrSfgk2wetHUuuy88BzF4XuebQyFjVsnGJg8ThxLzLt6nG+YtdpG9
rHsW3jNBW89FjH1pXXM57V3SRCL1CUyQVznaRv2BP3KOy7yl1stNB3j1K25F7tl9kajsCUNQI39y
EscLOfWLP/Aliw1pDmjFd0yG7bHJTRB9/yAqEN9EaGKvwrITdnyowkOj4Z4ugeWMnxzRShhSNGGv
0op4Oc/xmutB0qjLPaMJiJ2SzAdHkBrOv4ID5hj35Q4ncGBwztPSkM57XDbabtRMMNwZ905qKyMA
B0fyhX+P8k7+6a7pKJQD4yHz262ilobEuu28dyR7vEkfYNQK4cvCJX/fzUb146gAfTLXLCJZOeiJ
rTcgbFIhnh83g1DeCkshHY2V21dgjYTyXL18twzzuuE635r+zAx6YqS2+oQDoWk0cyD6MU8rsEfs
OLAfhoAgO8ALfAuYIhD1SlWgKEOBp1BA01kPIG6W99HZBZZ/8uG+wdf9y9WGSWC0jE3ey1I7eFuK
Yl4ojfxAt3bywpDL3KGiCXBPgpRY3nHec/mmzh6rc4Z3TivPMOWNn7xRov3east/gGoowrGHtYLo
H0HTr23pRU5AyeVENGRMPLlolnXlN1PSOjuV5jf5H4Wx2WdmDkvDS3Dac1b/BKZoc6W4nC1dhF2a
MG4bs5wTMoQn1OW6wUJosSAUzzn9pG81z9Rb8L/F2JXU7au+qsT7+eC+Sm85YOFMAokhcO9ZF1YV
Sy73xEeNYbcmklumdXvF+dBBAvwTRtJURdpuk6tcMXUBMptUCucSDN3ufKvfXIFvPy8fWrJlFBrt
RoIT3am1TdhBeJ2iTR8WNQ2qK1DPyGIW3Q0pohcBAdl579zEXjTTaSQ/3P6nogR9Gc8M1uUHxQ+F
1BgdRgSPhMRKB3SXYgZ1xRQhX7/rhi5a0g0/7KwiiOXXU6AMZvcjZ5t4V67Hlpdz7rGU8GtEuBZv
RIvNc+tmzsHRf2fn6uca6tLlLQQV8T9s6LBeKmtPkBXLe4jm4tVQRk85No5z7h2nFXSbmm15Pg94
HtRb+eg1c/4YdruSBN6cwqykUeW8nMT1rMSylt+0Vp1pPSPIWbieMAxPGyGnOTo3QNRC9CYh2HTV
AZXDmy1Vn6daEOLXPLXtAj3XMALhKjb8JYp/Vz/rne8V491RM/JyZpkOscCEC+7JyV/+b359KwLJ
w6r1mW5OqE/7aKymmvGgJbfggVW9qQOThJwLDl8rkBvr5vdENAUN8AxnS+jpcELBXNq792Zf3pfh
qFq67E1D0RRrpsTc6qJIZjZp67WcAvgRs9Ruxa+kttQ2g9R+1yq6382XfR2lhnaig61KYksVcqrQ
zBH40d6C+m4VRFTwOlAgVXKMkWuvCYT0XX/ygCYDTzYKhwQc0Dg2DleL0/cl7jJM2W+AbCmz/EzY
k+gBxNWUHFKNAN+ROFTqOWTr/RCWl9zPqNK7SZXiJ9RXhXgGTeR1CnUdUajgo1g0k6t8c++xWgyL
hbB8fwYmFLAK40EXc6YyPJQ3f2kj1hwYkYhOTUOqpIQV/Sa4KeQcYR/WDcxvdkvviuyPL1xxfuqC
bZbNPm5w6zVO0/gmGRd1iZy1unbyzHL2uwRl5b/dMSJVRW74j89AtbrGdoYPm/jf6D+rB5Q7PDfT
4g5YtoH3cfKdKOkVS7OAhjw9YZGi+BPKMMGCQv7Qr7lsnPRNGRLdz24hn82RDF2skNQtasDHi1lf
0CAbo3muJUbrRhfk2nHCtkYTfG37BjnvHr5bfqQYXuDrYAhLqnyaehVhW8EpuwAKTvKKv4bev64J
hCHOtabGcKbsKAUUZyjfAHkO27/YF0JjGH8Wqp5JMNr5c1f5KAO/c8ciHLqlUeIMJaji/kvqFVPB
apg3Q/Rhv74itkBH8UfOkhmleX8xQrozk6jleCfjjgTjbScJZaTtwaQN5kkM/h5bzAYp8mN4ilnN
iG4fglj2SaN91eaOolOc2bzEKftOisG34ZYNWmG/5H4hrsW3j5sn79sj9zEMnpw/kWCCAsfmHQHm
+ziXWe1PlF1TsvmSIlt+UvKF657ftRUn1xEaauSFlkMZAflR5ZjszNR+0zLfPwD233bJT7H/yy4t
Vi8qRCe9KkAAoJ1rFh/1VXUf3AkItfGPjVyev37vo4SksTuTT76Q9KszAUx+lTQEghomgP6yZY7G
0JoWS8QtSZu8R63I48eo59+2+vU4bMKy7meVQXbp1T9iINLImGdBM8M01Hlxw0zo3JlYinxUMip0
EDHdHb5pYJgdi7brAG+xlSIlbIeFdjLOy31cw0Q4SlXfg414YpoaVJ2VfjUYhPJBPAP/RZy5vj5j
Vk6/8dQvq1V+qzfCgtYiS0uDoWkF0Ti53CJLhVavKFlo5Bxo0+4wAADqwb7rw0Df5O/9bi6esXKr
Ahyd3QzQZN4Qd1jzYROoNGb8Y+HkXAPLCRxsu5PxYb5kBApuhMRjaNoHFUFlfaF5aZvikxVGI8Vk
bAshXOts4X8fjtmGSvs8iMikUDi3mfg4insajC6pCRU3MvHhJhQbJIPY0tXrYlkIX9VFxxEZfKZ0
DZfoZO0eP/97G9OcYUCOhobc4ppcFIE9d9dxyShecVA89EXuddGFas9eAXLAiq7XyNpwR1km4GkM
cxYtwJpuGHeYqLDzS8NZoSMKN0AWJT4PAgGFqnVOEpuL/Bg5QgFR+3CQW6OJeXE4nDvJJrisLUWq
EWF0xTFZWteERmlCEbxV9exVtRAoWz7bKCXQp/PqUPU6MKCWomr9XyKnRWraG/HFIdAGFuAxlCs2
fD/9sTHqUlLJs35uiiocMDtqLEmH209xf0DExxeW7izg0Si7gEZ1oG0E//ARb2h1tSZQWbs46Jfo
CVbRecu99S8nZihsu0qATeDfluMM3dqGuEekIZK5L2prIPgrLHsgmEgz93jqcS2WYBx12khng69n
nIOTmQ/xUOEqJzMMeoZlVym9SeopnMstAa4STdNCLntsSqw8Bh2RvmjEmzEcWkFn8BzIQWhmNcXE
SjnWvjI2Z5PEarBBRsLIhmGsxZWGapwTom/V/UOz0a5VwQpXBlhCMKWWZ83JGEl4yM6sqJrSo5UA
FanjDIOKTsCbr5H9NLa5gil+pRxyJRNyUnuib1GvU9/9f18yW9KXnTcrkTTYbkCQNrizdcjFyu3q
wyMhpLGnzwMqdu130L6ngsgPorwCdnREsr2AY0KvS9bD59gqYv5Rigdp4gnOSy15PxPony79+B3P
p/Fdm0anhWDPihaAzuQfOxXdHpYCyfWd2ShVOGSmRKgWP6mboi1DcmF7KR5sdKVlrtpazP9K4PL0
JSNai/MAAon53g2rL7zX+rklnAv7fIPtbjTzP8glE1LVMPwqvHp85DY2OlVjftOcR/nb/6W9E4h2
FwtREIvALdsNhFqEGe/g1JfGx4hGEfB7+qCiVnui47agucWJ2H85xH4t8b+A2FSe+IqG1AV6R2nj
vq7D7gAIrr40Yhqq6pcM8nd1jczyyTGlVHjYcFj5oIEoayNYKERMLtOzyDeozz3sMxzvj73KhUQy
UpJeZH7HxOeqv9UDGOudZprZtjUufZbelR+2TqCi6WIRhyzsnJyBx3PFGkn0ibFI8INPqM/XW3YB
RQ2ypHQ0V69Z99mT78A1s3F+g7EHyUPWbIIvfjczGvZCNQm3P2+I+1B8aklOADHyWjgwMUNxy8Pj
LRvtCTJIEdTSgYhd3Muiw6IGOCuzMMZwPWbLSRKrF4zo9lo11+JiuPrMNML2b0YLIOYGSsUPMpUt
JYNVf7k6OiG+IDbHxyZYnK73m58OdLor5AssexIPsbs35jbon8y96PDT9YzvvZjIHaK401LxUMXJ
fyN+mv5DOtRgDw7MfRnU6CCXOpYKMQPkCtwKVqxZW7FC1E6i9pnp1z3FgE/esS5s5uPu2hLPB8un
sZP1TqSIHsxWmHg1Y6l1VDzU9PZ9nf0VCQLHI9QXNidkjtL2aJVR+xjV1OPcYTPUm84S8y43m7/D
BzTmbVANDrAtu5iGxbpxkukRMKa3nFv8m9DeHxl0/ufgRdqbloHIqm+Rs1egV8Qkq2kZt1fUxiIg
yBlmblsB++sXWvr5rjTHO56gKSEl49Mhmnt78LQo46qxICeACwSprdpAA9zUwA20kuvITzokRcQe
VYFrzJf7sh5jsTiYCsklJjp99p/aV4FYRxKTT03fhP6JTb3ctekjDqNq6c9/TC8TJzC1iLT+3SQM
2EH+mc+QYyiM9rlBAzay4xYFOmAf8QJAy4gHmkGqU464QF6S4Z/z7a5RGv1FTr0KVTkipjGQjEYt
hMF/C+Es/x2cSqhKfZfJuKqr+tWbdgMDFv/kGBfgw2MHx+jPn0D47KQbRJa86OTZNGdAfTrML5SA
0UjmSfvEPn3psU1C3UCD/89BpOA+NXPcp9o0D7lljns9f/cr4YTL90VilqjQbcW5xC9NXCdIj7w8
GjcAHCpUFFmkzWloAJN84R5503OM5ywOCEBhtnewhGBscwR8HBI/3jENxIphKCIQBD3oQ0A+aIIc
Pgz/44HSmdbbuYr81EfmtSGfLyuFATx7tgId36R/YAn+Fy6bcmMGYhTkqY3gla9WDkvBbp+2CtJz
MHZtkqjns1D3alDPFbkZbyN1sewqLsXbQL946HfDoFfxHRBEDWVvsE57rYu3kBNK0mpIN7lhdD6p
2FjtixB+1ZfvX7uwPhaoI52s6BVHpf9Y5YOpti7Mfzr9hmcq+s0qpTTs8JtNM/1BPEcuSJJuBoJL
ubm6UM95hI0pHarILzbOXfBEtGl+CPGxaEsX5Joz1bkruB/8qwdcdVoXp6GPcN4hnuy0+XPkcF4S
cuuEkg0WY19BtFnM2alyvMq/msZzOXbhxPafY9gGhq30NM1/kel4NsZHcly3l8wF6p4lMOKYrzJ8
lrl4AQZEzS/LtxDGvCl8YEH498pktGQv2g6cIQEzLOcyMn7zn/dQc7gyer1DAXjPfgKwTUAU/dA/
lqtZ5NuB4Eyg8jgoA1yi/xNlOZcFqD9x1onIbCM3gBoT8BfOQ4HfBDGL1Yyy4oukxxwfnCd9bXUS
GK2AvGue8Hf10iqv7z+tQCTlch6FgmtUC2CVNkZzUhevRBuCAyI+zUr5QpIve4XVjpAFikAFf+OR
11Qc1D2Zc4VskWU1CZKr0T+OuglUEiYvTLNh9ckqQmvzkjv1nkmFr2xIatF2i6oKCs/OULV3v32S
KW8/6TvrBm+nroItg5y7vQSuWQCHh9DjwNGVDo8iuULWhGk58wiIOlGVXPsrFI8GJGpblQIuJDzy
1JEcrMTn9QVyRfwuiZET8xBjuR75EsN8u6cpbctLQj22OEknbUhA6XQCyjjFVmjG06uElYaJFOHB
ptHn8OUEdCFEz+uYKM0jO9l+kOaYGo7BkJkzC8L1vBsFvnobUJpc3oYIu8oFOmww3HinghZyi3qa
XLTsdl+HCOpNyu83reL3n8JnUhR6e2rSoBoVd0Yfs32pk6Ev3q680CKlekT7lcg2PUnd06UWd+hO
dDHydF8qf5XG3YkB2WHjy3F8YtTn1wELM36B1VyR5jiMXEE4XJh9rMBjgjMEEzimIH3Jb57w4Xlz
R1R1VrVR16WmPgzEuM6eGWI5LWeJ7yJOKScfb844KdwqjwUCU6mHo8yd66Ne+jumHTorOuD8Q3eu
VctqUZBMlhnYIVc4gmHymJa/T/ogqdUAzVrQLqkLJDqKNnzwGE48NBvgw4V6tsjWQs1XGK3ta7Tp
mE2w5cGAklqBxekRIOHWW+xTTcb8ozpfP2ci+DOj5X3OeLiveSHGHpbgqWmokvuPBWFIJFghVg1P
FJDxkPJQuazbwlirhd61z7Ba0VLco1JcFnEX5oU7RD8Yoemb5NTk6tcienFDl33NQJTHsS9e+0Mm
PM5bnx+7JtAL7nuJz94eGNi58Vb5rB2yd7KJgUPFDAK1Z4g1NPmRZZbHTp+57S0Dhrl8f8mso4+n
tZ8Oux2F7KnEn4Z5UYwmyl+ozTcb+Z3Qz3vzBk5IfvvKG9CVDT/zOVVrCv+BZayaIWmdBO6oOlMf
+dJn/puEhY1qyuX7x+LZeJFpNUQ8oNmnF3XuV05WPF6A/y56QXhzDoY8B7Wxb7iy2eYUXsmDd9P9
K9QNCz2fEO9Nx0ndpA5ZFh/UNyTrmukOsorTrmK17IS7AYAAjPtZSU2O6JM5mg/rWrE9/lIChYo2
If05cnqBJ+9TgKtW7fkNTLyNC2py3x9QQASQcjmJRI9Rgl2uns0L9ZXukbtVlEKqJqcN6cSZE1Jw
57U3P6AM+tkbtLLPlDBb8PszWeKJKTT5pb/CzKzcbitjpbrh/N2IAV/9jL7NzsboHXhtCQhdaND3
UNpiWC4mfawtHfUPy3gK8WmFO0jDDIek2BDa+MMty1bldOGlnf/T3prhgga0E8KH3mJvUJA7B7hj
iFIwNtjAvcURVEpPW+2J8D48HuHufEGEx50xFp6SbWosh+D5kB6IWbjlvKVrXD5gysS5arTDcJRh
7GoqNOVyhuRlTVpHY+TmF+bjhJvUSzvuFkvaG5evNHfedxuh1tWd+gnO4KvGjrAuBcUQiiEeBL7r
WpshCDHAbMnLtgV9pwWtsPGQHZcVgxUfBP484xrJTsE4wDAlYxIx8gjANjMUbIoNSlZDf97Y7doy
0U53bwRi6KRy8nsbGgOdsntD/Otkg5XfjkrYXFPQqMDX1QTNQRxCLQGa5CsWO72h+3MoRm/df+3u
mntmUSIw/9nNFjb7pL1gDGxX1z5w/g7lrFfy0WBSYyh0WVAVESoh5quRg/d4os5Wj82WcZbo0kLD
pweNUYfDguncILYKOHM0ZuzteQsqixZEYMK5vVFn7BTg8HZL2xui93GFAPC35T0hSYnx9YpWtBa8
/y7RVN4ua6b1Vn/9pLCJUHDN1nWeiBlmVgIKq/GUc7OknanBWDMWnoZ1mLx5F3ADiQ9et9FJZ4at
1I8DqJ2v6IQKg/gsyHpLPOkOHoHJ3tBBOGWX4MJEw1sXqeTi6K/NcF1AHoUbMAjEXWlWXyWPBzx8
LVeqi/4ZHNBTm9dCrS9mxX3/eWcooxe6KQoMhKWrrL90muvtl5s8ywno+WtoCha10s4W5gS+49Hz
IhEruvHZ5rXx/NjS5nueKDd0pF1GS4JjteiM5gsyHEKUDR6ff6QyYXit8OawlTChm99TlZ54tJnh
edgPQQLKXEre3N0crrMAnFhHd9GgHlrYfFeRkZADoCkLPGSJXIMMB+DkwCAOSVwYImP373qIdKgf
vhw4IrXXILARIhk8zyojFlHwlDW0xa4rq5mzru2paQB2mAgSvDdMXYLt3VSOP6F7FaGjewSOqTOW
jU59FRwDvAzzZvOLVb+eTcUglvCUPt1NVFpnaxJjLstILGwCC72VXD6M+MwLzPYAPjSXjYvzB4Ek
HljmBTfOQNTrUu1HzCElgeq/rC/F15EHZ1RTnq3isn96lFlcZUwRZE5Q5MHVWy530SuiGombzscY
FeDuolPBWoyfNjUbVH/439ppMk379m2MqA899dtosJnkbXvHvkrch4I/CbWPHiXVqQkgbs5Ar1as
gSa6/Jsqf5SKVT68eGdYXTLR2sbhA/bb63HUMZCM9ZqxkjBSM9vJ7H+G15sE7tlEzCX7hqPSn/HC
PWC1aXGcbS4ZPkg13Aa1CSnt2rPF7Mw5R8EOQY3WakeIx7dMu0PysSY97UMB5ONdWUhCn5t0/FnH
55T3/4cVV+Y29o+gFKbz3fkm8qd8kKiarIVPdTZUQZM53w+XYERKyY8RyB9Uo0kOtrpcc+0DawbQ
3BMUA/L3UJfo2yT+woem3gJXT7cUnb98oC4bzn3k2PIsjgrM+VR3GE/h2DUZ/ZwxUXeT99woBXXf
V8VLsg7TgebHWDlNylQLry2aB38Cy1YiV9k58Mb66f/NWWnQRDF4haElJh59736ROzyjMD6Sykpz
WylrkRE0T1GTfWUruUR73Iz3sRuFRs0PC0PsB9g4axYm0Zo75dVPcZIt22q3bodtp2NChwzlfGhK
+FXuDbkg51dwuzT01Ee8O8Ts4Vg74r0rTE/7jUrGElB66pyQ9l/aEIvydYKoosWkntEJIt7ysVyo
YIUH69NAeMVI5dc+l2BMUz+hrw+lew18pHiWcUsIWbllBT3wt59WHbLmZij9dPKCxXh9FUpParCn
w3uKVUlXBG3KyRQUFQfAn1S6R67pbtHI7C/zkIQG9mkwSfz+J2PODUog10TlmDXiGF0JF09cvhjq
m9XVoGPSieSviSPJDs88mrhPMXYaV8yFsFCx/dob/dFiVXekzTOPSo22SCllDWbEigv1Mx7NW4l+
Wydsqh7QAW2bkHQ8S+2XEBAb2nk/iasa1Zxc8kV6xSDJZdU8gxrRzbxkUMuZK/NElJLlRxyx9pk/
nXi8WV7XdJkSnipzK9s8LnAAgJ8VUkGT0U+2cdpynwU/1vD91XlXy9wbwIQVoQog6rV+KZuXdDal
GRLkbtZPrLepFMp2YgVurwUxY54Ii0nhMYgAAHADkz0M0w6j6xAy/UFXtmUL1wJl4abuY/m78fEb
wgC56nRUnxxZlXuy/Emo+ZfO+XaDv2/syS07ccgXSmdXNFCWwragkjtXpF9OyQ7YR3a2oeVBjFLH
TvxlG2ZXh1TBjkdtgS1NAaYFctcsN2L5WsoE8oMybKFSj8rXj034Q9tW/FT1TJgC0eNIKfpKbe+z
XPNo7W+S6QDjpWDGMtUcUV/2IFCua6ogj3K+AEgz/fFp4hasG8BYWaBtPrjlx1GQSxSaIFATTcMN
tkwz8z9HpSBaXZl4++tfDMFrgUFoM9f6oJ4NTX0Hhszk65gIO+Njr/2jVGHXI3aN8lh2t3h5KPBQ
3rOsZrG61pOqY57E5QCmNuUrb4ia3WsMvEjQPRtCbVberZQxXL9E9LbrB6y8VJVUi+D6D1M6c4dm
mJOyMekn6fkeL72CyGB037jIpLs5hhoznbVk1zvE6wp9REqAm2w4ZbRRlLsEximHd9UNKy71goWN
wNxRGk7QFtpjNBfAivWmSnUM9dua3ftQVacUkx0mG9QkyqyIjn/vFG+WoyH8Sj18xEfz2ggygcuI
xHHX47CLbtpY7u0U25T0E+nriuKeUNKyEKq3TwCpj3zxcKhy9NLyHerk0D3EIgWBCPUekBAxzpgO
fJllDrv/IJB9n4I1l6biHP2dLwlxtgA6v8D3g4rbzT+Ajcsmr2oEmAaS+rosD7S+0seadGsLhe5E
2ZCp4XJkW3YL0IYNTnmvV3A8AMtVVTDXV6EwznDuutT+C2k3AMRxPx80xlEp1Nwxyw0EXPuvVYFT
etIx27EfQdgQicXp4Cv/jAC8zARfuvwmIGwmhelniuSaf7mH0g6sDwBdWWweZouLqx1fDHgDpBWO
RTxL+NpO++gs+7k69xz0ObiBjau62mIHnESco4ucpj1zN69Qmxc828WhfnwEB8v9DbWE2lluYRrQ
g+GN8FfwBpZOcli3XV7ibLqHAL6bqsfts6D7ruuXCNb1saCfpOQd8ZAD/aRZgVGLf37LzxV9iAUl
MRbaFF8LRqIfO03F89sdak8K7C3/v6hLIcu6kAGgfo6ODS2F9FO89P+ePfDWeR0Gi0pUWZd9S85C
d4+HdcrRTRnnLasR1qGzmQEBDYnco8TXJ7BYi1QJulwZrDSNnBKr1P3FJNNyI0NUxpXukOmZbZkk
fZKvhApenfz6B2lCDFEetAp4dxProyceZywjtzJp8qhVNBhMD3xSqUL7ctndksdKl6l6pUfAfP8Q
Me2l3YvTzjRMvVQprCWgbRSoSautmlUMQ+JWBhuykvpTQZx+Bxxt4y92MpoQienOO5BcO3hMKBbS
Ukhh1kbBHRhNXUpabk5vgFBQGfcGKeo55gaNKbYzmg2WJcYy5HZO3DxXhhpdEFmdTBqaxNsiyHXs
xRgZMYASp7a1vMIH8q7cgCosVDllp75AVBosWBU1YAq2i8gy5Aj+zDcPLzbOQHX7rjNae+IMFuD0
M0n1XwMj0m3OHmnUYBL7Obt6OAHTU92yqXBwWHICFdAizMu2q+Pf6giZYUaIpkH//oMgoUafdtzR
47mDF6jVweU7rV4xrJJzNZuOF6xe0FfBuOpxISwopmgMkbWkHQ5JSR2RVMI7rixo9W63WL3DAOIZ
kdcKyT+/w2eGN4NvcTwqIHz1tHyfA82l77Zl2/qF5zsYl6rJvU53vtoH/1vgknBmFnYK7o9Egs5O
q6oLecOJGfhekPDxX2Pf0c+fVxwIavH42KG4tynVgnS2akph4AlWbJtPNRS1NoFr+F6j3/LnTG8W
ZNvzbFbwwhLa1Njz5ODmPZ0j+XQ3kM37mB2y+OoLI9hTNVN7iJXJqwN6+mQvwlh89cUsJEze3lpf
44Zo1hJ1ef7yzMC/5kEJry2cNlYUkzjPbz/r9/MIObQ986sEkNEwQhY8J7M3HeG20Oc5nhqqiYuM
bCYdMmoKIeKRBSyg267O6pAK4zjiCboO4aQvVWgy3GjroHDwRPLxwTf2K9AtmgU0amPwZLvlen4h
xVOzkbPsqhn2OoRt5V9dHIGXs9E6xMAhRZQ3YmnH5/zeSw/U/hawbkZWfINdkr1wb/PwMJyuF5qU
KeMuNWDjYOFa+EEPkhFInkge4RM/His7M/yiJr4itJpeodk7X8vUd88u0GvFPTwqScQSXJXm6aJh
G6YdtBxYas94KhcUgBXDfUmwjOu7by18Lmip7+OgH/prHywyxNjTgsBY88jdzQWK1wA+5VLGCTHe
oUxGdYK1h30/AvZmOq53rbHaheD9LFvlhPVgEgYnOQB/bDdec2tCvnrixNHcVMnmLxU4enZf+RGh
XJenyDIFoqNPakh1UKjAIgDAb9RK4xrJdLr8kJ0cHl2OTUurbEsJ/Ks0jxxBBnGcQ2wVgflIqClV
WbriLmIt/T0XNa0EZl20yp/mEvPiaSf0ivfzzaqVWvMOumZ2ZqhYf6/vV+2Fo0DA5cUh3dV6aAVU
q65uq8/91FSHphgxjscbBsnlXIZiPN5jpBAMX6ACY0xvcE1RziGeFy5oXolBwF1efaURfrf1I5nX
8gEpkfqcjdFeHAQK/1zoDVrhLYoh9YnXdRgbb6keIjGTNT6izkD2UtFJsPbHP9y9PdczkOIY8D5V
2YdfBlkUwUUfQRpZbGaPJSIPgLj3wsBTK6jIBy9ttCk4v9EWhHH5ulKRG6V2HploE6YG3NHGQqko
PsArJsPpDiMv1+JwYpRwl+M+k7WEXIhugIex3ouI6BzJonvdlzkOF4Cdd83sPeqEgP8PpF5DV5qy
Ka0cfPZ8rlg0Ahmo8mEmUjWm4/7+UBCSjo1GWMkaGDhnWsQm+0qvB+Flgzy5RxZd9Myo8L9Anzbt
wm95y0A0/wuskPsL5Es6TGqAht5T47EIxKHkB75dgC64may54Sm/84iB1aqx2Zh7low3qbLr8NUn
+idIX99MBv/UluA3cJBzkpOVT5UBFl9fF6lz5iihdp6NXSG4UFDFOG3OBMXYdi60HuTUa7AxmIVk
MCE76ktNauLMK0NJdL5OMA6s+CCGFFhn02tLTGaSYQgjcbb1/i3poSQ2nY4dy5EsYg9cGaOlbeKL
C/F0+H5QzOMdkXIbCltvzVmGAqXeySmkJNyvFudFk2qZ3f8dJtsYRJJUz/SWU09RBq8Kyw3C5j2q
3CpcD7ar75tM/qXPDaqG8LZvdcm8iDNWnRmlxJUT/CpEoc5qhR8Rr5EnqFya357C9YP7MWjUD2C7
mlCtDnbYGKpE3/4fg6OEmkALSSnMVh4K+dopK4Du4MdRWdeScXubMo3NU4VgepxIktSKA8qL6jI3
xi3p3+n4yH06bGC6D0px7Cg+eC2h8JQ9RRgF/EzOVWlrWscFEMKkGbK0DVyYuKYxHkclre1/YvRF
OutNe1I36hOQ3t3Xhdne1hXRqO+y+Wr0Ck3K53bCkaAMiKhpfb9akkWbo5op3sVGpTDN7kTMbJCU
eR7e/UhNpRbD3/MrkdUO+L49dM5a/oA9ROw5TtBXuFIHfkRQElzcVhRhPG8fPdw/AFj0Y9chKN+w
Ejh5C0eb92ZZ1agPXmDTZ1O+0lJ3Q/1wsdKrEz6smt+TIkw+f5pe7xZvGYIFz0SyeJozYZbRlgDM
pUt2d1oVLYOPQllRBXGB9UKNqw821e8kkgxPVdV1G0xS+3ebFW4sElPF5NaNl3MCL8+0hatnuMUA
GNmafvyl2yXlkHtYEiXWrreQaP8YmCUqQk8e3Ulcy8UlHscKZbip9pp3JNRAn/Oa6CkRbwyQ76TO
neFrpCrCjf1wXtRCABYhopsMxxgy1HgFhwPsO8ig9m/3L9XQ9OlWzwGACCQfkEJ7Wfuq0zMfT0uJ
b76eawkfX8OGjP5UIWiGsWDEY8mhhczMuFF6X9YV12bJvAEEEm6Im5L12T6wPev+lEY2l2IwMgA5
n2C+83+J87Z4pPhXikuyBOS5bour15ZaV1nMx8sSGHXXoqz0OEyjvn62MYvhHgAp+RS7zAQPQ6+D
zrEvjLc8mTm0PERp5Vh1xElXcxDcguQ9CvRGm8doUdd1hWEbUjvynVJcHElEoRZhTxRzkYyjBEcu
POX2jgfAjRg5FOJOLE1NUZhS2OUSGn0uNaNh3om64jYehk44m5UdAsvzqc8nS9v/7mkCVYRG6XtU
f7XSd42+xz5IspKNwzaiRbp+hsIsjPMfgkhIiN2F4m4Kd2aiM2/x/sOz5He1BR6K5KoXlZkxOUK2
yxI9pPGAmj/7rEe1KxvGKJvk/nK6sQ8DxseUU1rYVcQTKArFWY2a99Q+e3Hlstq8CbARHN2jdYru
3HCh2jqreAqxA4txEKJK8RCadvysAZ3/pCm1kwebZ5J98OA3+8FpCRbinR5WQEYwVOcCuvXThvOQ
PaDtHpHexSdlruxgViD/cltTrHaCRlT7Oxjk5ghy7b0iJexL2p5ysqE9u/IvUfgmFj7UPHjABWSJ
k+u2hj4SOMe5/VbYFVuXuz7zPVn7M/LGazd1uIQ5AgCMQXlUD4s6Ms8frqsQlYRd34tKHDGrn7Je
zEpZLKjmy7Z9OI/twE1SMiLKLczLqKHMA4Bh0k1xRTZME0u8WB22RirGeh43h+2jxU5wmgZFwrtx
TSMhS0gepbxo9ycdP59VGq0q7olIl6seKuS128vkbnxtVubciw0v+LdDK7+hh2cNDTAtyYdq+MAq
HDJb7ticTR7rdCMgzsSNn4TWRrH75pX1uND7UdHJY/+eA2S7LtF6WxNhSyM69P/tkuV3V7Aiy6Am
t6d819LvkdGfHEFJfDgTrOxq8RXY7p5ypzi9s/Iy+T81xrY9cVrK1Mgs32x2lxbIyobJ5s+IFfVi
m7x1GS/RGNgmNX64SDDNEjgEUTX+HtEnzziv60iNStbcMPRZLDGJ+lOnjKTpwuXSR1G4pHeCLoAX
76a4hdX95HhrluN6FzafN0sgLuSHytK57QElX7O6sepRz1eAa6wCiF1X7+OqqI+pRjRLiIai6GBl
q7I81csPm4V2KuxWy9I3FnQwqNLSuJ1A7ya+UWlZ1LoP4QijXp/C1lDkYgmCBdbFLXFie93V4lNE
wzgol91Dlcat4UDtfr8fVjRo8k5j/YEo6BDiEuRrB2wkRwdpwjd6qqn7e81aM6H9U2mukiuAqxos
G3a+mKMne7k8tVvOQB2WAYQC47/XX67aQwF1uakNgKvBmLVmWIpgcZB/qv67oxMUzHz2lC1H6r8U
ZnLYsiYPmEO/ro/uBjTT5yH2C3ARo5CqobadUQ6eojERbZRys6rHa20xWapxZonDHAqpRy6tvjuE
7ydQD8coWVUofzKIyJx9RvlG7oEImpqGihTEujbgN3EiEU965/FCeIKONWLEnc+ExC9aXcZEiLWM
OrNF/PqCkdDDf5t+nCPopnXf1z+vGVf6mEFZSCXFQnZ0ty5ZiZXgdFG+/i0ZS03OCEUPGQltIr2/
xuAoMmcX41Zvqc1qVSjPkaCAozH69co0T9dTF6SZA9SRt/gCCvxdBehsZijGdVVHilODRhSpMbBi
UuY8B/bpLXuVlor/sMyOcr/HkBJkKszHBiPBEWwMQic+QVzPrim6TFbxEaaPhmtHpRFpJB/2i5lJ
3/qcVWXu12V+JMh8Pj42LD1MSIL0ZxsVYfkK2+FKYgJTDse7N7BiE44Est1/A9QuDi1BC75StsxD
G9CNa3krLcXVjf3F7hhgz17j4MVcJubqkTFL4tk5oHdJnn9snY1REcsZYP5rl3HbKsNJ7TBfjALG
1Ahf709ob+zfkBEPzWoVbSULdGuspgoRidvyWVzEmgjR/8U2CZKLeE8NVy904Aby1cr6JCNP0A6w
W4mkwILgaG8h55oDAjg64SlAT3X+YQ2vbF9GwHHbPF5D07XX883c7amdb1lsz9SuUu1HiNHppoA+
puvlfiCpJ2x63u2iibPzgo0t/6ZGdo096fGzpGNpEyO9K7rhUyxSYT3pcLku/Pcz9qz4q2efytQw
t496itgouXHhYdYMUIWUHJr3DjSl6YurjKN6JnH80bxqpr4qeY2inDb5yOrm0LUgEWjXr92mp5qQ
rnbXGZJZT/Nmw7L9xFJ+nbhUlLsvP4aWbUQHZuufnCRiFTB5j/zwFIY53ZPgSeDalo9Pnn6Wh1m2
djnUulSGZptpyBJZgGtTQu/k3L5SfrvaWJ5IcImF9cUSdl1Z2wfSUvCDWuxcndiBnnXOVdiSEEzi
oiVnZWfkApbRjAKjwORbQhJ0YMw2K4IqtZmFZAsBUUJpdql4Q3v0X4+p6RIxdUvYbGUP+Uh/R8bi
q/VQe1/eyQLbEs94C/YMDw8yxLfCexpwr49PHTFYvRNSD+wR7VRAjAlOwLT9p3OYvAXzAQ7jBmvP
vCWyTAOrl8W8dhyPX4PSTCqkT1XrgtGFQHh0RE8zG1dYjT9b1hNRbEFYiArmjgcA2fY5U70pTt2J
t81ecL0/4L5X3Y0QCgFQWFYqqf4OQaWgULupJheG0RoO2dN4j7GSd/Ur55oPXZtrkj1PJgEP1qP6
U4vtsEaKsJnvD5boiMYEKtUnbWWfSDqcSmyqtG/barzbJSmcxvvr+yw7dODIT2rzwSRW7GEDX6Qg
UiRiZTPpPngMKzG9iBq0w2CPsszKeD0Lcvuy+ldHa2mAmsu+Nq3Vu3+vZ/SHV9DyDn+lZeEMHspf
AQa2TNObQ29A9bXQPTt9EuPWMsKyaWEvihwXcdqmwNUYaqc6JDSsJKkwB3AGTj3LzVNfwJeHGKpr
ApA6BLt6X3Pv/Ogw+6J/7qlzp9d7iy46UC7xKCo6HgNs5oosBEuKlNSt0JvkDKVisSqcJ8F0IQ3s
TWuFAIxrUKlZ8Pwx5h+poLVi51Pc7xg8eD/m+oeNxDeXX7EqDj4vx3o+pD7xMvFxFMQwoHWS3xJY
z4/jcPXBLhjffjSUxdFpM2pym1N93FpqL4GloR4qC/7rMiKC+C8jXx6t5cFw02S7U1x214ATWjeI
LaE7UvS/4zomlp6KTw7nlzxFXpKYSXTXUp72cPPkvi8K3E/09VwiGWQ27Wl416vnu/69S61g5tu/
QMecnmLSLRRpOkPt1f4zSMRQBRPrwNnL+Q4pF3LqVA2xaLdu6lGeNXcmUed4HwBpKJ0TE5w15ULr
R8WACJCgGcW1CifA6Gb+j3PX1xH3VaJLtq6pNmSnpO2LxvGnZ7WGE33qD3RBYHrJoKy567RjQXH+
0gzP+JpDvdz8+LZ7Bqe3lf+yzeMkyFh52qOIYSwJtKZLHty66uE58Gokm1K1RXVQM01LuGepUAG4
hsQzcNU2rGb4331VqjZgtSgr03eOhZGJSRo1a13gkWy8cfUlX/v/XU2D/WgCHPigCZaeMIgsP8DE
F7mMEOVNgRROhHFZpVdhMFRdef5wsr6RfJQbV754SM2vSAN6IqGoEWvtGqwvUTmku2LsyL7lG4GP
O2LXA1sbsEu063qnqaEvmYxjP2wWSt2n2yhitVpOMHRYjxb9Xf0PkdthSv4uf7pJgaHLd4twU2dl
GYxaHtOB64FerFrdnu1nY317wUy8P/3/82bKRTUTqhzwg/GJxsy8BaQ8myZmQ8a/P+GetX4IimZ7
bNqL8GWCNxTMNEks3OhG5Ja86p/B+hXu+OWIlX960/lAiFGG+y8c6srShWjMRKH65sDjVk6AR4Cr
dglUoWR9lYm6cVQqbTBkJoUw1A1OvWBXSHfjhSL8DFfifyvq8cVDm8zDw2yP59o5rDkgy/OuEOo0
tgrU3gw16Wq0sZuImOUSOvX0y6p3Tw+QIAWtFZUfYo6QsC+XOjFTXYffl7yXR45ClBjDNS2oyl+B
LsSUtWvLWw9I7nIuxNf/zX033hxn5yfIz00OolrTd9APrEusubsM6jLQqBbHFXU4O4nZ5H20Ji0o
3dIp7W7aiAQXFzGQhozjsHJ2xjH7ycsa72b7kkV5Ju55ginAPmrs0K/0R0HajGTCctpzv/rWqxoX
dlvz5zmYmcwzNsLX4u7SAJ/I82Wd2fI6dlF/SqBYWJusdDwp3gmAiVB/g4unt96uVGaf5f2LkefL
8DjF+3sSVQhQULggO7Z9elUa9dcd3C9v95cYiYm8YfuvUFM5Wo8Sg6Vhx5sdNJ6L/yWlMEJMCo5o
6TNyB7MBDflzCk/7RNR4TTgXn0PwC3BtoNQJ9VsTgI9phX30pHzgPUHnosOBVITpHHS4d8K74T1G
WYytv0Ufa2DliqO2ElAQjrSsZFxgqLOdJIHgEoDjJKEznd9pt/3N0pbU2lqDiG6IVBP8d5Dozkrv
BPWOrTgnxHnLp+JKtKa7wk3hFwa1VoNAZbNF60JLtXEx2Bzc+1WhnDOkdHc47Bk/QaEKW7xZZt0d
PGwQVYXEUzw42nBHjw+Gfno91coyG0UojkHGtiRYdJabdYe5f6+ZMwYg2/7wwO+LYuqgVQCiztzh
Kxl3vDWImYdUpucDCLg4bpMnfh9fIL74gWkliNBaQ4Fz+RNlbiWg7P38OV6rtlTtaOGPU7tnYw5u
MLA05JQBwsFVmLg2rJFLUI+pBYQ2KC5Pnsl2QeXWqmcH8WSLB6gSXFl+Bz9wElE8a5s0RavRJHpS
v69SBGyASSqvMTqcEz/2HUD8qjHXjvqFsApIg+LDuHiMws85+Pg/QmGg27pFRwlmI5Y0RhzXECGw
U3GygP3cBESn+skZikO+Q8aXD00A+Y/UJQSJ7xEY8trVPGgiC40xtnENo50jLYs7z5D8sl7iRwXI
b97uHh5ejAfaizhEdLB7NBmcVMev/X3x51SZOCfILaoO8P5AvNoz6w/RtDoEPVUviPEjMXrWyuvb
52XuTgVLQzVd0kv8vnmMgwddpnSgVZ8VO47mHZnyuNJoO36XIkCJ2Z45+/HSgt1/1U7lEzV9O8RH
BBpSWZxUJ7H2tl+zPYi5LHaZIo2DFja8/uOZhJmA2bY+HgV8IuhLfq0aAnXqlhOoTI1V8DA99hIs
M4SluiwZy8gTIjspL5UwUeXphPwE+Qm0dyd6NDSU15JKWQ6lF6fdrCYzC5gA1nzCI7JNLhonTxoR
rHLEFYpBg9psrCy56Ms6UpGtPXA6kvALorqd11fVVkN/L4Ah9vFBkRQ4YPEpyVIrF3NGZfKEAUQR
IB8lpkd9wdyf/SicJSQow4D2lDdMfql6ZPwtOZcHKEZwLYAZaNhTzZIXH+6FRR64rTlCKaPA+IZd
BBjtSUeSO8/rKbXHwPSkRajHUxH9fPAipxUrhkG3fEhR56BxpjSTnGLSUCfXX9Q2RwUcznN82vrQ
o47wxC66/sjkcv5ZDjSA1YZzGEp5ZYSV02psP/iPqE2Xjh1yo3wz4bTFupCH6fga0hBlfxl48cFn
diSCZuJYazJ6Tlc/qz8yk8zPZpuS1lzdkazp7eibQyVzZbp24jjMEX3prIpmnYlwC7a/VdPfKd4w
FBpwjL42/Iezgwa5vl2Y3lzReo5vHo3n45sSbuLY+F2aCeWfwKkePg096uwyjBsiXL8xWJWTr3z9
N+I9FAQboz+Y0DeGh320cI9IgLqaWwQSn2hIUKYq98IxTcTTD/VP3OkTiZvBLJIphWaYeBSKSYj4
5ZzKI7YEH4ILtQBrUpdEv+Jblw/hH6Bicp1rWCmZGl1JlHLldn8Z+guSmv2UtKSS0Zh5+RN4yeyX
81uJyMCQvKTCDM0oFcnDKe/A46viClwhuMAk/EbSSe34lTbxO8VgkqUIUld+ZuFT3RNApJU9aeKR
qCvzFKz/g1faLRUGBzj6RIovtSfh55M0OcfuPrLHES1iewb2zF4BD6jB557P1gOycJDl8LXhLfGb
StohlTZelG+EqvVYaj4x1Rtf6yVRbtu5e2mQXXrgtsQrk67YJzWMWUQhZs8bvbL4hMDmaIOcahZG
E3yKfADODxwnmNp2zukx9bMd/R9I2O+p8e59W42WjiAm/Mwvfnm0p9y+q8Z+qv0bsyesVqKNFYFC
N7oEnPWenrQnOhoXRI/wTRP6hNwAm+iX3icfO1AH93xMGDu86bY/yBdxCp7N+26kIqrQG+XRHTDo
ZkvbeZroiD3LAyC76u5JuAsJyGc3tPKFSUfj71keATfFtTt6WCkd85Um10CGJQra30gIaIfp+VuO
qRN3LhYCfcPgxluYQT9wl1aLXfHsFpG59avo2S6K6k81zEKG+Z5QwX/mJZWS+37hfocKR/z0dkQx
v8DVW+7lJMKHM+sqnx59dMb9iLHW6BOdRdYjn4fVDjXQJp1bRKmrNNJ4fIAyvPahilkl0wH3+4oP
GqP38K1q4dHqN+4ZEhcrBNklB933Szta7q3rGj+pTAj/L0QoxZ6U5FOtaxkP0lCP4sGnp3npgLbU
xgU18VLid5TK7qb0SBIQR0XU7farvb/916ysNEtQEELhH/s3XcRXchy2m/IT1f86CRLkKNNFg4+A
RLZE8ehiUdcgSWBWQGBNFFGaubm1FqcZZK3I2vc0nxgyUCjWJ4ITDGQ9tdT5sbuOYoDo6DjhmX9Q
2AwFXR/17ez2UTCXpdJ3VSU9ZzRxG1peHlxmQAx1SlW7CLbMWep60HiV0gW35lTJ91uxfHX5BDat
mc4GA9slD+5rGL0mckPzXn+EowQNmUvg8UOy6+LWKPv+d22VFBcxFjlvVGN4FqdjOOLv78J3YDAz
FMbcyfQmDdbAgBtDvSf54aMWTJ/U8scT7QnD999UQFASMnyIWhQxn44D76QKAH2PHEU2ikZNSoKE
KeZUftrinnLTmW2WNKM3a8lp18gMViq/GN1hmhBlUBvV6+/ROqGAWZcxNs5Gn3B7SddyVgzIfPkL
bJ365d8Q4cBt+oR7E7pYUI8yRscPspLZBCPbQvgO5i6+TtA7EX3niBKqJQ9DjAyD+5UfBZRzRqe+
HBe0S1EK8Bf38DGwoxnpC5tzTgLZLe8U0z9GgrnIKV618FrxdRFH4n0HGKvRyzGpW7/s5cWO9uJA
07BMZ/zNPmFBMjdM+VF4+vy4aRZfqQ5vU56I7ud7z0V4G/MSqEG8Uvbu8jDLBVlFkoBf0SMIMQKy
zwGTf1iA9UJAwmpO8/v3vyGcT71dbxphmO3WlCowJV5//dttdLMULg38P1IF6NhYCkHpkFcFi3Ml
QVLXon6yuJPSkUpNBJqVjBCiTU05NIbaJIbNThY5RBUI8GI50xhC2QsuG+OjyW1nxBLclFx3GYiR
kNFa63YCNb7IsmiBYzNuzTS30YSIlKA+BVLSumV2Ez/kFIDtPR7AOYBYtwpDuCgEhffbF6ByV+5l
vc/hZyYJRFHwpg561W45yYVbLMyKkINMlVl/S79op+tO0RpaYGyNurx2sgo3XB6BGUjM6U9eqG76
oR6VvLYYH256knzjPg+6Wj8Z7TtloByeTXiIIz3/IVqrRqZ4Hhkc7mv30sGtpxqz1YybXx2qdcsm
oZTqfr82Bpt6LcOdPvXcX6G/3hidHKAeIgz4qxW2ifwqKJuvTXO/hf53jEDKXWTJ4lBcP0Q9JEss
aBRmNerw/izkeMKncz6CtKE4Oy9CCYwLwTgcp7iBrZ1p7e5Y467YdTGO91EDoysJRnzDd9uCD47f
U9Wzuvh926d/JAZ/B2RgwRj6K/CEp4L7szafY64KRXJc0XTScGOjVYXTXaou5eweYlNRC+TnqsJH
8iS/RWNbGXciRneBy/LjJ0jxSNgT7Wa26u4Wa9mNE/YuKyw1aYQApeY9xmxvefUshlbVPxmR8oc6
+xLIDVji7/+sVwB7puJwEX2/Z/bGtWNod2cWlSyGMAbX0bdwbdkI+otu/ofW3QOtZSdiwdbamue6
3OYdAYq7ifhc5OeErpb891UMJV6Wr2deBjdm/aL34apBN6qK4g8bpLfigGhDtrWZx537DE3Tmg94
Ufrtbkk5Z/pfPtYkTnv5tUgE8cnG7SIXENW5UdtBTE7W40e7UybDuXDIsem4b3w12pw+9fB8G/qL
A+Mc3wKsZnBbSNWliKPJqDj/B+6xwWvpCcCnZ3l4I5SpmWgXCLbEelLORoUI6o8TlmpCNIkBTVuO
oWFF9riXyQu/cyrPbiB4axS/hyt6mCL2k2+HUdtXWul/6fq674kg2kCUzJP6Dx2gG05HiLKxIUCP
tvHTUbljUJg3/JKE3p6Nc9eoX0dszNH3F+Np6Daf30cF0hvhf1DC/bH5F/rjBzsN0aGrAKni2wSp
S8wMnTrMzRIMQQTuGa2KPPxhZYzzo2TsKfxN4oVt0uB9m8RKB7eEXpS+a1B3aG9s3DviSBM/GF34
h20gTJDPLTEcMZw9i0FL0qi3wpujO6y9WJh5qQWRVFu1nZuSTDtRFO7+yrqlPetFpR1BFy+3uoln
ZIn2U15hZm2XppsHAJlBm7WfgWMncIa8gMZGxrYsGCEwm2Fm1ahhX36DAuUEvNWz0vd+zgtK644Q
eaqzh7YTJAh0Q5D4xUDBAKjSrVUNkUK8qNSBQURxbkOrutAyoB/qbWvKEDRuKdkA78uxMuls/BY7
Jtpc1/PsMaKhGG7KvYiqfC2fljQ3YHyKk/u/Ryd8YPc/VHJ8difwb63ignEas3aFr0EqtUrHt/Lk
2/Alx1RjWYNDR8G2vgGFSaadgX3FfMSZigpZ2HBvT7WAznrwIdHU5DLPhGOAfROs6oSlqOi+IHaZ
08Uhe4viQMZgE4+psErfagiso60pDrRUoGEPz8xCOBYCyIXTtd2kMPiQ22sR95ReM86psp1nSI9P
hNOGja84F6GoLwxtEVrvZCYRigHWKF29vZorBsjNFi/PZDhIChAufFSFyMRoPL1xvtfbdJYtH4rt
yEzfl4laUr3ZiUYap7QXR4zWRo+ccZvNpnJTi8C2o0pRjHiW7QsHbK79Xqn0lSDRBjrDB6yVz7nF
A6/OsL0JJ6pf4+Pp5m45tXIp/EPM1Ep2Zihu90ILTfarmHpvDCF09WJxJ9HiI1IEK38JFJ3K+Ew7
NWnBmKQVwpudxT3Xf2Pdagcvbb66xzjC1VEt4BSflXxuW+aSViw2LxLlFYlgLO2L4ohVMoOhYP2a
7eVBUV4oC0kyiFGn823QwnPdhZrV6zH3nM65+CX+fHvARhg+b6z985QwDvqZNW7uDg/xzjQGkGUC
o4AWvov8RCPdC14NYnQG0RvU1FqZe8jV9HXQ1hxKA8EnNeq72efRM+9P4f/dzro2l9hWZhs3PzVa
iAr2ZWNAKa4eWe3Af6xeQ4kMHRRZ5/X1g0euXNICPNkLRN+kYqGXa6riWmK0NF53mR18u/TTFbVP
48FocBaA4hQT08e6W/Gb6nEI7r+yeabMqmf79jXcBpaVswPaqVmtqEDiVzES13ZFI44ZnPoBbfDt
WXQ1bmzX8Rk0alK0KeY/tsE9Wihji3r+uMalxKRL315XAb0KBt8IJR39zvAd+bU26Qh6T2ThPI/d
dsHm4KO8HMDG9WS07sFReK0sNoGJ6kTl4hd17H9NAgi3WPthYs4n5UeY/ERHKA+E2ys2N3Qe2i9C
fHnorUNKSRQLlFhn3cfZrbPlOwitBVHWr3AMS/+YLapeLZc33++4FV+slcxScmlRNlGjHcpWGALY
D72KPAWUcICyzWHBTIwdcqlhkl5Db3EWA+J8+A5Uw+5CKn+0jsxDtY5yhBrBHY71DXjaQVNMQfSl
UNP0dSPbLfCWTthGBdEHyk9keJJ1rTBUlyvxUPOJi2smj1gfKsv7St9XbqckePpEi38erMmv/PeQ
5spRut6Uwc76BIySMO7cl4ysABi9PNMD1XuHhuU9wH7SPY2ZOdPDI6dm3Qpz5P1c9XZJTbBPJLnW
x4a204xiIf9W6jya+7UBwzPliXRRCoGT9V1zOYfaZfYtGE8fCnlLiqI7b2Wy+SeEPakVRpdJgfZn
v6GRENWQgQC8Hg9CXTqkgvjcmwK7is0ecQuSGjtwCgMuB2ZQPkUvS9GHym42dcxmvBTve720N11c
utpB09NZtj/o01lgDyCh4OV0w+5UQRNMvCHX0TA9HMtMnLQmox75C7ezYdH5kq2Yi8PLDikF5lHl
dU2O9oqvJ5pO//yiXvmX8V2L/X7sD7c7eUyyfc/i2jWCY6RprqrktEYn1+L8jvpJJFlBu+BNNjDc
2BurDvQ3a3ZAAaGIBZ5iRg3f4V5wS0cCmWcACf38Wx3XTLwFH0Jr6/AWL2TPHzqeabjDllKWalLO
Rsisqu1Z3nndmGPlvaVsGFEEdOitdxyvsQwxX22RSfTH0PhO/lybg5KXXSCz60cuPzTieWIe0ccU
0RvR+w6pT5n0keXT/yrT6pycHxSS0etc1hMeZyvpXjQtUWuoA/qHPiSA5eWt6szoTbnUaqMvnI/r
DSMbycM0u2wbL5T1WcI6+cXak8OQtd7LwxDCahvytdhkHhTu+2cYjetUNiTFZAKbzuWlVFdbN8Su
6Jix3NL8tF+seldnKf4y2oTc60wcxBDGXo5wtFiokAT/rAR+nKbVfyCkYd2QNMEEX33/HDGNXX3M
XH6mEAOdvol8HBGv9bAQbbtVdZqUf4pDcN0w5aqgt/Clma14zambCTTWtagOl+TqXGgzT/EFcbcB
PAnYNBY7cBCkso9p3FhtVxNdpiY0Nw5KYd3KFFHId7d4OvCyTBYVJG4GMMUbVSQpeStLuMigrdYM
Aot6Z1rfuzVI6DT6Q4DSud6uYZ8C43UINkOrpjYLJsqAgySQSwAeOhAJKWto9xrJu9YQ0/RI74dv
wZZxqU/5KD+fZVb0ar/t1WsSxPPLumlidI5giPk4G8/pRwJrmKPWbOWueY8GFPIWSdq8nbZu7/Zp
2kE4JbesvlPefCIfQh/iPbcvOV1UcF7CfdxBPtbVW362JvRMjcWtbuqWOLtLe23q5KE0Y6wfZMG4
R1riK8Gg15C3vgTxDvgOaeG5Yi2si+bUNS7O3O2OjgfOmT8Jsu60ry1oLE9nA0sHqwFSwuZ3ZC9J
0FtjUqfffj6lYd8yYAOb9wPhEoZGSu0ifiQsMlDyq0CDvlJnEjJhngB4FARn18QEnytz+697ACtB
Hnma6DEXl5Jif54jItoaTg4fE8kXY/hYlxPhm/9la19HpchvA63JeGo3r5LQTmzxI6eGO1XP8fui
G19r8rby9tR4IUk0OOGU9H5LgGECmmJFkpl+TOWpBBiqN+kLYi9nHlrGnQpXapI4yUzo1LBNoQcB
LO3PVAia+2F6e/OaaEXhaoPB4rw89Evix5St51YJSjJJGcOLVq1Br/Ner2L9EuRyQRVK8IQy1R0Z
ZOE/DYPY+tgP0OG21sZyIPTnAUlQbBvCX8P/TQE2Rfeqwn+pGf5hN/ZWLcrI9hSZFV1pukgYRvs5
dFE3WUMYrX7Fihw91KXG8xbzSlQ0USbC6eucj2qyZi7nQ9WulNgqFa4nRVhcr+2zgYPzaR9DAAIX
JjH0wZyJrlVrxodBlM1kgvc/ycbGINVZWCb6VjWECKPzGLrJ6BfuFetvO8IjMqLEhBkG2YL81dxt
rO6GUCB9qKMH514EltHBesneSGf9OtmvArCeqX5RBcGIqzEf/kJV5RVqOG1ocJP082xrhzIIETLU
tTnYOXnia8q8brjt0nCnzS56zPLJ+udVLXsIAITFo66KN65sB4onTr9C/9sKC3QtQyXgJ4H6gvt8
io8ngdJ+qvzHMGISHAi3bKqWeuRc8qm7EnmoZ7NNsqlCdJ4ChOeefmlPoUKO+NyGbayHtSyPI8hh
+JQo4NIZSEE6DQ59z0d4jWQdOH+UbL0ATsero5H4BWDWFBQyQGCOCLDyldj7r7jyfoB4W2Wr6955
QaSXAMzYsgI9c5Ho8wkYfoJQOVQtxWdJ9AKocW0eRw8Icu80cxmul3Y4gvhXObtk3KaPVLl1Pedx
L13INaef1fUxhG9PGcTfWtK3qAZuh7RIbB8OLtcWv+5qxYEYgV3M0p7GJy0vUmZOTFe3wrzAAdT2
mPBAo3PslWQBNAynVYPpuXdEAYxAkilHsKyDOlXbjwLYSzfd28lV3eVfUwLoppWntbgTATvooSy1
jaX+gyxz+FmX/n+DIr3GLUdRKxcG9uODnLOW4DQx6jDOzFbnWtIDgVKqY6MhyKQ4gnTXnblLP/+d
iIw0XU32Y37JeLsVMoAwlOl26yl9XHeqYjB9XEXcXVhfVStsNsjVawhmJugOYvHaiyX++ge8xP0g
5DQ6tPCVFo3F/7iiuujuVOr32A+VfyfhkG0F9lJ4jb174C7aT+tCZAyU6ZQMTcysddJAgOEUcBkQ
lGA5AERs4nE7AegLhRqpQt7UWHGnlnJXoGr25d9b4AS5WLt4WkNkuiDAM/1CT0CJZIoFycW7L01H
GHGA6OEGm4F9nxYF7lxpK8UDaLlHlbKpQGa2fPjMdLxa2Ln4Kq+cNd/XJ0hlAyzSsemrSIP0pUnt
+2gxZAItXTbv69FKGpwuzw4+EQjAR2JYfyNt/DP9BSFHeAk0bVua9hsNOh8sNHFKThXI1LAmh+Zv
X/kPE5dMFnKa8YlAGZktCpX74LEs2HjE6Q+SSCdNPmw0Epgyb2G5dG8eYSy2sYM/ezRE+HTyRHc3
x6J+J6O1zxsL/IOYpNRB2u0/8LynUhBm7TRyGC9AlERzrqN9iX7SV0v7N0kdwNppxahiQ5OB75Sp
+t0x/rFxV2q3rG+thoI0taM7OsL1TQMHk2tSmZQ/URdrr5MnGvMXRgREc8APE48J3tfRUYbDGQYK
oVFr1sOtvHsvAcXT3OD/0S7u4oLcbQxznQN50u8EImvHbSzIkaYzR20luIGGH/WYRwrXlRdeoBco
fjOq1xa8msw9jQ3Q4gOUze3AA4gE21QsBoxxQATUT9Y2ZAEnXVi3FKGdvN83jm8im7njNBH23Ztv
wf/gSsyHCRgPIHNLowanryMnfhIy1x/WSFheAEvcVlIcmp5gsnoqZZ+7Naqv7/5PwuqfafqKj1Eo
FYY6GsJXlrA1JtUAhKC/6eQUHQfj2/nKNW0K2PTELCmn5fWtRMqzxGqJ58d/WYDXC/zwmPxHnpCk
jINQBTTk77Eqj6HFIls+TZ1FckiroIhbkCf17flEgQnv6fgHIQ3P7Lcozz2+kVMPMMY6nrxP51C6
hjcCMpuXq4xfZXMNuIjhNoh9WnfjZMxaK5XoV9jTUebzMXfTaZwlLDbH0VAHCP5ETjbN9riRdQNj
CF1U/espMXtTc7o6cDoTXKHRc7u//rE0Mj2ZsHT7ucIlsPe5j8ejVSBdUXN1B7f7qhaS6K+gl99G
qinxiDwlh6fimHTY+Ll6BAWB7zcSLnl6l8IB8N+9AooeajrI+qxqTnV7Sd/F0RRi9nP4hbsfP+mI
6+/AiJ1AV1Ah4LdXMsROpRVK1KUoKBsH2DY3vQxdovr786Zl4XqW5yPS0EwPP2LjuASQhor7UUUx
8b1uc7CqbJjx363FhMrs/JUUadhpUWshRvOd+5dgeRDapw/kV1+MEychOgzO+qkZ7PYjny0DNHTU
NBBXiGUGpwJmwHpIHlGsaWS3PItt4bOaIPxg7NwQ7bakcccJzRqeKv7dtTVGny1sIqA7R84S6Hbc
sOz1ARQ1u+//bQkpwC4tTtwJhhK01WLdCLBhnn2yBD4xb1HsMC7PKB/R5EWvChA/PIqLFNhn9sU0
l82d26Jk6ijFiwBDhlaJzacQ1Br46ahBTIY/vuCeJ49jUjNN4Ek57ZXnqDMITB7PcRpIZLffh/Ou
sWMGf1mrB+nZcdh15WAn3NK3rJjZ4tX7YF1TxU1tKZ1GnZx1vl5+LsoaFCz69+sxfGhzZPPLUugL
FryBqSkQCJSxbdZ7t9FFzkGwLzFfT1rdnMl5oPRdnvws7UOI2BmWQTgn0SiMnvJrYslYy8DmOpMy
rL9zL8rrDZrWFsAgsXVnWdvXFVYXrrDw+3ZxdGYJtTUEln4mKniNzCV0my60vZX9I2teI8NnZhhl
G0ggPvgYdg2uiLx3cFqyGMIVU5TWJ5BqqHK9nozhieD8rLm4EsRvHKB9imtPPZNf2T7SHnL4ToP7
drCIn1bQtjsL2Ig1wifperbsoJM7PbSzxiB21URhwRBPcDGBh7B0ExcbgzG7GHS3MupfNTaWwpJM
qTAs8dtXTsIO/1FyBxD8NShct5akTqFgldNFDUquLYqOxz060oWdNB3NQTmd7lFeVZ0ny+ewhQgY
O+7c8MFRr00apvOT5OYewFgNoHrI0KEwHG69c9pWUiwPb8I+tDVg7dZawlj5d8K48xTGu4PIMFLW
phLvXP4POSFRjyWX5pb6x5EPisfJ7gY7K11I+JB8Dqa9j1d1aivCiHnyR+DpnVeIqgbEph5UrUiU
RYpzNV6/usKGIQDRN2M6yOl9hJip7FVIeJDOt4TiZSUJkKGfjQ9d9TEKNxGs8RFkMq9DC8kbm5PF
rrASjUIHtOE30OzYzuynWnHcCasOXvceAWXzPbxyFa6ih7B/2Tz62CtKgY4xc4gAO1ksPPSTldXM
YcbFr8deDoY5jGcs572XNrgDbmqNdPegPzJxUNuHyQkIKx1127SCrWpQcx3IvkRLFDikxYVI2iUD
F65b24eAuuKeXlZ07qFMEd+f5KwdkfTJTmhw3JlTzMgWat4xfRW2GHtqE3a82qFM5eFvInqNh38Z
btGpjsdRKdRYA/ePZRRDDxuGLc8W0jK1UaMii8je5b4bN06tB8tetTtiRESg0eLK4oFBwNvewdsK
I5Qwguvv4m1gYPhthmHsclIkoHdcFwxzyq1Mnm+0qqkiJn/Crz7HHkMEs/ulj9K5t4vS70RknomW
O5r3qH+qnLEun4O6vFgtkkg571TOLaRaZwZtplKBemDD4SAy2NKfyl3ZYVm+gDbsQSuY7zjwsYEh
lFu9WKepxj3SvxcQUgku58e2jR1eQ6xbxRZUvPJnzotydv4dzxGu63NR2JYNqnqW5xbT/DDx0Yu2
Hd06QQkETt3TTiwy6EQkqmn8V2/T7WzqXDEtmgb5P9ate0hykhVAuBXbdbrDH1o/psvNO1DPI1xL
1sLEXVg2UjEegCbqJRKPb2q9fxYRzqIQ4ucIRP5H5d8va9ObXUFRBza7tuCjje+Odf7HIvgBk3HN
npXtztdKRAlQuTeSb3fsMfciTNhqr6e9TceSP9+ht4G9FAcviiIadpyjeU52CawN63MysIClWIIs
qwRux5S80BphF8lvtuuur61MX9FgXoz3Fa1rvSAph13rEoBVOd9THB93yCIuuQGIgb3sO6q4nEdm
NNTQrlckINffI9KnVI48AsR5DycHWHLgj1dv5Zr8JIg+GFT1HUqzglqaK+ItA03pK0FoXgnpaLvv
7HDtk3laooAwdxihsjcQLbmPTc8cNE6+aVXKMMiexiIza+gfjKh9BDM6waz39nRO0s4SgV7sjxo+
BxEeGZNSWQd7h2xJXrAvhM1r3qbbasSk9F4zoidkHnSzL7h3BsxKNTt4R7XwWBJ4bOIwi3Tv1Fj+
/ObQP9D7f3hvqVwo1bpvGpXWulYL6WKZK0O/LuZ6F0SXn/4U8YI7MPXMYiBKuetuVYXODq9nMJHP
zQBJ4DtdjwC8JAlbkYXVYcvj06OikGzEP+/OytHY2+Zun/PHt17fvgGAsxEEFuGJIWPpyzlHG2MA
oM/zNgKQd5IqLmXTqIxc+mHOZJks9hmkxqiHJyexSiEgcEBjoTvxvx31Bcj65u2jtaVJCd1lEZoN
WeFejeodP4OM7NbulI3O6S7sWTR1AxEGP6AtXRegvYI6bYV29sySlM/xWKXi+EjmSHKPo2zhtAng
MzvbgNzVK8IHoIBjgPE3b/5UI6QYktoE2Udydtywpbktr8gW/wNGCwmOpbahkDzv1D7akvEG2pdE
U/YTZ6bcLik73H7kL3hRleQfodU0tByGHkmeOLo0ZjtDbDxwhUTdOFkEkoGGKgk3NnzpalvIe/Zx
o9ajQXqUpEdwEylUm++eGEUv0BomGMo2C2bpFp2kf/MOm0gb8PUFTyZ4lf+8lMFNXSLA9nU9oBTU
7kcztZqNgsKORyI7HnPFriviEsv5/8BU2bgLmeVXtLQYH15E9DOIuphAUDObVM37nRUty5Xm8DgF
mdSGUXLdCYLEgb2QWP2zceDBs+yXUuyrqj68qq4ZjKBeQ2IeV4DBT/DvdrLRpRVr27NFoXi6KmfY
hzEAOUqWrh0bgH3A/W6GwU/ma8kf97J80bzC3n5OFgyiiRVu59q96T3bSNs/cfKz6HGNV95ONrBF
gRWAIr7IAe7iys0TYl5b4ueji58YLkmsaZ1HSlJI1dsDY3NCq/cU/WQH+2SRYCOdCe6cS/WjMHrv
F+YZQb8fxHTkvCpxIBb5eVnC7JnwmT8Vab3RVhfYQ1xoT9ckhIlBLRUkU5O081+gfB1e2jnKjGxZ
UPk9ScaovLW0tVRxIwprrus9K6C8pd2jmeER5v7YlS7watgaZJvu9x+eftVeJeLok5suHPnR8NhR
O9PW2QbD6NWMCBl3G85GeoHLnhVzRO2OAGHOTUzLOV+ME75BLspcMkcuSLsS5gKofQIeQdx2Pi0J
x+uKfc3IRKb4uJoCkB2n3AMt81ASiSg6zFLWEWPY3yyjU9+B4xO0dMkVxv6VYCPA69d3X3qP7jqM
+9R7ChxvHyuIwH92IJ9n/oDzSzVSlNNTUDheAgvJ22+fw3yMa3eM5EBr3SJw7bOJVvrwkIvxS2lk
N4jOHTef6AsgbTSCYmKWa9TZ6fMHkUocr37rpGjSbJ5xQmMDrE/QjUVPtP+EteQ2UYBGTV+xeL/M
B3R3J2pVxVmU3HnDi6Bbk9JIGmWqvbMCYFKmk/H9OwGnNRvn6ZAjRCBTo7X0MNIVbmu+oIrP0MdR
X5knX2YhNlTfHEEkLK+H+rwnJX2I9V6CUf3TWby8uw1uUWi/GGZtoMX5CObOi7mStnx/tUKGrLBq
A6S314b8PSBdzu0M/5C2B2/+W9apFloIJjhFJ5nW4ZDhXj5+JNpqxifsXW33RtnMpngnCWUJVU8a
+VNBnXzbPOSD2LA/kDVql6wZr8gfM5vSkiPFm9/dTClECsmEpJVyI1rno/OXgPvhbIga5K94qRfe
3Ru6TlZ/AyWUMfRe9dMy35O0IPox153lIeaV8wnjN7VO0GUXFe8tGyo7uLF/3+moq+bNV+yxKGv4
maMtWZMGmi7uPVLhzRsB6TqBy5VunYuVX3BNLN0dss9zxUAlYiWdPFYWNTtvAjYgDbvg937YDrE6
upnjg7mGZjqOXLnhxreeiTFfcOeDbyt6UxOnyYlnAsuWnG9zVNYALhNVMWcrlkYE9TEmtjd9rElS
1Ups01P5cD3Z71Xr/KHD5Hqmm0Wro3mdvw/tD5rOPQzAn3v+VLs9TGc1oTnktFGXTYwFQdAo5HrH
5oJZqeGtjNpZ/eu5uVNWc1/vFzNYgMeb7zLrVy77YS11tClMXSJYiQnim0qQg4eBABS+Gp5JjERv
+0f7FVV4pYeXZHhFv9sIyjRNaggwho6kgRdROhpKJ10LAiALUBQ2EqcJjgX0BizROQzvDXdVawqD
1c+9zutqa0Foc5s1M7qaSR/EKBFChTQGJYa3i2h+It76fbavXZB7oeECjz7pkBdUwKP2CtmLJnfB
eUERoJt4sxu9mZNotZXvZbfso74cuiUQRpihD+K8Rt1faWwC7adD6qZ43JI9ggb9WMk3SIXOAyl5
MnSPIVNy+gG6ZZtQbO6bm7YeNBMq9BhoZqH5hyDzlgLO7sS95LMeWbnUBXxrvmzn2g2TUZmItoVA
8K3mr+RngiVgntSYStzZZYMBKZn2/lC8AQunUcpI5lk/GV6NzL0zOn88p7GTjBMOKLhwLWWNeW/7
hdcnblf1p9D5Rh+G+xmpfJdRbFsfcOv3dr4UwEgD1QuVJNlqFCK8pgBHEBFjSPkNfRAlC+IqIjb0
DZP+8U0YSyl8qH0XBI0S+Vi8KDGhjth36Z2H0lagA2Olwd1nTCYks8JXXD5fSpCdds/KhSUtnDcq
IvkLhClGDBTcE/pfELk81xaz1XZR+zKFS/hRdkfFaeLDe9qXNXalqaV/YlWFzR4PiqH2bIvOOpsV
qJSLlrcrDt2QS+oa6wuH7zkSB7jAo3ReeVNO4990ITSyiTaAYl2eFIXafCrASDtKKYnv2uT1kac9
SL2AaVzmmTF9ObZQ1+8M45QGGcfIFjnzcijzmM0NZ2GM6647FoELN2RbnLN3m+9/9d5af8V7lnQV
CvsnmhtORqh+HhSHzyeP0pp+DqrTCwvBS5XeGWIrp0kOmECXSSa5vwskDj8MSLIlQQkT2dgDRI1d
hxovprztDavuL815tHFHXN+2nur+f21JRc305wf6OuZdAh9u34S1plHL/dz6v/kwe5xW38TAhLm+
+u1Jklm2+CE7bsP4cPsQU7wCGJ8ETbsWaD05C5/4En9c1TeFoZYT7R+/pd9QLK4V2o92Llo02brx
whVOgIqdoA75n8vqfYhg4BEFSAZumrYcOAQLxYKZgXI7HYVyR/GHxN6XGGSOkygDajF5oTLmhoNR
iXPYq8B7kOePP5g0Ov+66573GRuRtcgFCxfzVyuOcYfas6/RBBdizaWEOcT0MwyVN3bDCjtBqjX6
hpp3FF7AJQKzhW+gjnBWIIK2Vj61tGq/ICW4lc8qKH11Z38ueSvw2ITBUJSXabVDjlSYDEyGJ0LB
JN2Ia0X0Z+8llfA2HM/9lo5FLHCadjiw668rwK79pccmUywK7BMfZM5or8vEOYuzEf1BOmm+mzsV
8oFH8ojPiOwCPrXB4roXRXPxukabcf8fOobuxV3RZiHC+Rl1WYCN+r3EuG5LWTjBTycP+SccLdSW
a21+xvN9uIGKzt17dWGg16HY+zFH/siKmGjCMdEAeZ2M/qSeu5ELgjfSxC9rQc2Qyag+mTGcp89z
aHlkLftgOMYvv2CK57/K1+fnaFJ6vP/PX5IczhbCnwg3uPYMXR+FaWYaTe/yG8HpDwzCIkMcYn59
2i4o9NRYuNUiCciSTK7mcu0lnTeZ4UPCfeu30BwJ8uiqiokIAgDIS1BUC5zAUE/9luANzd99Xx5t
lbOptsf90jZcKgHtrXck7wnM5Kf6241sN29x2DHDukiASV4YDueAQdVzPDhsy+maF9bqmUpytBlO
IRlWkBnSGvToOWEdKRqMWrcRzxW3pG4zFZBQFErqzRYttpO8oIwuzqaVQSkVUVkFlEkJZoMcyqLW
UF02PtnrVvrGguQbIp6S5S42Fs0M2usBjlcNEfWjIilfF8oxx3yPxLIpDju2X8iokig+sjSK0bAO
nAD1Pe2ZFh4oK2q1eEBT08LsF+kdH2nF5O9OqMjC6GaRTH25ywAa7fGxvSYXfhXGEfVx91R7wtES
kw/gMQ9tWiVWJdiwvY0ZYNBqm0Z5PKcXz/uDEU2ARqWhOG4Y6asD+aHqNc2Yw7psQoViy7mBf0oq
blPZc8gxGYSQeLPTjiorawdRkNECI6G6aFoDcv8qDpJkZEqzv1w2azDfAS7mDG+WZKS2PssTxg3p
mphX2DLypjHXPDPVzcIKWJJSuDDtREfM3pmN7K0aqG//6WWx5Zsz9v22luHTL8ghLybV7s3fjHej
Js5kcbv7dP8KO8OGVwCAfb64SdZc/ty5ATtuk3ehYgq5piqXzNdrLwT8puU1D+UlE0gOR0xoDBLQ
XBL8oVIc8LQIk+sobd6tLWoxF+GT9S10W7VGcRgNUFdSsMRddgQQ7r7XNz54BEbEqkEw9EWLXxq0
vePNf9S33djn4lshMffY251HXwDJkdoJxY3uDJFcbzyU6Kj9wSoKn9e8fxaHu5PAXJPuCseX9MH6
buvC1T0tdOJ6IRszQT5B4JtMDXlOrqcco9S9rNDocNVO4zoFFCZ3N6LUPCRcMob7uWW8MYcKCTlM
cSSuU1ZhQe44y/IXghS4RlIewtVpujmZnjKIRi86+apLtpQ881sLKAajKwETOXHL9ouFuCQ0QYkW
Ylo16Mcksny5wpdXwzOmXnF7PuphSbeG7Y5Us6S2DUW7f3RRtzKe9/Xfqlh6E3PdWZyfC/vq4zgb
x15RdKrujCnz7KfSvTOYEI6Q1oLiiWilFzc7GqL/B5n37n9twv7M6uysm2VdZA//z3wRp42GJI2V
jlYH7F8/v0LZaUnCqBwumQBlYkejICbC7zP9uub+XvWwdiyHT6Hixm4vxWSPVKLRqPgodsGqXLTt
Izj9xc3OBK++FxLu6yzSeL42bNoCfoZmk0CQz3NWyyxBKE8jRhYVrFjHj8HMdroXp59fu3JR08r4
856nyrMVqShjKR28JQwzPz63o3iZw9Egb/wOTU7X1U0XcQW6KwNJJDqg6uCMpHYRMeagMO7UpJCb
csSx2U5IPiGi6Y9WHusiE3v2w+145ZD2KBQ3a+RP0ZGtc03BIL+T4lOte99Q5WTPGc/Ucz4dn7zn
e8IqdiI6KXEs+27CWyzpOHUs9oQqsXEyvTbwTg4+2jRoC75hXcj6kME9HyEpIY2nV/3crrx37fDR
ijqUolNiZUwie+ENyCDVRrK9zB2jV73j/fL3449n2tfHbPcf0p1BLlJwAUvTQPTWNgTqoP2XyCqG
AjVpJwnMJZ8cBSKMz7QuhFIOduA6o8cQjvgjmTLN9lh5uqYFjxp8nYYvfj4F61BxXTQx/DFAbFck
6uHIYAxQcy6QOHvttU9xeB14GnmR/kOr/INel9imV4A8DKd3vUxU8EuykpggxUgjQOFuZ1TqdHKr
AJ4bvLuzkSst/3hdF4O9qZvse02XazcoQS2ZobsU9Y+bjdr3UYn+AVyOUN/YDO2omphmjd1kOuRA
AsbE8hH+2VZ3T1FRUuBYc1RtvRGTzlgFjCkaKTucJB7SVHJmNdMvlY4d4DzFM4u8xjqn93fSgvQU
W7LZNsND47ArJW3v6rOtWZvw9IGiIahEHX2Go2xn0CNDCwA0xA9rr7woMQYNVxbmSUjFfHVFm6zh
emffndLwtIh9EU4GWpDNsMrBawZDQ9xyQSrBHbpWi5/9xNYM86kY5GosjrtQF4rQWYzSIO6T/8WE
JZqfIcnqCzGO/2sGpFIE6QiIcQenZGRmf5IfPB+aIIIQvoF8NqDz9KECHeBGvaK4vzP6rr5iF6/N
CFeE7SzCyx5RKv82pYAREJoq0Y+OCUTwLLCzGnR+FPFYFePUHMggkqd3/FhsEiJJx6RMJ3Tn6eX0
oBSthlHtN60a/Ui2YRVpCKg7TSDA9ZgLyr/0bHG+lgfqV6/uRecBJ3UkucaEE0G402Kk5rnINSSH
8QbEeT/IgalF6ErIjig+uFhdB9ILGuJtKwpVRhNbnw/nYB4Krz9Xt1MbyXkt9WGjUOp7RMS/v08o
Bs2FV4CUrcGH39k3hBuoZsO3temIE+w39MwL/mpnaECIWz6vj9RqVwKa21xMVB5GvT8pcgf3HUNz
+7FxB4x+8JioGlp9ogwMhZVFfEcVT7jBwT/QOxmegr+Dl+L0jUsXmQDYbMQeCTaA/1qTRPuH8VBQ
Cyk6y5MTzGCdGFmK/9Jn506nHu0Y8rCZhLijWNjtIFClwMHv5G2wHb58w0hZsiOzysAht23B78KK
tU7sJz8cCoE53bmzrY+uORfryUFWZO+jRExtARzXoTwPEGrnVNdR7zAXP4oz9pSgMKcry/j9Tyb1
eDx2G3+bYtEratee5B1Ckh+fl1t1SofC4tdyNZkjQUmwem/EhbuYXxBXWZTGi+DAMYCK7Cz/zTRl
FLHIn8ZgSG9sOz34/DQpXiWzYjapvJu4s95fWn6i/Fx3VNn63pZmGVchdhESa3aTisnUyP6pVmRV
ugkKvUtI5YqAHXkH3vzV/9FfOBMBFiPK1JV2n+0z8WrGZz+l5XQA/ZVmSPDraQfsIM4o9rSGvr1I
NSfL2jTSoaVoZpjfcUR85xSya9VYifdpDyNCaeYu4bdU1hypXOwNCB51XCoiKkIAkN6hPpEFtPlh
RJKbtfl0bgsUMFa9hKPY8I+X6BnGhPQA/TBKwfDT0FmiXyGXncGNm27nLgUHCgbO6p5/Hs1fjCJb
lU7fmL+M5nPiwZ9tVRwoS7dXnx5k/rZImqAGCin36Gp8fLz7AGNLBVIgux+iKUYO7Vp+ixJXOFrJ
6hZJjtrWhCQ2umnWiKGQAIyTxY47UzPixsFO4YsONNBiGLmvJGbvDBZeQGiUCjKxTn3u/5+G5Zgq
FCNrttH+8Zk0hedvQVPw+RMrBF+/xVrLoJj+JYL+PX1h4mvziRYLUb0hRGHtnQ6qK1rovr39aeRj
YlshWrmdkn6diQdz37gpGyeDDgmOvVuVQ7WrcUPi8n5ZdZ9mELjsLc8FYjNBUDGR45tYKnt5mVhc
S8c27u4L04XvPcK5oirKxxbhN+Zw2UmDz0pYglNe/bBhSWE1r1Ynihq6zfOpzba7h00gdvYqaBpK
Eo7OJsPlWvWoqbK7nkBI14VJ4FmngUCF+msGXB6kQe1iO+ZXPOImHt5XTrNy4B00qzgm0ADOSIoW
yk938cQsfjerxBOwKc/ngP0QxNn/p7aSCbs/Y6tbz4EAMwn/Zfgw4ZR2uwR8dPF8gCiygB5h4aqk
RA6D/x2xYkQ1W9Yrb6gLhrzt4MXz7zPH9hq8mCvKgxtre2cKW0PdC3bYQqUwZRoOOkmXLPD6bZpL
m+up/H983zfF37iCWf0a7fsn1ipcq9ql5PFoyfko/kSE4WRmIRtmYh8qlKMvBgiq4/bt5iNvGbjB
oNjUNAQRutr34na3NhdDAYMLM6U8g0EmCQxmG2Uw93OmY/noEgVrKU2NPPGlxURE0z9pk5AAmD9c
LnrFsD6HZnA5qGoJzXJHBye4LgiLTpTDfYGNquRLgqo6b/HMAyKFtGTlOG37ra/XJXxxJX40Tozw
+g+xwDlvUZNyUzLPL0nAw1Uva2I9Dw5mTH/JdcWFdPAJ3mp+2kxA+kRkQU26OeJHoHXVNfDK0SbW
QydUprTpob2IogXxgCnvMkWfJ6Ww5EvmJjUye/irIZYndjojbMmOv+2GCdlw7+o0J/kQN5K+QVHw
V82GoWXDtWUM3ct6aXebrwTa2S6ACHkuXSxWc1+8tCmN1Toy2jXYsKiWHwqdzjbmhHNYNX2AtHIy
HuMGNZFa6GiUrGe3K+GbKZSq1/pUs50bfmCoZgEIaXJuQfjBuqHP3kTE3q0/p+/QJgzgci8smzyB
jjSKOfKSx8LBufn/c9fHCYxIDyu4j1smKrS/BtrH+ArTuIDsI+fKysRy+Yri0h5f7PX7PkpwbckG
zMV9F3hKub9GYCAtACtsX+dMFx6aI15mchVlV6OmGd9iAvTd8qEE2YmwY8WMGzMy1dk6qa9YclW2
R37EgsTTAJfFJc8OuqnLlfpz1mkIp/6sVJiupir/LmL0xhvgX7ZvhbkR5blKmU6IrnRIiSTqND6g
51bV+hK9IzbfIxaD5WkOG54T9vF2KMg5BKjQYc2wFvbMAcjDAB/lo19StVZ7qeUF5x12+iCZAXzg
zZP0aWRQzaqC8Km1F32vgruAeTGzuzQDpD/6w833sD2AVuHHZeOS8tIv7NK3NzDCVnIAMXWqZWu0
hDtNAK6veVkJ/I3eS09nvlKDysAzFabZ75BqE/f2/PpsnDv0KeoGlO6fyem+2NTnW2+j/ZVLf52M
WQMAVJb6UVa1a+be2GLZ+jVohY27PwZSmF9TSGSOcAK5MVGZauORxUkgT8ckJaXos/eLJEzUx30o
PO8i23wMN5/FJVDLwvl5AtiInH8iOK6MJOU9TAzI4a8xZeWx5ycJSpTRqhff0lOo0steJsen/agG
wtGEvwQBkEOeQOHT+pmJIII2c26NaRJpNKYoTK6AOQUHF5k7PbW92Wq4onZECtFXCm88Y4wIzw7X
vSudv7DLeDbgmHHGp6aoNkD3maf6Kp/7SWNUkFe//r1jQ8BIw1KzBxTSH1jVlF4TxZ4WFFNQXWSV
hhvaAE3SSH4Pfc2srHZs/+Z5/cE6FApfj/Y94mMk+y2EmjdkCIaQ9CzuE4FP3TaLnTW0ZFSHmION
QRTC2XbWSFoQJ2C5cfWyQX0rJoxtvoaEPq5DSvjbCaNaXXuZpwmCjJ24SQtsCTm/1e/LtqVNhV72
6dl9x0T0gMpXA6wKjYHYQAbVebcLJ3cSS+R5zHeuVD7fHFxjSU7HJzHO06MRB6v2fB0MN7jpl2De
+H/VNQX31NfaekrVmv9VC0fD3MQTsfItL2ywJ4O32IBD+19w66uCUjg7Mq5VU3dMj+kGKCDJxLKe
RuMGMkrI3WcWnKiieRIU5NCKa5RdHpbD1zDtcboN+d5aR55Y7Y6Zg9nS6HScEou+zgrX1cRdqiJo
7hG+bvTiAsxnQ92Md/9vepbT7DHJUCF13ONI58Ntg/kYJVJu64iH0FEJJ491IeaCRmbL2La2p/uN
5hX5UgWJmwGIVz7fKq2hgxEYZYwDmLab1oKNjjsHtAKvxiwGtwhDpyNGaXXAD6YNVWvD5DGT86Gw
JkfigulSxmuNNELqdmNT80XPhlq9puKFh4fVInvflR/Jdx/wkMNLnIilsMnj5nkQsgXQcWqRYRZu
yOIxaTano2yLlmCpCcAqQtfF0OpSBSK+yyppHDLTmh/W0x7e21ILqVRMTBVTk+jT0VHp3PCfLZh4
TWnhcbdE61A06MoztT+WERVAKpYfsKJL6qPYMk6LOyLFD8o2RuaZwLfLTnu5+oCYYlxsrrgWMHZD
mhmU41JCXBvpPObPw+4fZgFra97ex2RTA4G58LthszyC7ELQEeDU8MEhCulCSOOUTJQ1KNImsl/s
zDN4NRyGvYkftTpuGlxi31n5RMLqiyylM0I4MYFAfHXVTpkQDTHExEtXfKrLBxgR4bsgvd0So7pd
m8Y97NlIMr/ANq73QJT0JkV98A/v1SlT2eElDyNuheQlNSFMI/xoBIFsg67u8maNUpIKiepFYJYI
Zjqw4fPPGtF2KIHmTrobOHWAfSo2uLfB8qdBNamFx2+8XnJX23AHQfX76Ai1FmHYT8j2gXvXGtwZ
Dfi4GkwrOlQB8TZ78Ac3JTVfHWM/6ePz+7tKu5Ikg/IsT8McvZFVQXZenNWMspXd/1SeZ7cutg1i
Xmo6fZCy75IIILNt8RFYWY3kD6JIPZXDdcPJwtVFQejA+nBha+G3SKL5ZK+q8Yb/NeQxRuKjBn8+
Dj2vIFxCoja+Fz1s9uOSlK4eNhC8Qt0CR1EjE0jmmnVPl4BK7eBEblRl2qNA8sPgf+3PSjL9QAPs
1Wz9GEaZH85+Xs5gR/5y91wWN2pyg+ASko12JG9NixjNXvFWafXV44kmPvUB/Cf+3Ga5M0EKEdq8
uZhqNg+0Dvnpfduo3fd4ckyeeN1d1qCdy860k8WGgB3MOAjcHBXx5l/YPM1zgdqHW+kQeB0W0phQ
o2+tArRr732y92H9MVj93BG+jiexdTZsaSCGW8yEFnG8JX5/Fc4AyWofutdyhHrZdlZaSqkQw/wO
ygywHIC6IglUTL7jvigyGPCTDVywFCvhYHpGEKkLHdXfmtJVMKNdhk1APQESA2nrWPcUEuT1jLUf
ULrpHNKBt1TBg+8h/yFp9TUOi9Ft4XgxmoPFcw/ZxGXtVV3E5VxhSI3fWwmTZeZ8m+aVIFrhvkyK
tKY0HPkjF0LuSSB10PLlxbdcdzZyzky4pdibRxGqQFYzQblI5zC8WVQPIdS170GNkSyuEOUA2WcK
IvqnLd3+u7M5ZTgDPjm1JeLuRYMVWdNB4ZZU9CiJeUqj6zmKZeEJJqK/m1NKyGAJmXDXTD1NycGv
+enQ+Kp5MSfLUg7LLyR6tLLxVw+BGSdTU74wbKPa6zHgz/3QimLjCHrCOJn7GTIfCwylBeOg7UCq
qPJzhaScP+nZsn5+iaCYztZxZU9UzPta9GGh3Jfgqc4hWCt+SGxwxXrN7lwRf3dAO7e6EbVIbZY1
MAFttRLGlSgrolIKPr8O1o+AI6m28Zkb7m70TvwLRHJMaamxni+HWU3MboOPZS5yV5hveMUleDZY
gofW8vAJ2YtqWMefFqyfOgNyulZ0KwF+/y4sJoeCeewRx3hXiYdFzwdH48p52avRnVbMWtBy/Hwq
Ecq3H10DUWthiqzJrt4EYAynZdkenUVIAdekPaC8pjz7cN9RKCnwFXcNrC5t3rDkzQBl29VCYpIm
ti/GVpGxqwczJG1NrI3OlHsEb5lIpRj4lHr4ui9Z33ugX/dGtY5jPFfRS3rgPtSGOpU9+4JGT/9n
J+ZspShJFvK+hjZCzxSBLhNMLMjPi8uw8mIfxR7kWb1ywP99VyrMzxf+agvlpkYtHAvD048smH1+
zuhKOkkrAbuwuDfWrsPRM/jeUnYlgeoOhwQ6y5ub4VpPfP2+1ROaB5jNDgB5OIIo4A8dGtbCKX6K
qB0msrN0RONg8RTAf0Je+/Mrk1nFeMhkXsDNJ8RxXcqskTsNZqH4zHLpzYoT08IQQCJbtN5M8vQo
Yo3jaEoJNdRAalrAv06109wH88i/EiHkuPp06NoV/d2J0EOlQsDGhBaCrxzvOFAeMR53C2kY9lZC
CBEvPR58yGQay22ds7k8BJus8B4UA5URQgsIEFqGbvknoTlwnCZs0GDgIOKxILYluJtrnoary6dR
FbmrxTr63EWbzpZP7rljaVfTY/fVZQ1E8ywg8LEvWXntaCXuD7IeJJfYZQ5wGpIfv91ywsGlfOAa
b3ckyfT1SHOm49RfOOFcAkUIc7fjNLs/bnIIlkf9DTVA+sA6uaarEMjmFggYL0VjcljCiO00Kqec
0kD/+gHcY2c5P43wxSk7eVUrSPO/WWEjQm4uKpp0K9iYJsR+62i0l7YdYa9MgGRCVL3E7cBbI0uw
xy301lOSHduqSFTRa+/mfM8yggt8ctcDmZ5iBo6O8+yO+Pa4fTMISTHa+J9h+RDTr8ojeqA8IuaR
9vl2kbRJ4n57Jm5+k9Rejs1jckIJAPSVQTFnnP3E6k9pHBRCGD/Rd6liMi0QKLc0vzPiWj2DiUhQ
nATgDXtueTnLv6NqyeRfZ/5xv8Yk1boWZOuWZsqzb7u8R2UuV1cLGUIpHiAzfb5DCg+NtL88VBbe
w5qT+HUz3QliQP57Dv026vdg9s5cQJMDG5xmcLAnFX+VDZf2j+VX/sQyUH6/vJ7DxdvhObQ3K8j/
Tu5xv8o0qZ4gCZkQYahaZMb9IYQl26VH7BeRTu3RcXsOBAOO1803G5TeNkxiZ8uL9HPvCpI3dVuN
OZChL3fDe+L2fpDpwfMy/D7hMRuV8nNlT8hr/60Nu9fWZIeZ2BhM2lfKQCs7AN0XLUcmcUPqhg+a
KqHDQhLXiO3UwLemDpcalwfjLX7l4V1EO6CHtBJIE1r3g1dtn72YEebK4L8/lMDpaoY7ufDoanFW
lvU/OgKWKvYKMFgy2yH7cGsehcuHtGUIbnZnN9t6xFcdtSsLoGUC7cSB7E03CWe9mDeyh164SwB4
KlaDlotLLseQyjdFW64OwBqdxcBVap/ogrPZaZc32ZmWUuWf/y3AlIYAriYaplOifPAwebe7uyXj
olN1pH2j02Y4D1DZ8ZISEjTQJ2p/nwSb2IeY8Bymmiw4tiKvRPOSzPhjnGlNWBng05BS/pPYHN1e
aW1NPjZNYdQbWdb9woFhJDclaw8qNM5nD0YMZyuRckG61F3sAcNDqDv7bPMBpyCmrJ/TFscuCmra
BAt158sSWiEgmYaA5nCL9wduUNP6sf9uuxhuNnOiqMkdo4hqVL7NQ57Gg6JOSkolwimjl0fk5AxE
4aguFkVfx5U6Z44dB1LG33UVlqPMfX2Ynl7QG+rm0j3WBRnHQHnoZgZ+5sc7kgwMzTs+hLBEMDfI
2/Q3kFegwMaqO4Y0RMWa81RVeh6GMJA5CRgXgO30dFt4uM++CPMA17XcwaKSi8GruX0quE2sZx75
dnfstuKBfd7OO7Db4+E5SFFIcjajD3O3AE1ZidyrWXr54rWkLJ7JhWeZCK+D/n7G5u2d/dwslzc5
Wqtfyqbi7A6qrRJgAhPORNk3Ss4ryASE/gH2HD2yn0FXj+lFJYMQkSdloCJWHwzhnQIX0E6zLhr6
ieQlaREEJQyO1e2BjHmOuZDJaKv2UX05fmcuq15vZUsSFcPjkmaXl75/HeG5t3S0kJvTIXUMk7mn
pBB6hen/5HBDAWM7vvoPJoWJ0x1XcjMgGDN1cvkyBZG1qKVQOBigDLQl9A3494B0AQj1pHNBpvI6
9aWi1cisAZaa+iMO17Dlr+JE8MKdaXLkvhagN1P2pH9sqByGNdE8JbxAuRKzQULWkp7otM8oZ0qW
lFH37z9e8Og2itD1mreokJYY6qvUUKArJObYUDprWXWhGTlTVpm+Mvub5UEnOYitp7IVxxB9bsRi
wyi206E03tOFdZ4QZqDzY+2uyHZORHTOdVBtTzS8+zGXPAo0TsFiS85+f7GJLisz/E1WkrOc7y2R
ncoQ2/oKjFpO9FbaPLPxSXccXhMO3Kmq7BMgUsBaRtS8vMofzkgYCies0WPrZKWsC4eWsacdV4Fp
XUeAbz7cvuSjI5KJWVxCVvH7vq5P8lnjMbPScOX04z+g7PC6r/ZGlqkYZz+l55QDXbQIpXiUyp2o
/McRXTieHsn/BL2u7vezUc49TW8+rdD2498FA/IzoxoTpw0GXhCMTkT4+d6gLU/PuQ/LVAo73l+S
LNXlKEYIQ4k/M59i+JxN0hch/Oac35sTk2YxmmYvdiEMJpceQFuXTuRR80CXi+yt5vNrV3vLrUqI
eo5iEb477LGWSUF5kGl78+9jA4dSXXfcVJZUfs7/V0wtBADv7yHEIYMP8MersqmOg4GCbY8MqEVs
2mqZLp2X5+ICGLskA76n2HcnOucH4XvyQGzobCc94WAYYwt/6m/VIwYUw3XeGJQem1RgCYJ487C3
ZZ9dtv0ecyua3hwrblVJw//MGdyZVk+SgEYDNeoXvLsh7cZnIG+FfVknBzt0iPxgE4s8fZEFFHKx
Lxq+49CZ7EkC6D4QwtAnCzTuEKqwUpL8TZy5VgYoQITFnSoK2Ohblg2opKK/lyWRpg2IiDhtu1PA
6UWt5bCnw7PW3Tr5UAUwgqDkmbvP9KJmBrMJ9gx3A/3uDfyU+CuMZwMe83jgAKMkezZHTaAkVFd5
pG9QLbu5mh1ri+BslLker8UyOhLMfPIEsjiJe7VonsHFrmuX8efW6A2NSvOkJXX0/d49g7eMAeRN
Ixg79LMAsk0dlfd78/Rfbhr9g4yzgo0x2IaffiK3SWx8QL5M7LW9PxrTnH6UeCYKv3heMLtiPLTN
BK2vvQAnd+mOUzpPmXfvQO/JSqXaB7udlobYbIwrrhuqTmelo2crhpr3R8KpZgIWPOU5u5rTKd7n
g2z2sDQtPb0dpwHxQONmquLyojShXUSI9nQ2px/JxNcishtdKJws70cidJe0sHzMpHBubIDGXrmc
QyTaT4a+W5lYuJwz+nE1TBzaS6SIaNeBa81bGBbANvMzIpWHP8+ivWl8fryzkSrzaOEjCSmeEesk
6FaQ+QPm7cbeyFlTuIB2/8lXabBCJWtogN2LY7BPVFQb2TqEZGWnGirzfA90Ke8PQM5zS8CEWfam
kiDMBTU8b+EE82b1EBp/muEt/WeaTAhqgydVCtm0U//WzkWNlYIodJeAnlzEoLCOdiQI6S1j0GWy
5FltAUjQ8ecY9+hLaYBH3cXT73LC7gA4luxiOD8NxE6WAvOttBbdRSDJaoRfyHuLFRRW/8XJDN+E
o+lNvTGH1E5ZeiGKMhBzzNMy8kE2nRX+M4lDgEEgfoMeFXUY/JC+TKNO5WaSIOzWgMT+vg7OfrIf
HiFTRxWY+ijqHbvBjlD8yueZTGqyDZnHZphgsa8MNZxN4WM0UaTDUFctRb9+4sodUjMalx8NgjtW
7FfMRfn9D1DJbltV9T3GpunNnB48foKKzIvDe8H8vyzY/6j+jflR497ER1WGqCXi1l//Pf1W/QJl
GCN6I4FfPc5YA+bcmvL2Vm32n0Y9RBJAoYBw857ihVsBYRkQBaosnW9jM3xcWXvA1K1AIhGsfMHZ
05khNRYdGBH6wJRCEn6Rz1qvxyOiL9qAAfjYBPFLZrmCI95xLMd6knCs0+ynWReyZjacz9M9wlqL
kR9BfhMTCOk0EwE1dGhv/4ELoXlgWT4wGGrZlkKiZkUpWz0db3E3I7LgTV1GdgRDzpStJM/cmj/u
NQoyXMl7pzNdVsk3hzgvQAKC8hLptSCYqe+pymoViWITk68JR6HST6iF40urwMNyrrZQy0qjPuFU
dMeIGHsPO3+8RmwjrpA1+UtUWPTpF1XKFS/xtIT4eVD2k6NX36Vvv2fo5d07+TNP9BYjcjysyA+y
PglpCoawDFJ4ocUB+qtSmKuMb3G8CVUQ4JiyotZy8/asnBPmB2O9Z3qrwEvotCpCSUZcSsvoP3nC
FuM6PPYTABsl53NLJPfHzNETFpJpmbFe7nCxTQC8FaOj8vkcJ/bobuG8bKf2nuv5MBBcl2XZ2807
SuuINq15cF/BZ9nf0cSmpdVMipI0fbSzoptGxYzi783sZFYa9aX5+Ay6xUWUWFdKCGVNvMbr4SY8
JoRbNp3DteCpjo2Zn9dqOJbtWYYWKbs2hUO6Eyf5VW2Y+DJoMQnDXxzA7YBnoOv+hucp3GynMsMB
TnK771KMrfAQXgjZyLbVARxYjd7LrCe1Io6WkzXN1eavppIDjSHWlAG37xQiEltYSPqNBP6VnVB4
tkY4qWM7RQe5RQa3XEE3OQTllq5Vs+PQ4URYjUh779K1QIQvnGUg9TaXCsnhQM264t0IoFAuKhJZ
K9SuRZZKLaHFyym5T2Ub5/tJFDKqqBSQ7PlwtHK4hX3WefXkc3lyxbwGHE3OyHkIiNNGSSFiRyUQ
I2B1B9+tWIzdhasVf2GRHmsN/s/T6jZu73ISMG99cYNl+crN1LP6HYwNFo6h5dbC1DBWjLsAs6Py
oJxtpl43hjrOwnQwargQ6+I07BLUSNM+ZoZPQ8HEXcrOR0N3Pn8s0EPdzXvgAv2Ng6Bgl0KZ1Q5C
RI01mn6CXNVgJLrEOJCIL/t+UOs7+lnK7D2HczBaHrWD/t12vmsOTGEae/zJtgJW9reCGoxhUlHa
aIySxFDdjU/JKR7Qv3Gr0JTf+HBfWlzyge1GhcFM6W1B+YM/fgKNc3MN/hHHCiY7uq10qiPtHVUb
Xi+odRqd6dJKq1dDEvpotURRLlX/HT2lNAk2o4n6fxvTYK0paFhRLbp7ubrDBljm4nxum2C2wGjF
DDIqQj05RnnWA4+BnpQnEeMj8ETw631sPMxfPFRRWzTfzcT/mNcRHnaoYjOFe3pssMV9ua4d4kJX
yM+Ri171bhrqeUR68fFHhJk7tKot4hS/VEa+T6aRpGZ8O9cH8mf7tLO7+au6bz/inLhQxwAMUZrz
tkcqYj1N9+eh/vGczcZ3tGKRu3euB4yPefewSj6Jj6/9KeaUs+4R+HvOENK9fiqnDY9nGGzr9KJ7
46rPl8pKkiLG7gGm1iONelWvqdPANsumqehrW5DVRJ12apsaY8iUuC58/8jnzoj34AcJe0ihPEQe
nG/2GckDMe63UzPgsjw4rr0smxwm7dw9oCPvfF/j7H06GDhiF21CHPlJmXqFLodMxOeHWZIKK5IJ
txQgz9cE29UY/uGoa1T5NMgT4zEQBVMjqc1XpD2LocsUb2I5w85lWh5wakJ5e0h29TB+8Qdkdcuc
TW1TRsq2aqw00G2Bt6miuQpBWlrBha+rLJCBB5fTb5dyFIM5PpZJyDyW5+jE17Yugv9XX/7CrYq6
eHEmycJ+4ct+UTnffIWSWxHeVFQ8oKi76bY7iukrKmM2fy1aKyBf75np9i2CMrdZbMWIsCC095hx
aZbPsSno1O8qaCJ+EDnyKv5IskyKghuZlbBZRdOzfM/UETDXjRHNsFK2bc3xrQRiWN9AdV1VGx8Q
PuU8RVluZaImEh/pgVrYiZhkOOJri88UyNm6OuNtmEmDYfRW1vLkKgHkt9Qp+iK+swMqDm2fLUII
r2+ANPdMpl2UB0x8yiJGRgbmD5GgLC1i2taGVtyXSKe9nVzHz6GsIe+I9gTwxs3nBSp7VHD/rUkR
YguxFk95WdA4QsUp33yMq2Q3kBDoEceGXUo8UTcEiHYi5s4umzILBxmzSuUPqOz1t7GpGZOxwzWD
9VAJcBEeObcne9Tn7MwFlBeMq4o2mYnIC/rBLwF3eM1MLeCXL789hGCuNBdR2lL5sCnk0ZbZ/Q3e
P8M3XJGcbj20fZmhsfC4DS3j2/d+45ZYTiR6Ciad9ZYsrT8TC8Nra2i6nBZpdSbJloleAUzVyiSO
i8D3eBOyLNrM6rWvZOK95qeI5emk2jUGlxc6RcXyZ4+JAGsO05XoROelrkkKcI5CiiYvjj7s+rfF
fDrTbZuOCzdB0U92GM751mBWalbGrox204NqjylidwCjHTF1O+2+B9qjXIUDod4Oqjvw+yIZXyLQ
+LRSJrfxVcxTQMVkiXrRxmCJz65MTjrBLPT/yby8x3b+Y177Khtw1AC1FFMa3xkZtsudyyE4dCNY
cmE/NxmTL1YNvkeZN8ztsAPzzqgLLEEDsEfXA9ADO4Bz+0b4irHE4u1hz8H/LtP8Oh4kpgWyh0Lx
sm6tgpYDbx/UhWXtXHCCsamLgugA2+bHiINxI/gIPW+fsEakiihSqpBHjkqF3xy/zhR4PX7KPRba
wo8F1Kwuu4MdtH7lfi21bSv5fiOHsPJpDtuln9YI7I241NRvucPZnJT4agDX76ucANILh1zojJnd
2rQkK/k5nQ4chh29iYgvPeK2Pv96yaug/U2mNrXycrxV79seWA4gIsXI7TkKD+rdQ+pqnZI/d73m
UH8o1qCYyDGt/MG0V/3WYpE4l+ikmPleFc5H3iyG3LpQR8S8ri+diSkCZ3JML4A/Ll9NgsdZP1l4
O0hwjwo43WUAWL5uWxt++bN0FWX65nP2du9iBtFdWjpBDCJnOBRm/5WlLCy3VQGdn3X1FnKOtRvh
o7OB+i0CvuHNnhLn/iJeIE9yYJkfKeE6oyMkt1MyBH5mt/Y6LAAe8lsRZs1vtnS5Pq/v4KB33gjo
8CKQFku9TqdkhHj6WJxkHEPoiZAujH1EwZnQbkln3VVtBFTUqpBWqfsPiNnmQcaiH7E8Nf8ne3xK
wLuTcw6wVTXsz+pUjTrAfIMpQ9covS5TbRHdPk3omDTnA7B+m3fNDNBdArzp5/o0UkAToRBDYEwr
MuQEp//16sdWWlGXwTbYTDbBgPuSdsl5n9HKY7T6xn+JUJoEIgkc43DqE3yfbaxZOqSy1RuO9JAY
wX5UJU+yrkTkcemKOz8aTPa6UN3ANBcSdsidg4E2aKWCeH9xQUWN301jdLNzV+pCYIduEwsZv9V+
KLZ/jJqLonLyV83JTLl6K6Zh/VT6Sh/hJ1VqU4Vzbf+zLw1AxNBpVB/syKIKsW5cGEMnwNYFQxLv
qgvCL1IWnq3rdKS9XkBZzvIwnP6xLYzM1m463YlUJChEhU+fi1VIT2DlVNY0LymKky0aeRWRTBnZ
S4h2rO2GGCMytS2uPbHXHTRIEIskhsgZ/m49vKDnkV+m0QgEPpmS2KL3rsgZg+JSTLrvKy6IxDCX
4U8qSRrKv0xjpKlrtlX2SsiCv6qPbuRIlOdgC5H9uh5s1JRRrHa5c/uH9kBRjA++T34+qvd+CM8Z
hUGAaL3T4nQYOnp9Wplgu7O9OfH1TQSGPIGxVZV4u+aXNbwBtTSRXwUNsI9/dcXN9avmPeMBFSOA
YFO7t3V2/DI5kjM1xKC5ilynFTboZ4lY2Kkg2O/cVZ0hqveBZh3dA0ZXxTFem5Qa/4x9U3Jw5irD
tc+onMqJ8+9woi1PomX6yyRmVqRXX7HjWnQ9X/9CrLpzCKSpWGLdNqJmGfaorBHOZr71j3K1ivUf
/mLue2AMZaEeeCWXgSLKOx8hEzzEVl2JqWKedsSRGRRTcfxLK8Lt8SgSMeMOTKHCiE7lIeHaijhM
slI8yTQGFAixH3TAnJ1K2cqj1hUzEXTtSehuBeDcS5INVtrY8fVyLsfwH/h/o04Zb4cW99FqVZkS
89M/rBmZ9EvseA3Lv6TyZVp0j6wQAaF9/WwiWiz98YbYnb1mGsjeTxLgFr74ZloiJwEDUpCASq4e
4COEsh4OLCKtHmqndR41SXb07o9yIwGGTrxuVYq/xXTsoge+Tpyc1sYVwlXNr6cMiWUTBPxUy/hy
HKTTuo1vp/y7vIVeB2Dper/ktA6W4BynRuS6lR0pryf2BH83TjIGQuA/gGGdjZ5S0p6a0M+dwElO
YTNcAYANCLBKqpGZegiHETaJHxpURgx53IBRH0yu5cforBNHpbLQcG//tLspYgdwmc9bnUIBbKj5
UE3C6EFEkxKoTUmoglZvSONM8SSJ58LE26VTAHGFd+LtDLasHiqQAxvVowIyLoGAtPvlwCmG5I9m
C7EgRIrZlqm40Pt3x5UFqu4BSWmm75WJp2y1tFD1l2urn/G6EloC1ZrIi/oNqGFIHb6uK153mo25
rIelfGpj2dpmaO/VzXxzo/bC13ayvEWPTzeqg5xf+q5wZCUX77nxskTwRe+GX98TmdosRXzYr/zn
6HPp1bLNnrVKVLG9vLbxrpxintlF5Yaqx7PGWDVKU7F04tPpwlMAhwxT4pX6k2DPI3z3k7nmKXLR
oGyz7jeM/+S5Eexk6pZKZd/DSnVR6zhkEy8JDQXNk4Iwfob5vPSYywQ0uUQqtlxVruaC2VHtyMKN
hXJx7K31d/76kVrGwE4f1CienVUgEGtJxHZr7cv/vd1dbuZV6FjNkSidoli4OinnQYT4KuEKE5zP
1GsPHHx72QZ9f0X/oIbjK4NxPsKFj/Mxmzavo1kemQifAkiinu4JpOgSgop0tnfoROZU5HJT46ft
RLrvZBgf/rN1eElSWqjB5x6X81fCpG2FmtQh4f71CBJOyn55pu1MnujBzaEWRjR8PvlEOr5SfhNw
UPdgIaegx8BIyPBdoJqjjgb5b8SYEnqxxzIdJvOqLiuAtdctks34oLOUo9BekooMEaTNgh0wTJFg
7AyT+ybdIgYcFRSJOWO8CG8pkFVkWW5fYltkGemmNJCjjlWwUjpVOo2fOvhZ4lLwvzxxJ3Pv+f+w
+0Ag766pBlnLTg3SBDqxBzHQ6n4D79ktsFTjiwylMS5HQmhlr2nkD8hzZM+B9ITghbq0rQIArY4T
AAr2QYAfgDG82u8ak9Beo5ohUcQMT2/wHp7ihp4QSkAKCEkYtSbzMv2mGTdXP0JR9bNRytKy5tKL
DJAQGEdXBvB/Tz/bsnPZ9chbrCpuskXaf5nK6/VCHdldnwVatWAH83HUVEoE55gSPycK5TJ352Gc
LYq5HLWC5wXLONXOR/pATnw0bBtEcEWXOMl2UKgJxAdpgOygcLFC29QXSHM3qEdVZvcy2/HbvTxg
+XtB9UWsyTV3HfyL9TlFMGynaIvac5QASQOE/IHX7M1MdJ/HAjlqtl4wCzLcllxWjY1iP+uwJD0W
3UNRMegoSFKKRqNec0biLVok/ZQnM3eFyNCW6/SsKIBuHGLrcIXhwKQpSJeACko1OOKpSajl1W7h
+XedBUzd67EEqr4ZnC4qQa/hPu/n4O4lRcVACXxR+7AcWfbsRsvUyzg0hwyxEkewYCXjcJ7mupNY
bcUL+mmunZ8ZGEiQ9NTAttyKmRF9zooVAUZYJ+iOoYYTIaRqhXevzBV7fNS7gqr9ewlpwKX2sFbp
+tJYiebRvh8gwo4Ox0Z5cGLIHc01lCinmK6V7TDSDE3zK/RbiTTjlcl3qak8ZyYaDlyXQYJP07cB
g3if65N30fNo+0oGW7fHQHItRnpV6GR/PlLRuILf3/wRlbzQryPD47auXjXWk4cX25IqsPDGierg
DaC6Put9HTQnksbtS+3k0OaKa0YsOGXVpgLv9G/wpdu8oCIKx3yovqOR+hyMx9nt9F1ur0SUoHXl
n9NJH7LWjJpszkkc7O4uvdhwyR4ty4naDkZlzFXG/7htRe8SAeKHBzCS71Tw/9/EN3MPtBTj3kIJ
GJLcw8lrL+7+NaFNgUiR4OdV5/9PlBRTE+Eq8SHU9F9D2fTvr5+tW89gvx2lnPvGZCmZfQ7qq2EP
FsSbR7scgRC85bG20Ef35IyAO0KiXHK/tbU7d/WgYGP4zUkm5JJM5rY6maDQyIGIea75W/WhhG0T
MdCH+5qpEy2i2Om1CX0aKTTUlJNsgwbzBBKmkkqwdBfwZLx97hXBg5t8Wuys93MJiW3EpEUj7aCc
pEwT61N+ozTFhfgWtshYOUA97Xn+ybny5waD2NUoK0gQVO+psGkoKYnVQ5ZfFdQUMn3gOaPQzNaU
1flLSPDZ7yrLTgKpUgDEfGCE5icjn6xr26OB0mvBsspmkEtAqJSMV0US2lIct/vFrdZvKObUNy8S
iw7m55xyQPhAvlGQrbBqO/JJ29ZC7E/2RYqFeTq7SEJxcFrXWQqGqn87Fo+Nxbm2LsEzNbXKWEoB
Ykw9T+lvf0C5IYqC+npIhozoj9VJscvUTOqKAG5QTqbDEzHT/icD8Xxhe1nHQi9MIFhLduBi5EOH
FMoOEKKM9Q2t51ofj4rF1uz+1WvMw+ISkPmqg6HEoKkdY55pXurgvzdZH+0ULZwphIHBcrIwr2Ba
1RDUOw/8mgw+blGEyZ0EsBE89lB0YAaf42ul/LZZjDFjrKPnn2ClLZNZ6MjZIMRb2op1/L83jMfa
6EDm9HOFy3CxEr0z1BuGN+SWpvBrz3+IroScjp+HRBrKA9mL+R6hCdqkTz4CYm5d6UScChtKiiIK
7+6VWUtv2Bua+imwXkkFSUTiD7NV+yfGPUwvKNuL+3xxxXDUdg7TGi3Fj3CHAZTzHR3Y4j6Z0ZD2
FrvrPrUdQwtP9Iy/NcbMplVm0AILMCxPwLRGIxZ4/G/Byl/e5m9AcnS5II88jre+3JRm5INzez1Q
kAhdRRECAcpIigqcp+AXuMIi6Teufuq7izr7Y6GE8JBe38vF8jONuMPMLGJ44XR5WmcToKRYI8WD
EVWUnb1AwIwFsQEf8jTHGscUou2YyD3MKIU0o3NhtXSrsH40hJ7D//rxtMcYFpey6FgV3kbRJefC
QuspEV7S+rm3NwGZX1JzQnn9UXgn91DghsVLl+tFI5HhFnCN19rRS8/jQYMi5oSBrpjqRUfRABCK
D5dkV6+fAXb4VRgZ+Gwpp+YoGOqjUYeb1ARHQXg7DGTa9iowAFBo5wF23H6TXK3USWHBauhJI0Kf
3r9Z+u9HWhTmhmldjavrJKJYqPfS+2XfQqQbpzI6oRoDoZyoGQewqfCAblpuxtuhrEgdAraGJ48q
VlgBplS06Q+E+JxfU4d+WnO4+CI/khVv6GxNclRMmUHpFlC4glrqLc5NULAEaJHrYVVUanmiwtA3
7Tgjv4vUO41/P5HiRginvokLf9OEYeXD+pot3Gocrd5Zbl7lQjy+Sk10tgDA4POWGFvfCRCBZ+9O
6Lb8Wz1ZnXchgQfW1UXZefdbPaNr+tfQc7EAgsPVjD5QwYSZplWeqiP9ZFgKv6bXglnevrWRp17K
fDt7haPoxfUGhuLU/8ctBzM6ejRS0fD05eyvnyLCiisYR5h6OHSKozFsvPE8cbB19cMqMDB+UJm3
LsJ7FIaS4XEP7C5VbWNp1L2Mw12uCeIPpXFck6ayWeZ8gFdo2me8Z99rlG4OuctayDB5jj3ba3Nn
bO+K2gw3tVIrxSe+ZBaY3UUm6qzRV43Ld9TW6/Mih+twPDZxmIfvKd5QQEjn5s7K6B4RlYPzXy/o
K1kuuvrBe07Ql1tY7Nd3MdgAsgDLYf8Hq93DINCJxprtcWblOogSg0gXkPno6I7YyUjNLPLB2f+q
tj/0alIcRLBVtjlx9SPiJgX4VwYQ9T+gR93CzMePNY4Yoe1hp5eEIyq40vWdgyjYihQEOj10K/4t
8r+QbSNjsvDfpsnButhr9Ujs8J+OgdzNgMLFNgkd+WbgDZvYDzm+9W1BaHikHGEnR310+j7e6eEx
3D8W41Mjdwuw6XwUnffNgQ4UmZJjibowp0eMEyLWin0Ct+ckwveo/vq8JPyzfqz0iBvCgpik93E/
qB4ZqzjOLLmjkKf7CLnPtaqMislcLu614ioJ0UTI0FXm4slXoT1GtTl7PLw+B3ycBPBV07QSEv0T
FFZMiUBjVO5j523kfJrWMqtwscl+Ab+TQpSeZPgNReek5xtWJGXF8mZM+OKytetY4X1fEL7tjDuc
RFmwtTyX8qeT8CC/UAONfaVK4KEOLW/RmjvcDgbmdJMlJiI5rUEiq0yA8NTx8MHks9sQfx03eGr6
sanHL9cDmqLilKJ3xFEQNk2dfNzzWF63pKMwr6c5lQUQzUTevTwFrDceVjW59DItTA1rOETTBXOr
9KBT/5dSokh0wVmrC9sBYSTBft91ItoyjHCZ6a+QxUQ1r3jJbpye0NwIffUIZL39zO3pWoGVoI/x
RnvjYrp5SEe3LVi5j3o4WEND/2fkUjRWr2B51B8hyewAVgiCyAeOAuqUUv8LKplGbDXvb3iCunhs
8FyHuoM7CW1WFwpdG3ZOWGf2ZFZg73pnKyjQ/WFbOFJCuUqmhRoVzWjH2NZjoWTsvv2vEO6SsRZP
bjggqgr/KJFHGIEqoWPr6RmhOy3fMeesnmVml4Tfyx/nCWcA09LE7uXxIys+3QrcE6Q6N/7+cctZ
NAIfxWjiM6/vrGHeyg64T1zuru6xHgrVxZuRtp0tU3za9dtbddmd/PWE09ffhaeypTPpqUw9Y8nx
uOnYWSFl1sG49+/LG1f/w9zjaCDqhtY44iRKaEzi2S9fdanTemFf5POJDNmwTfYtJgWMBGKHYMui
Dqo5oMGkUeQfG1kyBVLiO3pXJ5e2G+AR68LV14HI4hIddhIjZy2CvpaonLOGzSKzM9dNSBFCqEWq
4Hl0bnQiSms9rnd/bWAgjgO76ttFQIMOeDe64y3lze/wXw8SyYYrEGHDNOk4YFzPaNfswcf4ZND7
5swixEOh+Ci+Iq7tN/wFeYzNFyWKzvJb6htLVyoB3LjeSysrh36Wow5CKaHfNXMEFMsRmM6uw8MH
RaSOmS/97j3PmAu/+ecKPiAT/X1IdCbXqX55+OQl1nGi/3YJieHveaUEGS1AUDFHasH27+5IdLur
cCIu3JBOJhEVaHW2Fug2Uu28DmPDpiX8wHzfY5PLPdPNGoqAvtRNt1TlTPBJ8WNR+tqvMGYpc3jF
oGiG5BRMQeIX9vp7XOD5WZraRu0P9zyz6+EpJ2z7uFEr6W6bDru/rQYq6CCZbmc+NAy2TKwsi+im
s4Uy63KZGveFDboAsy2wcd1oqu8xnE8TN9/p/k5f0bxiiSHGKqGTJGl3ZcU1DKGumvW7Zy9Sf6ZR
nGbiXpNVDeTOUO6zxHzYNxTrzF0rFxzYgRMuGsm4KQI2VxdewVj363cNP10q8cN0H/0vXcGG5lH6
GFoRcG3M2TbZTwAoW2rbNUgByKHiy2zyuDk2xP0I974oZ9HYcuugkTJXjFoFiNbE4m4MbsjVxboX
YGRR0m47q1HTUcWMJLRmP3/sZjf793DpY3+CkhD1aXo/oB71iJmioLo4/aNiuV3T9D0v2XFbTlkf
J8H5/aPOEo2hCSBWjMNIepvMzqE5lSWi57RlJz/jPgNF2/Snn/6RquYyJClX05wo/pHk2fw2vUgg
hN24++MXPnaW6zWkt7IT6rcfxEUZ5cremMV4ZTvm5e1YhMYnccVDEmm6U6AsAiQiJjNirqaG2I7M
E5VRyNR26o1ctOL10DqZe0+2wGtKN9UTISqRV6VpvfSXK3U1Ox+076iMdH9Y+yJbalb7VCazbz7C
czEn7/8Ob0wgeoaNuXfATwIfrrT4Pih2TlEViRThT8Py0qJl3S45zePBpMr0nYJxz9WQPx0PvXPD
qdSlo5YoPW6wTIlBsHDOBuAD3IJjKlfjjQe49z2qoUL1rpZ77ACFhUp0z4VDAly3oOatrKgqrX7v
Q3GCdZfzrI5mli8weI4EPG1wT1/lJwHnOn3o7nZrRXGIH09d2U+zqy1SxK9ninD75/Ep4foyxgJh
+BjOLLBKs0FtbVVK8/p5RwZLRnkNEh9jko13Yz+p+HbR4Dv6rNck0qVxvLO+UHpbRy1xmkkYUtBg
SS80yC4ofPj3xJKvXiWlnU+sZIH5R5RJVXpHZIE/wkVTzipvB4K3O3eljJJ74CEAt3FNx7wLrAmy
9CdUXPCb6YK7MZ+Yz0LTrcdHGa5QaZMKLyesyGmXU3SvlCDH5CaUgh9QyUIfeWwI0b2/CnkPYBvq
bL+BytpUldCl04KHFW1HSoG372hFYfHKVtM7v8WONo/cyeOH0E90aUhGrZdYVMtv9EXjXXKQAlm2
Rx4kl1NYmxp5Gk7Z/JHgD9HKR2gVuMnC7jfd2FSQcg9c26CwvipDHMT/pk6wsDnOI+zNZdRdVALJ
u6BiPrKycpnFo7jIuPGGvxGyuXmMUquRk5V+hUkBBsjF9KlvFsIntnOQgkRs2JmPCJiygc8cYd40
Nc5M+xgvOnwKbdq2tK+rhQ7UN84kesi8KXwtGNLgds/8MkacSQ87r6iQqmLs/2c/wvKW/V+mYdMn
meREytdBYmsEUztXR+jX2IhW/G2MndgruJo0/t+lB3kuGPMkL8XNg2aS7xTjpNTAElMBvQbme3+G
4MMFcNezz1f5Xl/tqRhU0Yp5fKGCQ2WD6v9Kl7IeqP90aW58vH0zB/FTa/nMUCoKLtRk07vigymj
8oQAuD7CXt1hqtgJpmb1kmrkCJJvNAhWr2QXe+4spN5RlC2R6pUNiOOjAT/IXJTU/M9haW+tnRt7
eKshE8B5DVu/vh3iax0Ec1HvYmQVlr2bOzG6NRWRl4NwbZfgJ1v1TRtL2rcyPmQsfzD+uECb/qgA
Bs29eJ9/e/yjxQ04iDlGcJS01VpmwLkeePNYBaN7NxelybjSHsFppaOZLtzYTR9bYnEYOOMEIu0C
KT2oNMAbZcVcgQiv94Ma/FpH2l2QkWOsMcJqCRhU4JMezOHXAtzV+xa+1eUg2GdA28Xu9MbhwKo+
H4azbIBcxga68+DtUM//qKuhI/OeH8klI0CmriL9+NrR9KSzVYLjjSuJdRo/PwnElKmQJPMSmzdP
Jx2GhnzS13OQp8ZTSvdQhyvcehZtZe9YAPxvkf+QYnyQwNOJdUx//ycKj28/F3V2qzpTucbckKFB
OfG7+behBkEG3NB2HBVGZsdnkUX9D3XiLGcizmurrtOhDdIpPCxibVgv1NFi64Lc2D13Hv29A5NJ
KTqqLCAJusUNPhkblX9zMdRJlGDB12MdLLgZGawI6V43einsryUJSgx+BUxgKTyLBkuND5jbI8BF
dSUEf4zeoM1ZKzGVmsMnt0x+1JvNX0VY/YOAXfz9QODBO4WPVf4l/slTlTxZGIc0FMgUCXXY6uBe
uGehzfCyFHpmvh+130nnHTdLDZDj4vNYc5j+r+BCMsE4H2PuFZs3KY521ec/pVVm4S0999Awc9Ci
1V0czH6wLeISnov7ZCnPu0Ws4mTFyyzANleVO876TGNWRS/ijciC4mDXTS4JhhRx7EONAou9WidF
nvyYUY1ky7FhSmY6e6jbfkBHr4tkepeBPJRhryBOAj4Z+OIh17IsC7zXrj5U/lfchJDcrYllZWj3
IwvtSvtHWlVer9jwQKkv8icRcUvfzbaV8imuRqnLq6+wS3h1EbQzxpWxJeNyjvvwOI99WuFv4c8n
5lF8NusWODVvrm93naYl2zOXS46CirPClUviflRd9Wu+ZsCr/8QoKLSAbNNr62sR7IDVQ3HhBl4v
rhWqyRW7cSOr62t/X8TpEcr9xjEUfzwgf1FRrsopScDYKUYBe1cWouwtC5rxG9LhoyeWimSngEQi
8hYp5/emE/e1Tl2fhSoD2pGDPPXoDv5QefU8wL8mbGopEeoD7gJueV/xXAnXv7Yunob5SOHapXue
C8Kxvm4qV92vWSot+RTJ7O7aXYQutJY3bACQpcscvziDrSTK1dCOWykZ762yZuaXErMka6mSJ6UC
4KexPldEmnB256CTIv1QEqScRFM/X5l9gZkDowm5+bIS+G5aJEvr3iBcw+Myi3LisjHif4qMASmN
ywoVtp4+3aWOnvAw46YLDNdsEp7JzPlxDGl4CT/DvYGNXGBYfF9ErFW8F8qK+4vszEawbGhvtoHl
2hCFrIw3OYbMv8JINehpMK3UC9itZY8oAALBnZdsGMeBvxUInUy0wfqxdivDf47NxfJb4lDMCfbM
CwO/5AUacDhzuNCVetLrwt/c6m0hRlUnIN9TXH3daBOOR38t1Ig0AXuOVCJXTRi3nUqIXXmd1b2p
G2yLe/o+1ChODZGrOq1Eu3ad8cAnd+eYKLP6uqg1ZN9rsdJC4KEVVoImQiFtT8ZVbV4X4Nzlhc1Y
+s6kTpOsYEuYx/l3L7t53MIfqkQK4lxkiHqzBtBUYtEezH6JcoYVWepeqtZER0kGe/6aNMqTCEX2
tkcUo2Gx3Hcugmczi2q2PGlsk7XaJxzecoWz0Kjta/gDTvBd5tKG2l7EBjsbWqqz5eQ4JiRPD+DH
OcAVAwxS5itjf1QtLEWDYfnHpnVthjzrkDhrk/Gv+r12n1x5NU3Yaq9MWoowAP7bbuZ15FRmke7C
+3aleBj0dfYvGJBSLbFFPSSAP1EmZsLCbwZ33fMHM4keqV/R95+crqLiluW2sQRN9p/NyvkW3/By
mzsBUSsGQNm1J5ZKBxinUjDvZpnttksrZ+12U06Hd3BYr1vmSC1SUic0PDiENXpmj7CFNhjsOwxj
atpnqAgbnqNV/+J+n5bbiP9yEowYGMTml38dCPW6N+jcSJ73gjNxrYSA5NVMqL5UH2ZWi/pLMfo6
C8BmQMJQ8QcdXoYXk3pTV9IO1AsvtbFlcxgKfg/cBM7VESsKCFQFYGvIQJGuaeLMj2xbrC23Qz1W
VDAZmaV5zN7Mdn1PIqQc2XvDR3OYnKonRKCd2b6idj+et+bwSFQiC+E/5BdokXEhNROJf1txzQVR
88409K80hdICTpR5SB8aqghJ8A9yWG/Kf6pEMwGfV5O1qNVfSuGSB2Q5MJsMu06dxfDNNzDTiYwo
Gk+NULOsBgQNPUdMVuiH7NScIXea2X2/d36rONo0xGQQsnn+mecbKSAea7+1zuV2xAkZrYE0IRy5
7UvVjXJ4p/B6HIxNdIuzWsAKnCd1nFLgJI3z3BFqfCPAyAdsW3vOyO4EuapBIfkf+kfs8r5es25b
aZSzjDMo/LbwzP5oXy/UrOngnRJoKkB1/f7y4WVxYdHni4NreoATo5wKGO+mpZwW+lhlHHv7d3Hq
QbOMmJp9Lw0hsueghy15dUdgMHPHdGSKR/3jWrG3Ie0uSMCaAeYQkXCwhoP7vOYijJ/IN8pJOoz8
iu4hcO4+BP7XPkuLAeaT8yT8tVAVos8BoyY+LyTk40KjEhiDFOSD4BOA3htF6DjjmtUFT3KlT8Nm
IgGxipL2g+MHw0MkwXPrKPQ7OIdQe8/PYwm2XZr415CdIgzdrx/kYcea/fK+SrQkek1Ew40D5MpI
y/Q8XIXVnvw/XTip3BsYD01dx2I3FBS6CI4pEf6GxpKuCKhPSLsj9LPXYApBg9W7ESgWPdP7nTm7
wWLk9o/ZeJ+TnUAY1EmPoFU5sQ42wg86VS40ThO7HCXRJH3O6y8+8Lk8KT2SAsmIqE5vlbusjYkf
8Ig4gLn3DbZfSE8xOygpzrMkl8YDpFHuhLeGlIqugPW1A+azd2angIUGLeamC7UljDmDEe9mPiXL
z8By99gQOA7rPXOoAVGJR4E+Btq1PbV3rVQGL+w3P1Oui2lc6UHG5iuaS7tq14w+tobArF86EvMX
5HSMB4B8zU8ahEI+hOO+ApG4D/es0ZXVjAz+3oo8tUJKbpxiPzUpp8lOzsDvjOps9zmUQXhvC/BT
1NbcMzvY8WOR/2Ty22KY/z/V4vhhpZMClz5TR9UXnlXsr9QC42cDhqg47pMEqLTKN2E39GAmPKJm
RL99r1/oIgIIxG0I0MZy55PRFPhMQ2vRoeQ6twNDJGpdcbEq4/nIjExbvEV4pOgbJJ9V9oGSyWXv
IWhpeWtH1rVUFVfBGxHbsWprwKx939q6/ChPQZNxPA/9rJbAGhXTC8Q2Ow6zTbdeRKCr83JeOimO
x8e3iD9VkfT4I7hiEayc4JqDCMAtpiioPsIDGe/0FSRsDRuMnSQISJ8A8cNMMT+3pEvcsdqU0qYX
r5JqwmhNW2UE4OFCpfuhlaSklSv5eBBvzRJ54q0VuArAdhhaVvqpTAfFtsnDbTa0xiXNH0BhzWUc
PldzpB7qxCIP+KYicnAcZELyvNtagwqywzDwLq10tfXRfrv31ine74+KT81OCo7e2EowG9/lBzKv
wRGLqBRiCNYo1GUqgPZvOuHxn0GeJxHE1InXn/jdLTRc4/sImEf87oFBGiqDI5RDdlJNsIQ3paq6
rz3lpzrfTcYwWezlnVpPTkiaj8fchhAW3VdiSskMtgrfUIa9TPrDMq/mW4zgkAHrvow3ZXLcMR+I
N8Nsm/+EXoMCOILSY8lY7BqAlCXNMSIdbFNNWNeRKnnqCW4xDfCU/bwREIib4fd/uV1N143HDhuG
Yh4wvC8c5z2bDwn9W1b+4mo1MeOo/DTGiUZrXHE7Nh4PfqprZtdMA2YUqiumGKn6vJaJUXKSv9NR
lDQf2/EZSypKtuqvCNvZ5pvUrMESC9hg1Efju6A1OHqMuCwEmfEF3psfXqcNT6ZARlll6Uhhjk98
9DydIfr3V+qHGol7AgTxuxXx4p00OvTxOJqkN4wRfLLvonfLvUyo42atdfE5uqJiF3JSXp3zed0r
ROMAM3PzF+8/4DUjZBvvRsKlYHyOlLe7oP4w8ywomz/8zIbnPhzbcNZg+QmwlcTEEeEIS79T1d+s
wa8aLLmoQr0XAKNQucv72CHMwvboaaKYDNFGG+2uxRAzmvkQ5N0tZ+BoObFaN/ZAfGdur7WSI2Ns
Mh/jyEF6QixfMrOMKTMFZsP/dBrOcAwzALvmHoMfIlpwsTG+cRnel/4oSP7Rw4zSIEANTnBfVllg
SkOOkYf/spimWEDTeFFjL1JF2HMterJGPeEBFo6wy4sOjYWHFsjwTTXn6tNipWG384dRED6z+KW7
R0Ex/iK5oglUoiwZJ72iargz1MHZA48DK4A8wTxp9hWJlgOqmSxeu8vo72pGgiV/Y/jWT4AJwRII
vZsycWsQM+vlVQCcrGZ8dor7pzYi02EovKI29WqaBath1/TxXcTFJmvzB6FxmBa8u4r9T0zOB901
DRBUUpS8YNh1ZC/iLlf4/zYPCXjEAgx4ediY5/hNg9hCPDANeky9P2sdF0xYACnUVQ6A0TPSVIGi
xIGe5PIx+IlwJQEyZiWwG5+0LqSqYs5VhwIhbbvDel2HcyFBw0isisQq/oeASSGisGsy9bOUrqMO
VMkRZBO5S5p5J+mYryFoCBpRVbXE3obz1j5uYcwlTO7gSe+dclm5ewsgSQ5WjVi2fKLLx1pXu+F4
Xp8TqWFpJKdy0SH4auDVgWNiqpi9ptS9fIRCPAmtrQPBtbKuJDNUDCrPe+0YgnDCVR/XiMr+7UU/
u6rPDTuu7PBSdlO425fLM6WcfEd4vWkWGvGqd7XhZWWqeRJ5BM+uPpuRyUIs/Pih0hwGIbatIHKr
QQwARIyLo5QUPaKbOa4YPzdZJWj5yeVz+m6OvAAYLHWqloMoPjaz0to7xd/NKR6B6gjQFnnIM2d3
/ThzTvVgufrmlcU/n7Mf0Lrw4i14UswHbMhKSFldQeo5WTTSWO4HX8LBP/wOV1x9VLMGH0X40Nr6
vzXrRIq1iZvpxNKsr3hjNtWOEDAIYTWJ1fkK0mIjwPWSRNZqNoVbNQaJAppZSwjDF0DyytGzWZg+
FnDTCYlTml43hqq6ScXcypmkoWQZETgOIqG0e5MyffyPv5F1gEtp+BvtSyKnLwzNyPaJffrJELcY
rfCZSRfwlc+34C7FBhBjQQxQcjAS0GpBU+0j1PDWt3lziL8ORdKoXA8aQt8krO7PvmQMIR3d8C65
ypLpPAxzYYypMJIvu8jAgSrpi/vHsiHhhMZ1OmfQYKmGmzDRQCUb+V+eGOjFAW+NqRp11HEH+omw
kUDTw2DU60jgVRk73AzNgjKHPKTXTRSkvtcxreehU2i6EF0lY0BFl/IMa6EE8ETgbBooR0obXjjw
Rs0F8wSrE0OreuCDJoq4jRhfdwtsoYprXUjrL3N3MLc2ttmN7p4FVY0aa9/whjkQZKanhTGYxC0G
LdsoyB7BXfHHZ+02m79bNRv47tFng2ifr7/slA1SzVV4xp3bygWBCvwVBCrmBQM1e05L6fCxzNwU
2BQDg60AznUA+etN6n6THcmxJkiM2MkoWKZ5GQP1FrKdWQwuY6jZ+XH61Yr278ClKGkVmTcV/nyi
g+1m9R+rj/a1D3ELv5vqvmhGMG8/2y0iGnI9q9SUieMMo2NC0ouPRWaKsAGY5kkW0R+9iwWwfDiX
+sQfUujw9NoffXOUrVX295rw6Ic39Fr0KkuVceHfX6g1ph2rj2Nxf4oXizEwqiZqLKjUHdKgAphs
+PFTKfiCuf/VwSFP0URfwwzVX2JsqbtU7RHddYHYbRL5xqqjXEyFjQyQSUfDIoedAHaw7aWsfn/o
j/SPJTjmmTPf78S2PThEbvNhwNHD8N5rgFJR2Xfhe4OZ4SEGiwZKOi9i4IHBEN4TNPl+bfG/lbDG
LOO/EP1+M+k1FBxXOcaBS9491M3zLJeKcuYyhVIQc4XtOHZOqlgYzdentcbtVvjWD5IiUvtMh2CQ
723hWJaidujWp2pwPZhiASkipuRy/RCXiiJj+PG+1v2VzgGHXfqghN8N2wb4g8OOpUrrESwpIBFt
ySxCMD6xOp8ewpNrZiCFvgIdzKpZr4EINNtdOYyTPmfqLyrzaLJ36rlT/jlkTpOVhvhy9l9ccQC4
Ij5ZbKh+EhBVjNbzJ5i0E4+VV1GhAhg+9j9+fROziO5IpDzWwUyhRBN0CDBaJIY4LfHy0RO05/IB
bS2DYOXagGLJB37nhZUNCLk3SQZSj1hkMA+EIfjlRCQdlRAESn6sLIN5/iHE1sqaLUazUo16H3el
LbnZoEhfrqk0z/Oc9ixivFbyZrueajBw/baYwoy0G2CIl6koz7BL7PkrL8C55G1vri5YP+81SpGY
AIyoY/iXab7/xNhiz1Sr4mqO9IbwkhTDXXlbfdzQLID3V9STFgdVZAFKFcsdEdaeyGDP8yMXHlf3
BGtg3UIGc4OZfZp1R+IbSl5anKwWaPP1ZO7OzvwXqO+B5ONstFifr3gXp5Xt6Znav7fXyfB0ZCJd
JX3wPOhHCTeMJNBhtfRiUjHcpnEOahKEeyodlRYOr42mskmoQ8JhtJZzLcDrSRN8+gH2TPGOdx3+
zU6W+Q1kva032E8hTSCWCoFnv3CBJo4/9zjda9j0SQoVFQgKUjDrf/UxxPYT/UCM+/vF7ayLY+rg
NZN8YLD2ZMOtbwl0Dj+HinPlvhmo8BED6fsM3ibrUqskYBpOJONTF+lkEIYdWRRPP/22MC1HEUP9
FxZgfdK3RnXFObJcbvhPkSRl5kK0kEmQNGUcg1gt2dvT3ytOU4v44i2H+LVBR6msNSr7glcbdoeU
+gsPI61O6M4sIkvO+/cjx9KVs2Ia5kJlcglsgaWBpXwYPgig/EdlgCZryP9jgx/qgoOuCk1j/L0U
b8j5ez8k32uZGXYAfGxUXF4MLmcsSXhF7f4WQ29kc4mOQFzWjvYTzk4PM4sKud5MAJFzL5fQSOVw
DGU7y1G1tGkVxI7XG8C3ot+1GRa6vpAZy823+vQVd4dyp6McSlsRwI2aTkLlS3VPvRZA+9pp4aHt
vvkLq3Hb5g5rqju/Ool4CUS7TE80RBvlIqB0uxilK36jvVgjCVcHL0udCXmp6u8Hydlmf4HETgJf
6kn1A6PXbHAbqjpth/gEZ6M/4RCfKluhlR7KSWxZuurpyCVKT60gNMZo58lm3lQnhKxPi8/BvQS0
epckdlK+m38Zwfo2xumiuagtH2yHO8+PeopoCev/cKOI5lXGSzX7J+j7QxAR1V7irVlWjudFeTBF
8BCqb/YMZYyxw+EX4mKydswXHANYDuGFaPuOLZnATCT/AFHP+svZMfUscGCGMfEyghocigo3OMSc
lwzGuHszznJQsoDBvAPNlzEyyuJtN6Ux5eIXf3ghEDTQo42N/kMwFOHqAWAsrd+/foKE3zx6oOWs
6LtOTgi5bldzAXAB3DmC2ZSUVlRWQL+BN5hIXFBDRFFpq4Kir23RSMKfH0FzyiOk5Q1X7rMYwUQM
VfFK8UwadtGExUVWYD2w7HSKLt7WAo+p0K/HjpWR6IP3M8HGfqk1yRbaXuZ6mJ5UN/uIJn3XPLtk
tu51B7UVJSXfN50RQyFM9YVSMVl3htrZ7VkiwNspNuw54ZaixDaYrFzUqYeWLQelcFgUxMGPfbuE
NLRJ57X2aZNNKWVR7nP6dIz3TUQ/aFvjC+OETmulYkeB7VjXa7g/cQlqlMpcFswX8zQOt9VbtuiV
oXPT5Z2l7mReQCuLDTufwNRkiHuo9y6CGlA4KFxN2dHBf6Uv2xjNM3yFAoTJJ+inmuf0tO0tXvQl
PoYKlVlKQWBPENzyGpB46Zali4k2/gF9S6DLp04nwxx6zpGiMlpIojQTcz8cDplRvzvShYYS8bzj
1MpS+f8PA4T90AH3S5JmAaguuL114ke0/2OgBSEZW6g/bpNL7e0r0xkMHSIUQ9BOzqWT5LToteeq
dSbzhCo6GjqYf8g+oGrelHdGjDp0Ya0SD+B0kuT2gBjxe4L9aMKuYdyVjUqZZPJ6rVNlmsxGeBw2
XBnXr94b3uqqbxJguecDsvS7rznmE8qYOEmq3h7eGNIxVDu+i9hJI4gN50Wx4U0hXEDxtjOQPPfQ
OcUqI/uicsQorMFw/o2ayQ/3m+FpQck+wwCLWE20IpPoy6zo8GRvLzf8octaVa5iEy2JbTe5UvLT
gPyUBdMaJNyG2/21Z3r8z4Tr5XvDNuld9Rc2fn06mvC8TInwVFqbayzKBVXmx8Sh62IFH+s75yL6
qFaSiNYY1hKOhxxLVgOqhsHLc9kbhQ1PiXe/8p/CVgb99Gt9vRVC47G+AnvBwiRy0GJvnK2Fhi13
i0AwIMHfwUsOL/6/FFdqm3ttUXm0aVF1hBFVcNrtRB1POWYupiKouLuJgFpGF1sCueHnPpt/bciN
g1vD3Hsu5nbBDTB8n/Av6Q/tc2I5d5FrO4LWylQN+MaVud5LGRfr9qyxLts++SoKm9eFBC7aDgaE
f1EChXBxfSq0Ll1skFDEWPctymYOvzsC5DiH5fAtlzR4S8oXlhB579BFu7zM+4C2o9s/KUhWhrqn
apKx24X4C9Ss5i35yjz6CRFwSGsTCJV/vj3K0co69tjVpNXozb8R3hzx8L8zJfUQCz4rP/IkwDK+
RZmr29QFbDF2Vsi9JvmST91/Y0HdUSqMl6vEGECGrf2897CH+kwXthLMVY6cfnRw6mJwIPgXUYI7
CrrkGjUlIDm+kmhKpAUCZ6Xv8Ba7Ymi9avUo6rtZexdfJ9TV21C8MeB5XvpkIDokfxRFW1NbUNmi
/KmSIT/ZSV4DimkO5rZ3O1JVkH5mrWVJIpxWTUT8qTkmnz4+GuE8rrev/q4YQ3pFkcpc3P9VcvZg
iGrxzG3JRNqbCYAvl+dkVgzlvrk1o5kz9q1ilcO0PeH1hQ6iGP9j/uzjNgzXpFnvVNPEIp+UsGCS
632V6oZPGVOQoYYBdanEIj80Tugs5G7qBauFwFz7gQJsbz7TdqljiwxTWv4L+HtcIi0ME07fbPuc
bKlf6GPar2GUx/76330cu1/MXSXy+ysqVzlE2gGrYUJs5qdaAqbC3ohPnovqx17dkbel6tX3rPxZ
mH4fJ+EJUx80tMnhCLYznaiUGoOMRrWO7NjRIe0wdz3m6XA8SMa63o6H2TcAdLflDqWgO7f+8FcG
pN62/8SG55O6jvjncZ5tFIh73tZnyIHU+sXfukwJZqzbJfCHbf6z1oFfcfWatzwZmSqv2BcSw/nZ
a+w4FMyxl3m1QhlqMEUeD3857zE1CoK0EHk3MgFlpxNMh+8quzdedyG1xuTwCzPDwqLnoWjhfhtv
MvoUA6TsJota8PZl93z9+E7unxRYjrzEgQfQI+9hqZIwc/H61tFRT9gjMHFEsJzI2ZWaCj4p14sB
C4PhuC7x4yELD6atqLfsDJI7N+jFuvNe+Fm95B/dAhQDDH+PIrRP1R6WAN7ampTEsX5v+wHfiidq
cLi1wpakQfZHSlEYHFSK0nJ+bufW2lbXR+mmhv60+HmewQxwGvoz496KKA0opz9aIZfYpA3iRJYv
YQMfOuoXWduKvVsRaf2JDonZj/qSXbPR4Hr3OzLgEtLTBHHdQjiVthYGIKnSDKogX1Qp0Cqhent9
aV4ATFxrbI2jmdK/laIVC1V2M72v1ZI+NLAxF6yAWRZRLQ9EvBubKBiRIPQEAAMmM/zdU2+l6hWB
se9FX8EatghILsq0uDpxwXnr1O3zXKqANftmJh7MMJOD2ezZd4aPDtF02ILVSwIT+wFiXmSJA+Eo
fqQgtXCdOOkVanCyDLiiZj5WVsldyiZq79XD+blfpj4y1pHU0PiMBmQzt9LP41zBIaX4A6QqkOpN
CX6dmwuOBksCmulWg/nCIetlRCTCKSaqgJWnWsyM/J4iIMlES5iYGklGU07JkJ4RR1uk/Oo/ZAiK
MKKIgIyzXsNc3IEkmlV1xnQvyFyhVorPTOExSDTdUB0TqAXil0sMtZYNYMZLG0Iw5IndxPEX9Dv0
j2aFCqeoLehIxTFvd3zG50xO4GSrkWF12R1emxUO0jm/nfA3trIhJuTRB9w4dqPItFsYeX4zo71b
pMnfDJg+NQDE9wZujqh1NiqxgcvWuqm4r3HqXrYMi/TVHytElrhrxZFviVTJ4SnSMqoD2PYy5iax
hc16xg7rnFF2G2wLa+98MK60dq6wJuXWgBYCVmXd7xuTz/hVqdRai9qUsSngtT7UGdDJ6yF3Ycol
FaQD5LjCgxA4A85BBLNfICNngbK9qLhFsTn0IoEgfBLYLKi0389ZlDzv/+xOswh616gfEjabHph/
iRJIRbJ42jw2AsvrOMpmqS4ZvGLHlBGe6qBjX2zgvycxD52zQRR5a1e/wIWloqLnuPn100AWLe5t
0DPrzsbtFWR5pO4H3qhj6SuNgJwLVDnwYaRzRBQCbRFhejlQNtVs+AZDqiHQsl3kwn0kWhD9P11g
/+SEM5UtIm5cZX3PmaGGhhhFjnxm+ZkdU5kaKV6YbxLBl73QJh/kQr2jU0gAHWvWNZe0ZECNArmj
BNmh7Iz8AVnOeqnEZsZlm5i/UpINAu9gA6H8ML3YhUrhFrEzep50VtnHSxHF4h/1g4iA3Um0LcnG
9kFsMtoYx/KT+v8v9j1VNad/flpmEBC3tLDg1Jr9Nlmh40GUW+0hqajHXX2d/1xKok7wNcYmb8zC
DCPn2dxs0VYJ2IIO+G+Tb63dJdhEXT3gHWSIyZ30dbFWJshj0JFZkQIjjXBd8GKP83/tOZSfOoPu
yaBZqzdF/fRteVnmfoPCmnbjRbDdPP+M5cOSu5z0bvve7H8TsjDmx6gFhoWpRdpctQrIkYkjpTmT
g8FXcf8JJl3LPIwwZU+O0Wyeqdu1SQU7ATBp1LFDDUCgy+dGeRX1NdZVe5CS2cZ/lZCpeeq2GuHk
pCeK77lKgxHVKnvK8SbQQIG0tkrdqB/B2JtzOEgLfvh5xxmZJTk1Ss0OjDV0ow6xRWDmJgDuenbC
TZRrzo1UVJUvn0SPFYzy/aevD63t6pyZNtCE/h+ZKemPmrvlu2Zd1WaKmqY0oWCTilVUQup+WZla
M4fpnJyiTmBx0NWH2cAtxJNdUi37qqRMSzbuUz6WFRHKsJZehtUV2LS5XO3j+sf3hrLh37YGBpo7
zYtXFVFo0ybTHNBMm1LUNrbqCvCFEwz7Q/Tktdb6R5FhaF+eCXSODVY5GoSHRICJsZTnJOPGsSNb
2j23SP3UduQ6OXgUfK6r1jDf7SRikvRA9yIYWOYFK6dN36WCJU9c82vKBP1vYvBxB7tyjfV34QlM
RxxWi/HIKN3MFgP9i4jkYHUJtaoZfilQowrLHoeXu49R5qCoP795Rsd4HwICHjna2ZAF7i4bJhm4
4NMKbDMVznafScz3M2wIlrQmJ34WOT/n+mfTwYrOEeeJa7MvvrNjjAMqug6i0NQfkiHqf76/3Avp
SWcmRgdaPlzx6YpaDj/HEUKftkywCSnyQs2ECeuJASDeWI4v1ta/HjA5fkUoFOpF2976WC+5qaVM
H0O0vIHh1kOUPtPzRaFzfBmAiKPvhFZA6HO2E/0sjY6a0Yq9cnMRDQ/mWyQ9LDjZBxHZc2U6TLGm
rFT7PO15b1a2Ij3m/5ztn2MWE/TBqSifYRpObD6+z+7VMRXZG95iLZ224OGkrGmwrBVv2unVomPc
ORI44igX7O28RCowcpik3czyuClHm2ImkH3yzrxu31L+N/98KlNB9oR1VNNSMKnG6zxtKMNvZT6R
FLytEJtRWkGUYMYfBLkTEGyOpxYpAsvvJk5JcLQiVMeREKvhjOJ1ZVSmkMqkT/b+0WCAul3M78zg
McX/RZc+QwTmSY5O72S7SpJ0J8yJ4YD1ymGAhhK45Bz45yVOKnrfDOsQh6b5+YMS6UhJcyaqTv/V
YqEIAczjRTX3SHRNTztJj+AVDYRJJdh9ptMYeg1ulPm5Hp5afGwxmtTz6PrASoR46ANoDe4=
`protect end_protected

