

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DIIXDeJza+sKqBrj4qf+gSpQ5HFYwUFgPgXoi9a/661p1fOh7GC1Yxr4QhwzfxxbI2esRkgX+RWV
O70wuqmd6g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tc3vvZL4Z4/k9lIOYWoeVvOilMT9DFpT/2Qg9j3BlHsCcWm3A3qs8Rzy60Chth5nEU3HV6KUki6A
hRQKZNb1v/6vjwTmXalrXjELjcws7f/IYaWgZmjVdYjpJE/aoPqNISqRAxye6F73bRYmttkSLsKA
mpZhym45OoX2lTi2dYU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qQBOLNsTpDaTilOll0jbdzN9+CFe+2YuHpSZBsocYQBx4tFyydxFP4QWzsgkpKMVj+vgHsshU0FN
Wu3IvX6zwtMbic8Oj5a78zbLuCwQAJkzJHVEC33oza9R+KKTeRuoZulmj32txP8npOqkH//3iN6m
rbkJ5ZuVWuWTahdk1WIS1WH0JMwmkoMmZOzkIvY3OwyRzQ7J4JWsuGgUCQP2UiR1wTcS23zdZ4if
K5dX89DOQ5XLDZRfGBzqloRoc2KLKrNKj69bM6afBdivLgfZpIq8pSaRYrb4D4nQ/NQLMqKVQM7g
UtRkTmmMOH9irg/EZkbw+ma+qT3UysisXvIRjQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FnYKQSPwFxsA2Tic0BZESWi6Be2FIedgCX7009o+DpIyXr2I2/Jxc6RNA88ViWghN3LxaxRvHMEk
pR+MRZPIxTWv8WVlO2x5IF03WAJs9GAB6d9KbRe6Gs/fOQS8fMMkXpyEq4+6dsQ1yT9ckah4Cdmr
T2dV46kU3DtfOZwlWxk0OFzQSvWXEIETRCvrsGEf/mlDvxo3c99T8p2n/HDBiBrHIY+98bbLLHvl
mVYYFNZpsys4uRT/TVeQxVr2Ro29URGWoe0peT9xCIdU44Br4X8OPNWGJlsWrkooLMv9dYIUEfQK
VsblVGzcgvRtwlSZRK4G7ikWOKojLVBxgIsuhw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k/CEKtjJXdiEV2H3DdiRA6UDxaoZt303yi4S31RTSRFiDtNKXEWX7hAbczUxcDYrAZq9Pa18y/Iv
ju3h9ViJ/yaF+1n8xAYTxusQZdevYvn8leKkc+XbCxi8/TAYj4SQ2bTf4RMijly6zLqqO004hHo9
AbWF/Tq5CZLrvf24Df0yyJWZTL2km1BM5nTE6v8B0iMxEncPNncJ1g0VKySbcBDCh6+IdZeFDvjk
siaQTjWx1gj+MKrM5hxCdh1gK5aVhC9As2wDY0avEH+1IxuO6QhBjnWFKX5v8fUQvgp5zjSufCpK
Ff3Ce0pbO40TcP98XMg/XiCNI+dX7w8S194wMw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B0pRxV4llSbxSsgbT9dwcuzImsNM7Ywl/K0BGEC/Mw/vBjKJqOpZbs/20GVssjsAwFuJAwsuRvU2
DcscqGBWo/UUVxZ1dW+/mhv8EMGY/gglmOl/jSYwQ7g7m4z3an+lZM1T9/p423pPW8FVM8MYisbM
+tyxyBR/MgTmoxWxnA0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EHRObHCL8AfvkiomPbt7c3iNsMF4eZGxQ33JWJrsuaoV9trVmGm8vEcVPWLNhGAeekB73BJR+LiZ
zi9a08JnSoTsgO+46uuuGrEM1IK8husQ9MqNyNGRTbups69htwaKPx1YLtc1M/60smF/b6euaSYM
JSASlMnD29rew98IbsycQiGsHKlati+Itr7j9mPAlgM09poau5yONp8Qnq4dT11PG2FAMF9RKNCl
UCdKh8nmXtEmrpJH+V95f0ogErBgKxxAVi55Yvtg8bgVdXD9OE1BJxHTIDLs/OWMstM7CzQdhFwf
ujlmDvylJDwTSbP429MwLLobIYUiMwfATB7Cqg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
G4L/F8qNI66KFJu26EdCrtwixyOrCb/Q9wHckvXFrz8P5rHLfmm0oyMRO+5dVvU8xyDrZ4aEzAPe
U1GIvjbyZDTV870Xx+Tu1jFjsuAwsgtY4HMYvTFdKJDiNexHE7shLg2elzG42hW+H+p/9zXnl4WP
9udUHe7aoSaJxFV/hv7WQ4JDBZsg8r1sFSfuGE1HTHDJuU/YUcfXb3gkkSHFHh7Ub96iOcKC6ew6
fnReWw2zCm16dMr4G4xjxGvoXMDKUK+XMGtAhYh8oh8GjeYUwJMUI68ullF+rSItddGheIyanyhV
EwQgBEshWpgE9cIKVLgC3XIVb0Amuiwe6P3aPdLqptz87XgfLN/XgVrsUIOlC2MiaoRzwrOmqJK/
WkZTuoITqHYddaZX7vS8I9MCb4GaYg24Xcm4XuyGpLLvULEvKdikbGO8D9PiKhbEObauMP6lrRWP
6FuiLE6xfgLN9XIGLKpRwvBrI+Ow1M6gmyz8wOVZi2Ye16oxr6ySClr2PtrSxuZUtTgUKm7bRkbR
quPRhBR1hoX8YQ6JO7vinTzDZB5oAhZ69gbt+F7p6jmQ9dvz6NsG7x534V5sxdiiXfWOCg7XiJJ8
607hLIWPZQ7y3LrLcxLRSzxb/JfNXXhugIkYpzj+uLvhCZaH5sNAjGwFUE111kGxZISJHKARbYXe
dkgoRJxZdoqEpswOeL8Q4CIMAi9yoRkqCn6I1VaFrFLjZFPQIFOkTniknvOhfoaboFP8D+lwAwWD
f+2DhC/7F4ApVs30UhcKJJopUjv1+edNoQCgOAPomLKvpR3ssmfhrlj2StscGXo3k29LHiYjCc69
rHu/DwC/Dqu+oXQNZDGSZCiHEcBJj91pIAf6a0kNfSeloQrTXLNtdyDCuncvC5gkQ88OnoCfibz4
bsjJ/h6GN9baPIBpEMdxSLXAuglTAiCf/XNkgd3scf7KYj1NaW1OEI6wd8vb6q/G4oB+hLkPOm6t
SCGF9FzuYn1VIak6hx56+7L96DJKIgP1hSl9HfLsYHfcG/5EIKbcBZBXytv5LJrVgS4nNYQvye4N
RC8VpAtbk66zUmB1ehfzgCiZb6gskDvyBZ+dEvHHdWfAIF8OyPwQkzAn5sgSU3BPEv6rMdsLl6rP
jPNohYhKbyyo/iXqhHbBPoRYnlqbwt0KuHI9rtdZXBVxZZcSMTt2xpxEOE5GJW+xERzAh9TrBzXR
zsj1DJqGj8LfUrZrGJdZw4O3YDTrZ61k0SEwxTAusDEoBYd0cRFtBS2DZVuX2yUeCODzHNP6TOvH
U6VV9BFMVrNdWXiIhd2jf0Y0Dzv8jHmGNVJHv8JCkHijN0NCGkdomvDSgpfE9ATBxjghLtKS87sg
QDjmvl24YKXluk3ZKNU6DDj1YHAR4/6zRg4iJ4TwN6kLk3pMOPy8xnq1DHOeLj/iOu6zf6soTMq4
lb03QPIZe+tYG8uJGSthB78uIGg5wt4WuLucBX0gGQMzopGKqKNaVwSXy3gmPR05wz2gBXa+fseN
MI2j5fHSTA4ZtMpItUVpa/NsHFBj8U/+yt/3SIco8/NTcKKD51GDPdGp822Pm7tgGe4kOXLbnD+b
7UUSC6t8G4sD8wF/M1W+hj2OPYfxlRs4hgR0NOhivMq5d4NACgrTnetT4njulPxCp/GpOSCEi8/u
JeIQoS/bNAyykOcTdiHuJ59NN/HL6Uzgzd6rPM73NnntVpot+pP4EQl5crdqPGG0C2zsk81NfqUv
je4TesacIFSQdvZ0XAQUZIzqODJ3PvC0zk0CwSaUbo63NfZja1C/bqhAAFaCAGYhuYGIRMTku+B2
TXppV0NC4CUNIjRtJGrFWzOU6UXaLKAyo79+GgrKIfYKJxjpwg6MLt9SQhseFIoksSPS4ZsXunar
X1rWpy3pUIcq0i4R+i/zY8ewa73M5BNHc5yFobOHk8PycF1e7r+doKrMM9SDpFS1Km1NhQPe+VNT
Y6EFkZ6/SKgj+vb/aQU1DtZ/sHxc+QHkb3XQt/bsiqsZ+VFErzoFLbUMD8c90laG74JjINpNXmIr
2VUxzUpUO/gn/fwcL2n8Y9eUC4BAdCX1Ic0AyeG0BGY0Co38xvhY/elTa2IC5Jor/SvT8t1tsf2p
3MFuNPh87u8CtZpgHVSFChZ9OoGS6gvp93yUH84XL06XuI4Ui2e4WYfu6AVqvmN8nldp4EozKOrl
g9NfLTycs7HErHRzvrhw3uilidivp4H+JC1FfXB7cdV0+I7/0Ai+c6u6urFWMVmFO0JAgnhGDKwO
5221kUeuA9h8oOpalY1sNuYcv0i1a7DyhKiVlP2VmdFqbU0QBxv+P+cVPojxbWES7+8/wg/jOPOp
jXkhZkDdqtDUN+04peY4OMTwlKtQkcbxlCY69B+24YaXTs7IsaeER1fkCJnjJyfNJpmjDNZidD3H
gqWJDjXAYd/cRmPxICuYzYwfTtF60lAVMYkAMuht+y9SKm5hlFh9PJDD7NM96Bv3tDyd+MKrMwL/
te6/Zet6N90dtoJh5b5pdv8yylVT6+tW3VAipJXj8EBi+B2It41+r4nO2H8LWmHk8bxHsD4rWf7y
q8vQBPMl+P7G09cTBmyczX7UNJZNN27wbA46x68tJ5LCtk8/bWLyyDeXdD577W7KyZG4jDzJRSJa
UZA2l5DJmDvnGo+YcriUzLM5JTwN4nz4dq722Kgk1e51ORhbFD90WvQG3BYjdXQldLp+bIrvip3U
e1VnUjLnjpINq0jP5ldAh6WuXkdGggk2G3ys4KMFuvdDbYfRbIZPn1zuz0d3NksxTNhlu7lExgAh
t9tJwY5bBQ4rC06m9/SPognbEwzKg7PdGkl59Y4eJYxyfMZ9KqL1M84Tfb5WYj9RMO+3yLMtiibA
Puuh5wRfjJJSbMmlKljZQihZb/viVPKhAaaFL+iGtwhSsvC9u6rRIjJzRaG8Fdq0tVdoD/iB0/oC
JfQ1AFkYMnIkF0HKpnzeKttru0zR9PkLEC1Mj27SkVEqLCrcwqSfNBTOwRoLSehZaQb98WImNUtY
9B/ghMZ4Rgc8s/ZX8Hskjb7otEgHUs8IYEuQ5VETxIFVzbSZlSpRh+Sqc+tr9UIWueRkqxJTiUDo
1woMtRfC9/ckkmZ0pcPkejvL56AcFoxb1FHaKaeM9eYMfLftoX4p6/7R+mMBGhwBPaFUTeL6EhZz
72Y+hJpYtTiur2UOYodkmpMiuoPH916MStpdo69yE2NcZnUZsVp1/g+yMlh76cOcSHpOv1r42Xt7
QvQrUloDK7asMR31JGiHwEhMJngg64gAhShj+Rv+NhfukDul0IlpGxm8rZ/DAtbwDa8muFzPKkTU
DAn26Acpj08qp9C4su+L4g/7XkZpfgyy+CkPpUs08ISQ7CRO6hV55PsXKJVDBMHq2ZKEjRYYeCO2
kfOTki3ZQHbAI7kDgV1BQ7nVWC+0zZTm02fKeBFWb14ptClXe3D2DRKsbYXqruC/0gOM0KAWyMSU
uGDl6o0JjoRvFAUAn0agbwUJ8ag0ixuPlCP/6DXOSSbsHPbnL1riPQMANORDiSyxVMAGI2+uIW32
ZPLBU7qLglrXy4Y/89BmrXwXWtzg6E7OLdgaI6RK0vYC6RZBvQfqm7RWz/ZHAJ8Mws6xDlkAcrCe
nYHOS4PCCetuuQwbjt0UsZ+10rAgxUrewTnprbf0lrPZsMRmxUTSAD2CLFrmZXqn1rlH//odiH8v
NWYznvmzUteEM69XVlpcEUKJEaCmxJO0kZVfRpWpAmkZ2BQITi51w1O/NCG/Ji0z88k1PIX+taRs
X5nVgNq2hyXFfa2CkA7F3YJyGngGyLRpvlgQ9DlIhGidj3t3w5tAEzlW+CxeiqIz1cKvHzPodXL4
uLkCsiWLbnzoX6HuZEuNap+m542ghPxxVu9ic7AV7Q2VCidrJ5tjYohmkc+eWiGSS35kbc3IJPFT
xxE63K5iGsjLgYZerxrU6J9TI6CFGhjKhYykTcNWiB51ULEYRVv5Hn43AZjByJ/51kx89r8xIPeJ
4szhEdyAXRK05w6GqOkZ4wKviaVirR+8C5JK6VbvHcwreBpi3gvcdU4v2GvlI6k6f8bO9L0otsS6
bPjaH77E1ns/LT4AZvjU93qZxzWEXAKR3hVywlvNiQvrOvPi6nfQeRRmlBgPB3jlYL9E71L4faNd
L9J0RUqAmlJGg9YHDMKsTzHH2dNEcKikhLxGtgeMKkG1wGKOkcvFsl/M24qTLiWnTHH8KoQ0rNkM
sjen/ZSR3Yl9xyr/FJRc3C0nH01AaSrHeQguhahiqHS5Cte9qJQ+57JtZ5WhKhfop/0khj2lPDKx
o2rMt5Oki0XLXLmUVDYaxxywHElopZ18FMCangcw68mSbGksVr/F/Tx3YwY3oJC15HECSpnfrIIx
u4y4Mg7w23In877xumXKQ1iJGPgg79CHZflfb7m2FU1FzC8PhVSoe0/XzcHougsIgLu1seIxWZfM
5HKW3ePA5TEQBob/7h8ShWj2kSbAVsHZCMpc8ttuZyBJYglwF+9jG/fVs+SU+WUwcjObgPAK5Q1q
XKEp2NxRXnMD6xSiWyl5/kWQO/r6CFWRLfGdFicB/1TCVz0KQZk3KuLHBS4T1PjMB8Io8bN/D/qA
6Rn1BaY/bOBYLZo6os+1XCGejm5YtUl/XKpq0u5toUNO5wOp3L5cwVN5dm2BicYf4IvgHFtU9yQe
lIbY/qxXhj9y0INdT64pWmmXAxB+721fjNjULVcuXbAmypxlAe6L2n5nkrkTM8tmWPitzOMfdjPs
HlFIqQmAu/fcfSO6xHm8HmZxzwrm/lir7OgVLCBblWhtdkZNND+/G1pWoDaLZQTYSfjo3AsJQeHf
xRNB4MeI+wFobz36fPxbw9xE0FAQUTYLXi2n5u4BKZtNJDxlvk5sNOExw2e3bhKuSqxxFQJWhX/8
6Yvzb3f9SrXng0v6OP+O+sPv0I06ZXd5zBXG8qNVaT9xv9FfXEPs7cfuPdgfYLV5jUBc1YhTmP19
RHygFm7kfBQHxw/fdZmDsmX86av+iezOtyORr3QxWEPJ2vy6HlNA7h9PL53y7uAbGWr3JJ+wmWf8
N/yfD50GpN8/ZKuR96E5xzzsEwiJWCtL1v2V474srcHuHFcUN5JI2oQ90/RZ2q9KsRUJEWrizxBB
+okspPNsY4ajXQbOAgarjTnEP/FmoWa0b+qotmtmBu7tEwc7UhHOBGvjTuCQC0wyTld8KrdJbacH
1O/UknTIwtyd6XYtLbOekMz1cvlZdaO5NXVl/uHsWuklkH7bRpohnBHhelyG9aR8iEXH5Brns40/
VynF+rZPz8q+PaDs1HRVYWeuT68sRSA9+EU+Tu7Nc0EWQZuoI5Y/wbAfJfzCpM3kqByZ6cJi2oVs
b33fvHwKGhQqrg22YG0AKkQHNewzmqAMmx69DdNZbDqvV52jOX1PElqizsa8WCCFsIIOVfsNiXQ+
I7swu++FILNVGPeqsUqD1O8N0l3Fw7DaME5CynLYpeNzTrF8PDIV3L8OmFoZGQo5PNSG8liCsAVd
CeWUCwj/DtiXorzm1ce3nIgalJKT3MInOQhjDMLVpNF8obXdmnIeL+3fbfGbusldK3MnNVgBSFbi
PwkiIBY/V58lANLKszF29OoGFqFNFHL/ZVDAzftUM0XlVyBWPrBcOJLlP+VSozJoYQFI4dqZeBPK
XZLIk/msdOeRUCFAr9PFOmmIWuhgeNhJwHYPmQX7NMGF3nOfwbSPynQEKSRZ3VpOHZ61rhEpRFJi
npflkkeUdAUFcw2l4Aaf3/IWC9DtoVgMo5Mcbjpb/z+eUMOMxMNBkDM7UjxSpZuPdkHvncx7STHj
0+J278zZBLBb5Y0I0p4fE7Z0RtPa+Bh3umu8Uw5blP+nLxXVZaYbAaKBLAa5fk2vkmCItrfnqjAt
qfVghgjjWTW46cHxvvCBFz4nNoa6flIbW0dogEnJDU6FZzsxAiRJYK07E+Mk8g8s2xgmMEwLCBb7
gf7eBL863L3LbNCR1E3E+rPxwO4qm5CnORI7n2WqGoG5ZgDv9KKwpM5HDQMweBd3QQq5sZ8y1rnN
o2a+vXwxAIWSbGdAWw1fuBtk+6i8ThxT4v/CXFRzuQjLKgpmeHKTnW1fynBxMCrLu8WHMyBbG1XA
Ol9HTT0uytwn7HQp4U0z0Bgrly+/iYY0l+NoxJOIfj5IJO/QqDp/1n1U9q+dKIB4lmKNA38RiNst
+MfFifV3/uUK1sxysNZnKHOSURPwJJYjDq15t/yg2hfktlzVFWhgsgSMnvYTHBaI1Jw8qWMAt7aA
aDtYlrvVRFPBwsscXsDp1QiykOUmEy7sV2GbZYNrWIB8ckpJstnFXKOB9bgzFF9aLVS2FeXcZKRA
DqDmXBBer3Duq4AxshYAupV4VbQ1g704ckBa9a8O8CQuvgmrFH0oysMCyU5/GB+dF/uLDgg9bevc
LGYINr0+4Sr5mWGpovrMwt4GgSXBSRNCTmVLSA+ev/a9ru4KXIkZwfs14+WFPwHkmMGbIcyCIFOW
nMSUt4S5/J+QXVgMGOo4AD6Gt2AuJzA3UCK8+ns1GXjvqYiCdda56zCu2WyC/mohwgjinvuKsnCX
dmABbugyJGD1vYZRBBz1WfjVIabxqslK5IqNI26DDGVW6g1rDysEOOHjAgujWBVPjERTCz9nvie4
lX8AFgLbdwoIurZhwPkNr12fThmK+iPM6/43N1qs+xzjLpWuxmn3VQYgvc46AowHSOGbLaiBWHsZ
7QhohRK0EouUkV3U0PkZMh28XQ1O3tJ5RFNNz+x57EIUbjeqBN3Q2IxCiIQasvUxN7+cwYVHpZxY
7g+gpQzQhXQxcNzi2M6st/7XYgPcqPtqWKNABM7oCNkTmMmgvl+wW6e2F1T+9Ss18GGGf0aoD1zM
ZczMsodzcGEV3PZo1qXmP7rvl1L3SxWKEkCtZflVYRog+4OeaovRa86pcUO8RWCB7krcChDEOrZk
6O9zZoT8UpEh2ORcivDzgqKpsdaAYbEQ5BgwHcKV1FIoKj5qZBow4BEgbPdtJAuXvzZXT3Nui+wR
Dt9kXI47gxISk61JcO6Ws6jNdsbeNptZSO/OVFn1rtU919TuNVylH428YorGSprb78hPBlsnOi8f
due47PQTTN9tT8OWO40MtdG5xXbpo4q+f21W+in6DNZzgvTj0a7nE/9Z6V+Gzuvf2Rt0h6lqsPKV
i/lyf7e969Qim1ZT+boZ50zr/WxYcjfExUODgZ/8ieWM9+YrKV6rhFDDApbh7u9gGo7agMmt/NKj
B+I5k5ctQPQngpRHCqlTc2Jcrn0izAEKtAQUw+1CUFw/UbjVsOfQ6mpyqCvkEG/JW869IHXxycsM
PaU354jBFUGRsbVhVjYl/yADoK9RB9tybpoNjUOgIE9gAhDxOa8XPle7bAQ6pIqVx5leSinMBvxV
XkwwgHO/IUuTVVS+RWc6iFjim5v3v2VLKBoKbEDMs2OTrYFZNVeG3b1TAJIqx+svLTJ8QBLYJ9+X
ewJSyAjPagOh2Opd1HTiJS8zkdMjBmTR/St71+jaOlwZvvddd1UZv/xKxpQVbpGHNDttGwPjwi8y
yvbjULe2aM7dq9TBM3Zukaks3zghK4qr2UU4IXehp8VCBg4dQbb2UlEq6henkUiC4u3CENBCJrBh
8TWA/p/9o882x3A3fq+w2dBrG7wVzxBaLnonlaqGuYEQ3DIguYZFKF0Dz/zUPUYN3Dkh064LH6T6
wL2NrrUYGvo95qIdc/pEbf7RlzdoDYWYWBASc5aiNl0l44M4BMBchanrMrw8KZMk7XtBa7XT0an0
36TgYl1/epVfFZkrRpIRGYAd/f03Ew2OBJkJpdVl5yP6irzKw/03orV/ZPIN6lZQ6C9zarRmlDRu
1cN+IZpKY2d+a9NENJlyuVxFUmj3h+ID6RUHyOSV1CjJDEi1/xXdm2trfA5piy7CobzN3fxzltoa
mLqSE8ktM0/EMqXIBDnRxGRYZkyZRgB8y28CLzyNPtDYd6+TgLUiSlYs0g6is0NwFk9ISrQXycos
UVEbAhILpGkgVqqqDSUoEl0LA2eky0YqPW/oQphOSY42hsmsCyZJTzlRnhQ4UcjIAzTvEQN4yBrk
3C3orvJFZFC3Hco3jHxJUpuSbfuqjl7vyeLHgja+Uh2+Eyw6j+Xg6g7FobGdkcoc6NkQR0NHJZfZ
9jSbu9aIATd/LmqhIxClGPYyVDt/PTotzmSHLC6UrVNMh69iQ5ty6hWx8dwQFDRs9C8ZtwUzYgUj
kdnzHAh0x6oIYqzLb0IerYVZqLYCJ7fVkP5hiSfwj5rGQCsxOITOJEf1qastYAqXLJl4sOef4H3S
2NpPneTCGrKLwrWMtHstd/VszYN9Xsey7SA58UIu8RsY49h5BWKqo3xdN71Di04PlvR2wRSwVlWz
eeaC0D24W+aicXN4jNxbPbPaXFVqwZzpnQkDKyYQAcIpCUFzFJPk4ypiaxlnz4h1pTu6K31viGnv
dyHK3H2ui7ECGlrphfrPuR17KV2+7PYAU6dotQHZmJ3wEbjA38cBNRr3EGmDrYpomWMW0fPh2JWW
QVd2ZQ2w+TycTHFp+/Rfew5vG/L42+H/tmmkI9LborSIUDtxZXv/SqOiadPvx1tVZ8pfq955OpkE
LQg37Eh4aDa7NGJNvQcWi+LlxV3UZeCZCtFhmV4B3MMaBoIg2JQ0UGax7ZHZm2ZU6VqTWb4K2h8k
Bho8oU7q1/s0l0KpHfTuffl2XJQcND+kjhwrKgEfu6F9k+bmJ4BiM+ZYZrKi3+0B/7qE1DV5+fEk
i0wdfaYls8C2c7fth6JFumZKfnPh1dod9KrgjJfmlr8N/O2V/sZR5xa04FPvA0RBa+0gowT0npVi
lbfJYWYU6eCE0en5lXEAT5ulM0UyIAAR1GqjoNdf6arNpBUsdYMs8h5EhrufPwIgTKPpaisVy6yQ
X+Rs7jOTHU1IpbkSzEcudehQRYkIA/3xczO1e+kYCepuEFyqWEw//jomUq2EwCPFUnWJ4xtnKw+u
PIfCuZfIcJdx305sgGqr6p0tiFXjbWsClz0W71aobJs8GxWCAYd66+2PMI9gPqJCIX9RtMVQ9aCS
iSqCxn80aXtt2gj1YDyVn7eDjwdWh1B3NHHXNgtP0CBPciqFrMRi1nhMpU88qCqNXFPhBBI7S5BY
HL+/YHuwK1qMC+uZ4CYtLlLl/wtQZn6lqf+5sI9Ia3o1/0QLgLgp5b3hW7KtYKvKAeaorcg9lsI7
MhpECh+ESaRZrtOaXbz5OSopL7cnESh/3+Ai8g0rpW/zbeLcM1mFnFXCBhVNDQApub3JxkjnU6Ai
nQBbupZ0iJVeEPu051hehJNLe9mp+eWzaboAy3uYTYbr125gifKonCn8A7ax7V5BkzbX0upJKQJZ
vxmjXSnDZwGK+b0fMnOADYMaDykbwbZKab0jB+jG5zwY/gPltIYg1pi8C+DT4acPwgF+f1h1Jv35
36HCiO6BiRTcF3pfn7e8SoVaQN3QHDJpVOeKfc6Bz7CkdB5KLV/RcKaeg84pabzZy7Ptw4U4Q2Xu
kMDtZQmhB498LvLR02ooOz+7vSFjnzggTuL0oOuLmm7JXXSWUtpJ/I3xNG3nsLGooQARb3JxwhRT
WbPmqoS8uRXdfXjl17VvfULqJsyxNkQpQKbBh6R1s4Rhq8jzLxBkqtvn3Jc07bfjr3mTgJvcwFhK
bhUUJ08x+5M5fUtUQu2lf875JMK6PLUYx9vYMf54rKJzzuEtvBFhZ/uvmSTXT6EA0ivLZvIYhHw3
dtDFlk0Px9zJwZDEj5GyOMkqhLGSBfaRXgDjg2Wna42Y7buGDJcB0fMeSTpLp0zoGcj2y/FwCmHp
oDbaeesiDwDIewIzJnapX+ivXZ9VpDA20nVNMFN6uSYBo7DIUbm8ojeByGq717a6JcSx8fm7jSUk
Kvjluw8pizOJddCk1AGrkKILax6XoJlU4rlAw/kfZHjjzuIICuKHpY6ecpRl2Q0wXidXqh/rwLP8
lF0/3WSFZYf1nhexAe4JFXGexE3vr6NMzxhGocsJ7fnZjGlJRpgEybAd+0nb+Znz8g6SczjTazfB
V5Quov1ZI42jfArHbtXz0wjtyvWiNzKlT9jNoegmzFiS6wXPrDfPyObbSeRCUFCvvBoI4IuJvpE4
DrjBS/qJ7slRliQs5zopKbi/zeb8Nc7Mnl5D81eclzJ7Yhgz9ksPLiRo7bc2mf7RbsGApplMj8tO
HH4aOZVhrz6bFXyEPqCsF+kul64WiAgKLz1t/O/avTBNFElIcHTigVP1U3M5rstB6h/yzgUDC340
1kfQIBx3FPVwyiaspDFjaIsI0z57/Lb3SoI5V4tJJTNjnaqgysDi1xZgd68xs0oMExJmgkt4EO7s
UumwLeEnaIiQ5G+PVYhCsHQmJiT0xQ6qql4qHlS84lbAJTcgGLvHU0aOuW5ZNulv98Xobq2mRssz
lTvxhSwTxI03549ZSvNHQBu0Fe0n+Eq5s8M0BEkRHEDfWR6yJG7sCESUVpTTkqrCymggarg/gkXy
DfeS9sXZe9R7pWSuGlhjuYjf2qDuTZp3BjlfFgGfJoYiFTWUqRqHnlsSbV5syRtxzFqtnpJJfiAw
6kLqaPXawTGqvv0r2NVu9LmdZj98z3BY5K9mZf1/QwOW1h/29mpZhSRcKDn0I6csjy1d6WfNWCE8
xd1pKHgmKLvt8a1/2cFkZ0mcd48EPXsCSTYWKQWaUByrJcchBl8rMqDwzPdsY83ca7P+cMt7sFpf
+GRQD1sOwJkPgo1aRjFpp3aBi2URJdoxJ2N9XhqyDyRsyv2hdWXTv08ltl4okR5pj2RLxbrRpS7F
CJvEomO2Z3xDi/EAOQBNKGH8wp/pVUahpZ29NtO7DaGo4O5DzDb+xapl0eW7UlIM52Qwn2PisHzM
idIKXOM9OHG8h1750Ezh4+tB+h3ZCOYuN3gJqurXHPpdxM+EG7TPijeKVbyODhGRdevcrnOKUp7c
+buRky1glKGN7OgSXW266170/fxGVxw83KMAlCXJxF7QAa05CLK+NvL7x0hjftPtp4BZ5IYnkIt2
+RU8XYuhznLMUdirVwPmS/+V2HoSrK8R1+nWA6r3ID6d/vbsJy/zy9YIdbUPCzxga+DTBM50e/Qi
GtMEI0BsLyDhYe8YUydIMXae0vZrEirr+q7wypY1hDRFi2PBjZMWL5qlDIlb9yYCW0Z8VOea4s+O
y/LDn1crSsbdIRMzhDdggwrmEcBhhU9/Hjl+IMnrCd3t1a56+uZgkqCK1/fyGt+/syM3LUiDqVqA
TKdWzkJ2e0qHMdBz7nLoBLCCnz66svXU8QFgZAtw650mHAuGRGvRoN0TdE7HurmKzQEpwDLcJ9gv
pjfGn4/YQca2ve6YbOs8uMMgdIaOyvdLXB890DtldIJj2maQLwHQaNbctwr45NEINMIJjE5vFO5t
SK0ebxbcnISADD18flYJ85Zwud3xKxaII5LfM3ph/RPQ2B8Ovdb1OrYS/uW74wECfTekWEmsLkDk
01IzyLFDrF8qUeQrOZ/ATdp61E7I1p9UNQ0gCyL7KCuwwNY3BUDRUShq1ythu+G7iTunMOBcrHcg
Zja2RVKQmIBuY3fKZL+yciTfH4ZpFvQScOBsPep5B4q+fxzYUlTuWh+0Kxz/l+yYRG1o8fNoxXQ2
Fy57lpP8pG5AU8Yskvue0QSOCf3o4qnYISKnewQ3kRSOWuwRXfdV7YzhzdD2xVNIf8afmNQ8FIV4
Fyq6a978P4eevvYWaQSmRRlpL6WTTM974IJbTBXcOWtDjzYZtlJiZ+DLzjSJLLRTiF7SHXqsHtmd
ovx6q4nVXZZhD/ymszLfwuSWmBVvNfL41pgkcyz4+fdjYG3BOyh/VGvpXxszhxycqdhyDoaL+qEN
p3wsOtahvQYlpUSR7HYWpTn/XYoUToc5HTcQBRStftgOmOffbRPFD8NXam26rLE72oHk05q0CqrV
bw6hP5AOTYcWAMGbDZriv53HrDEGl8DWKSRa5SBoos7ZPwT8xFsST/M2RiF32v//EHtFIhK04ByU
mSTfpNX3sCbpNotQhM7Vc4tKXggk0Z7KdGD2JtLL4g/svpAccpzuXAhy0QwiN2C2iyGsMMX+7M5j
OYXO1TLlnctVN5KWWFURzjg3wZlA8J8Vw/mH2KwAes7k4VO8yK1Rx5bLgyqeq6CTd9gwxQJZD2JJ
uQbgTytHpyhEkQ7w4UolDtuScKEM38sQ57zruGAyH/ZnsnyiD4t4oVhxHdZpqF7EzWfPTqF5pb2a
nOrdnnEXBk5uLuEw+pbqAJIuchuvnSMWexjlaibBe7ajNasCc6TsZkJkIB6Fr2LIC6pxgc8ghLem
sjPCItW0+gspVvOq4mgCcmMWF556klp+zyiXFfu5K8EdoI+SCu8rr3DnEgO6Ln9UIAlNk78ES40v
XeNN4h/lIDcuElmvHP6Hfe47U7IiVg96Ahuxz+LZ0CDNS4wb+q9JP+dlm0GlcnV0DadPVy0J3qlv
Q8ywfwTWwATG+MrjYeU0TcJA4i5ui11G9rV6aC7+mEqPs0e7XrlhwppKCmQOSryIJNUtVPVl1oqg
APPtUEJpW2ZXu1n1z0IGH7pGvmzjQeJCQKxP7HZ6M6OExgibiRN/iuNEjlyjtCrpMmhtnMtynOgw
Z3HJ+KPliLgM92XgbaVtrMY0Lp3v8okk2vnLlbMOLBNh4FsKcnF7CzRuaY+fsstz9QZf/lSVC//p
y+8QpHb91m/j2U/7L/cEnfvctXwTp+NhUlF0ChxWXs1KQi3d8hYUJ2gXVwHA7axqeoTDkTbzkp6O
oUpNnQOSzbeJ0khr5qblAw0YfOBieETgxvRI5zaBlqIjKbUAAsKqV6P/6ASkSXTn/tPtHzNS0Zpj
bx8GrGYRJIsC9kqVEYdMW4mE9eThx9PuhWaLLkj3tpHOA3+rst7K93E9juKCIiZx/aqVetKiXYMj
kOe814oZxWhSyyjUDaiCZFsNFd09iOuFuANgMnS91JDzGbAZDvEjrcnG6RbE9vPRwmeO2QioTsmy
AA9bDErdlJqTpNh8dIc3I6wulktRG/KYrjF+0BLwc4DSa3i6DXzig0+/xlAbH4EK08r3uaJFImaB
5936Zl6ctreevKdMatQQDJRqkMNnVoUNV4OrKI2xB/KMWF+60xf5tjWn7kbZNfgbcwnwVWPciC5S
cgRByqnkT3lThLXOJTsIW+e0wMz9tfiKVSuFiLMqylvjcYqhegqTQXWH2q6ikffTs9eoTT4ViZXc
dmkXasjO4i4b2Va0dlT55Isbv55HGsj+sI82QLWVfvA8MSeqVLdPtEcRQh3ldkXJEgPHRgAlcAru
3bmg56XXAtOm9V8Y6NgV/hJxPWSzFB4sFuJpTszM9sgWCtDuHyr8ZEMoBX6uwbscz1J3MSbb6CVm
Yj8I9JH+qAo8ZIpQw3Q4KL/pAqzBzLE+hu4R568c205fAutE0shcJoQdnTPrR1RzZlf8I3+P2sgn
V862DPnUG/kdbb0zX3r5+IAijBvMO5RWmLRsAmojFX3hUFdbltqaHS19Od7YVf0pEtE8Yws0ZJO9
tA4/JgLuqV+Mc4QLUVdxvUQbLWm0gfinX/nHANvuB5+cfMYUxWbK8XPX4oFHRdNF4kqziv5y6FMw
ZwAAtsypdgVFQLllD4mru135pq+s69teq7YYlk+OQg4KDkEZb3sBwktGpHxI1U7rxeHLmtNgkhgH
SRImZI8inVZv2ieK4tx9UZ1bY7DJLAQ9YSp7Uvq/Uc7qUBlbxkkalJiIVFz/sCRJkH9PC/sPGaHq
ANE3YtnNvBCu73X6/cAqJ06vG4hi6AWdAOPm5IEHqg57QBU+bpIJUMVORkrQV/oGN0i2KiFN/6jD
WJSCa5ZRTt/gBjBd+gyDSm0sxnJnRgeV/F77NprWLEB8+n1gfuzZAAFJVrIScExMONpvoaShstK2
ffkCvTns2zTilCYg8R4Vi8gfhIy49tRoJ+Mz60yQc8cAXjdT0mUbullDnj4VN79ZCrlzo4dcpMlq
cSWAq7U2CaugF4/Nc2KneeKUiY8VFP7kyLdcaalqerGtQMDY2j/OT3ULUo5LVtUTbwzT8KWWXhdR
DVNvM7a7fqLLfQH420f+ISDSsBCr6tS3WZy/zRxds7qaPdUMN5HiQlbHncv57F57WUD+KegnitSY
6unP8K9+E3XtWcl/U9H+yaW3def6xfDqSMQspXJ2G76Ek2Hv8kEF2Q/W5VzelSXabtiqZkqtnGZZ
32hkszRe7BA5T0t+j/jRYU9NfrLMP2RvjRjgB8Z4kh6z2unjfV/Jwdio+CCKL+tFup4WhsYZdiFG
S1N0kWmgGiQyn5hU1DhEESp1staep31pZN6omN2PACGzTzDPKM2vIsWnXMu2B5wXVvW2ud7Y3UZu
cewPBCx1dsEs+RTijhYNQpTJ6a155MSzwzpJEfD4jlMX3y87DIocs9safR96t+P+mG2M1pVzvMt1
fBlnbkiYECWW+RoRC4C7Bmbjyh979/90XkYjZylU6lH6NL0ges2HAfje0tBgtDrIalPLP+nPnLa2
TwSlX2P6zlb7MdyVVT7cTW4KZ6Ebo7DuhHIxG8CChP2W+6DXJkZaMh6M9r1hbkpZ89+9RgV1Ln/U
pr1sHElKYg4uS1ezKMlawqP3S+y5PZER8XAEr3C01fs9IwceBJqgOKIypKbaFt8ZhtdFnvoVhaSN
5G9EFAb4HSYV/ADgn3HIYNWoitZQeXb3XNoVPOH1AMi/EOH0Oa2wdPEq+jZEI6XQg/8odI3Nhdyl
RgTugQVogQgUxd92D0R5DZ2+PU5xGOrZxfDopon3NN14TFlCSOxqjDhPhsWBIbNbspp3fYlQhy9s
6GNfY02bhAgLclDF+qU+fE8irx123udA5uiOmqI0Izt8NjKXp2bT51wx8ESFKHcUPz9RgBjLZt1r
S+LhTmcPLbT0pUI4acv+RuH1/qPqyS6zlNZZXANkXUd3sdJd8svSWlGYghpz56mSLT3kV79CzYlu
U9wK8J08aPZ1uJ5ZZNiGRRi8H+bzhD2nhdpbIiHqLMOQwfQLG7eNotWlVLzYULhX6gNG6wKwjKwh
THJwbrECTfFivGVrVuyHjCDSPp1xaEQtbwVZ6jfhj/d/89d9r4uVbO+3okuCZwO+eLgXOugTUoRP
/6fDLy+UYkeGfaTpWDb/U7cQG+tt9sssHUzT+P9mg3gdM88TSdUXU7BBNKKMPAw+AM9h41ilMaaO
0Vqp3On9MZcsyMC1P2leagw1epu9WIVaWDLC8dIdCcu/duVy0a7RoUO7iGNkgCwQwIPPDSp3o42c
LA5LfX4j9LoKdqgEOT4sSK92uUAkLtZSxsxI3ve1vs7gQfsVlwQ2orkSvWmpwEqCl5Npp+Zr/eGd
agKxYJ75bg6KyP1dhKPDqfZidlHMET7VQwMP9IAQCJONhOqWp1z8bt5JN7HXhyKlV/+lYoZ1JK0s
4EF8GISn3OZ8QO78ILgr9FvtE8dSRlCjGT/zQMQpgpZTHS9A0qSySSTVpUKadytL2iaIOT5a/Ta9
qLWYkDZ51ya2vaKmOWFEXQjuWFNDlDevNAajRxRUBtOrQZpzNIVSt/Xkq0ghxWnXR+IB7hfmg6fu
8syfK5dj4BfOYEIhzo1kWKbJxkUV3hYSPFQuUdgUcyDUTEGN0lmCu+I7AeKO1EdLJ7VAaFpoJ7cC
nzn+mvduYPrgRIimYuN+gRHOjiB84P8cRzRh3UZiSJUufUyafc6ui0RqznCeiJN3fPFH6j4KD0i0
Xe+5NAxQSoPbloZGVqSOX/cPcLn/WlfkYrg1Go3SLmVrv/XdyihtMFiCqu3C3FDCrAjLlewCUFRo
FkVvot3YXSsY9KdjuoJVHzRQGNkpMaXpPEcFnu6X6NeG1/d9P7HVrsLsFOCpfaMNdrGPPtUdfNqI
TslOJockmsOkiz2SAB5MIAS0DczE9UnhPenYqNPThxSK1JBfn9xB62BnEddzsDb4/5N6OWjITe4g
ZBYuYuHWudkovSLblwXcvj7hL3QmowkQssX/oXFssEWaKVDuRncDafTEfnelcaJGiSa/SbcsGmJr
jr/yN4M8RDwsJ0NKmYrsfmkLMzRApB4C/T64SXZaKcitA/3RrO7Noj7Suq2HiKeNTkj+ZpCP6+nF
xPN68rxylPIwTkuUEPd6PlUNQQuxgxBu/Mb9R6jDLfztGJumUdU3KpP7Y/c70Vf4zg7vnz4efRx+
FAJ1N+bT6lXxcmHxXCfxH+KgsWmXVexz3gkfwel5U/sTyOJb5otJMawJHzbu5FcbCXG/A4apf0zf
BA2y9XvPVPQRuOjSTHqSt9GDe+KJoCCKb8looqayjaYJwGNHyKLlCoqX15+dMNXgszrQk7OgLKJ0
Hd9pwl1jPB7zmP4ei9QHKpTZ+MUUhCNnMkinJx/o69xJdkp2BBjk1OIekYA/b7b5wb++V+jOIqz+
S8FLKWi6G8HM6Dsl15dcbFsJjSlEbtte5lGSEJvUw1KE7gYYT2xRye8bQqdLboyIvokLS8uUpOgL
s8RNLXJMi2ognQqDntH5KsIP5PE4xpMPwLQEu5F0G5+j8kkWl67s4slnxIsxYLDryXdoILBrS6AQ
QZGxqk2N3e3m9D8pAjp8uPFLyz37NBXntYj13yTnd8RNfngFqzUxJL2kjMvAC3164YnedOVvONVO
T7JidwlcMdoNDHfz76v/FVoJdb0HQkjlPCT6U/pZjMtro7ML7tD5g+2A8N4AjJAd61nGDP++QOit
n06TJulDqwCZeDO2SalblA/Ca3pjEtTQxM8Ezf0aU+adVkBacFCu2Ecb48NOcw8abZHs+tC6LJfG
pkoml0xr8cRb2hW+bwLXjVc7ZmB43uZZ6VE3jJqLLofXTMDTcS1UnMJMwtXHCMp4COPkem8KjCa0
raIr72MpHC1Jwu4ObAKstbEZpmb2kxxqAV4w6/IlwY2qKOpQh3lPBpSjBxtAgt2MqLvnsoHN4z/N
wfZFo7cg5fgp/X94e6/eKNs8DQKDC4Hv2ZmO9XRWpqrRz74nTLc9E65yBDQi61ExLbWhsa/Bsv3G
FC6iKIZPw9bKo9Ph1g4fsXMLhPlwtBzEwKqoWlzd8u/ZkyyCdS2sSUfwp3liXT6RFDWNsgE8e/sL
svZvUTEHis89H5cblreEjGeIvB0VpuRF+HH0toZ87sRRtUNLhxC2hY8QtZFUBQdL4btdPIhYTP/8
j8Qc11bfUrNbjBGCqBCkuOnGj9XG0Nv3dqj4I7mZEU8IMOGOSz69YnU3fSNIiblWW3Yh3jjeyQTI
+uxWGnk8QsxiFimvePQ+V5NsbNUE4u6uszx+r1Zb0fPKWEB8J/2bTHHsuW14JurWpPMCDOgDIZZ4
IU9HLcKkA0z15OjCOsK2ANCcuoES5/TOXmweepwbDfm88KI9+iMx/AJ3MKaEdXGobjILdbjemOet
9j0prXl0X4UOnzuDyHyqWJM5U/FcO2xxh7Pyxu9XQFK/Ehb9ET4c97DxywgZ8OSE7Ionep6wtC2m
v35vBdW6CHcsV+a1zZlg2d6k10mW1tGN/YgKFlj0MUkcd4qnCVjoByGVxUwkLREhF84RZPEZSnSm
/M9vU/eIjlZKhwCdNEiDdM0Zl837td4jlHlsg1QMKWwop9pYMvs3hd9oTj7ryoxz8iZplLEoIIr1
BuqeQwhUS8CPN0w3o59a4UQwHd//aiZvKXkq0Ot2Wwlyc4hu/3W4/9fV9BWf/YZ7bzIqhnxJQlhq
9s8mpk7lpg6YJJSgmldJF5YjehXdCdfasUFPHa/xPXw77fk3EW+0ICJIIBcbTdE3tjNQXCLwcOWv
G6G0hm3Qlwc+zhxKT9PQzo7ydQl5RFWTSKBNZi4Yeuz5xSmgIq8ynBJ8k5c6HfalWjUKuRgFHG/J
6ia+ixWu88uvX2icTkgPvFo/k9P0/AIKMEDwLn8zuVxwvH57iPFJ7C+VkwHnHLmQGD+pem6vbTKj
PLQqKAbqUgBd9TJ5OsRf8RA2IdPJQVFe2Kn9Gu2blqVx+Bfr7v/GNDvDOJthzTNQPz9gElUAxT3H
dMcXwTi0aI0yPziaWtSjjjYa6bgEYMh8CDdnBsoas9ql6L0sd0FdNAE+/EFI4BSXCa6uMDUvPfgZ
CYb8my1zjQiF1lVdsNGR9mDrgnoZSoWHhgU6cJOqz0uKlr91i7emCvKVOGUXVuNgU2Eft3K3Xq/t
fwjONCe3LB85uejqnpTE90BPb89SXkPG98XcIu/4AD60qaDMHQn34RNNd0jcC990Y7CccZNjidO/
K14JhqDcKphkQW0gQ0HvREFqgWyatEhIZ15HjJJl/lEd7TneUvWip784RB6cTQYVu1Hpoaw7h1D8
kSQPTMq/qEr4G3CbpLTNFk1aptVYpwWH8eWEOgKMUPD7n7jE/9wC54zx5kF/HPJu+XOhbmuiqBNJ
QhFj5srgTvX7HnBuc88v3Ejvglg6ULs3BfeDRznVkt5Lpc2bIyHKaDNOtGi4CGaueS6PCqPIrsht
8ABKFLi8oBp/Avz3jGke5Yx4r1qut4UW2FvFC5oNcOCD2aevwq6YIBss+fwYDFEVYVnh5Z90ZxsM
xr6DpCb6VL1siW6+5iib+OGmDs8EuvVCDPVTeT1tVXgaYmgmz1yU49eWlYqP+BnyaopxlfFHfoil
+rLJgW5AjgUP6UjQQw3UY9K0WRfM23rX8vz6OyUxbCuz/LmYz1m/C5oTJUxraGHSFCdc3oKw3zTX
1lkKLy7lUrKtRmZxEeQO76PSsA6tn0cX9yQD0gqRsnzCspDrpQVV8/PFL0C4wQhyp5bNTYi4NCz7
2eyOz5fmSPV37tQsN80WLUwGDeOAcHE/u5PYXhY37MkIWC3Pdq3TWwoH8XEQhwju/ZjQphX76gOQ
qlQHyq/gVolD4Et5iyWIHvRKA8QbQ7jwfbxm+tDy+DBzODF56+meDR/mV8+TcSJQG85UkNp3zgE6
yMuuOBIetlO9eRMU00glGsqVFIsO4KRCApVDi2azMUR/c8Y0EEAeAK58La99yIqUaNOnj7kwKKCr
o5yHl+d2tdWw7YaW/LyjZrAxWAKk925enoB3XTSUpbRBARW27w/kxnIfOnzYTaReMhcy0p5zFq5s
qFVyXbKleoB9wHIJ9p9oLK7cGMt6eVW/Ld5p7ojzYiVdNpDg17nQ1kIitHF3cMhUvNLl26HL6Sze
Ndfl8uUEfHFdbW/5sAuR/Fh6HAWBzMZHX+6cknW4C8IYSpk4AJoRsCaASYJVxTMsVeQocxRDF1J7
RohE0rFcbqcilj2dgXxTKauaa0ZRbzg07IIg45KQ2/mYvzp1dk2jqmDbQ0qbBf8mOZotdklXA1Oq
LXyMcUDt9fYIp0iby1W6S5q4oxdqz6rZV9mwQl09YWf/dljujHgHt8xcWTFzIS2D+Dx8v4CVAWBY
cvKGcbzsDhGDc7oPlyUk084fb0TY0tdNQNUOXLx0QCRZAzYeOdho9Qirz69NVNlSeYRTcQfqLiUF
SQGz8aDBlLabBResRSSUUWtX0fNtKINxb8ZgarYCaAOhKH39Sg9TSvVKnXUvNoYUvRAcKpvM3POa
ID6lb2EI1fbyt1B3Xcb/XwGbJbqYvaLVUJvdznjqUaF+lb8WtIwrCLNrFkr+hLUsSG6WZU4Z5WB6
FfLzHTCw05RyQ2qy6jAQrI4kj+7GrH8DiIfV1/g3MH01364s48bqxui3D/VbjsV1rB8oQSa9vDlu
FWRDSeOR5TGZSj2ubBHom3lbeJOBD/Qyl3EruSkX/Ze9PJRrAg7aVb/l6FKhbe2CzaXwuPERtzXw
I2y7r25wb08GSEIWdK9M/P6GfwbzSq/OHxfXFmPjrohAE4mSRrWpBA011YZcSyVp38dNVuO2R92w
phT6F0AOHLcBBM/jMc8IbztG7iEHd2m51y2dJBYpZFonMIO/HO92lkwU4W+nFJgBKw9p9lOhIcEG
hs8ynTmqmPfX9FLAk5R00pT2/iLl3f00TkUSztYxy1Iw/dRN6Da1GNZw/bR9EkSMlohLY1sN/90a
HZ7w8qI1kFgBeuuPTiCirsEFRNPgeIq1oD01hktCy23b7ayiyggMbxS5Bpw0viHQxqMojXfVXa2Y
jhnG5rcq/jQUAp6uA66DGzZGlgXvrWlVkGiXbBydK2/P0iyIeu1A7Ww+CPJmwfe6mn455KfCBIFl
hqdovXUZBRegJg5QAASxR/KLHkS+fCf4X3sgDn++G6MhOICFl7eks7VdxWbdKsRo5U33/k2cOrfr
wD8fLmDAyMGWu7uiEtMB5lJkBWlUID1xhEz9sUpo0QSwV1+XLVcbvyU/VIVoErb8FlmlfgLYlR0L
vejzpi5CKL7VuMWIoNI0kYaf5P8tnBFdqp+QO1z6YXDEkhSD9TdkrRXf3dw0+qoCozeUIWcckKiv
oL3l2076l1ZlIz0+2mGPRodUjmFqySZFTrE28+AE8Ojd7Me6Fl6NfbZ5gs1HsH/B78vUXy94SEEm
gJRnCdVAjI7meBk0Sn2qnJFjxtY/InOpaVIDoI0uBjXeFLNd9iCwxFKJWvS6ANES+BRl9OVYZ4LF
9A9FFOWAT0LSxxE3AHZJRGxAMDZ28BpkT0sCIgoG2NaZp74AoVGcgnm6GqY4POGpFuWTGOlyC4Sn
tWm2yUHeUKrIOnhLAWuVxzDt5Pgg09ZVezybE5i5YzAhwJ1J0XyPAN79HQZ7l2njVAbtVxbinktG
n6AwBVOY9CjPOA0JOa63F9vtS/ZkUu4VNf0W3o1vaUfvoSj7M84g55rCPzU7276tujyONIA6fjwp
5McazzneP1VpcFh+GzZxU1tkmgc8YMx1SSAtGJNjLsbZWPrrqbJKL5KhiBrOanZHZvq7OOSVIEzG
UvNdfWRwBS+MRAA/Izz3kZoCAJwi9ak4YRpAXiA5td1ZAXyUTX8ujHUEtiKH5owFxlxLSBnegT6q
u/pcqZBFWWuCIN7sa72dIwZR/N2jpDXPAMFryEgP+V7PBRWE6jF1j09GSpclaIM17OG1nXRFENWH
sl2D7k/3APbci6sGld+bxmqtR7YGZU7W7gChAPnvLwrOqX+cLgi05nnaxA407AfFHHQScWXZinD+
NbOTXWWJPZSuB04xbfX/lO6VdEPEbEhQMO3oEMvbnTHiBgjf1c8AyhYGEjw7kbDgcoYME2fig7pF
ch7VsNHl97hGI842xMbneRNwpPJnc+gc6/qZedH73Tt0V6F0pPZMQt360HRn/3tSVJiSPTH9Ui0i
pWZTxbHEpSslAahyYAJzKEslprtidZ5V8gtXGoyJ4+PtrV7nHZd5OhVr5LhD7GDAmvsTPUPpCBpt
m4QxZ2YsyBCm2dZTgjmPk9kAirQnF4FsgEoqbVZc3LjFVT/g4RbsAg+ylKBxszwIRc2LU76W+zad
3sZU3K+xEzmq2wuuVbMubEx/7vPpY1G5JY0mLE0MJorMkPCtBfedai2rgcTX4joGQ/2nZ2KzjgzJ
in78ibXRJxp5eFeIiJw4bpoDhsg8Ko//xW+tHrao6XG4ryPExa3CwlXEPl4YgsKRW25k99Ha1DTZ
QlrWPO6kHEdYTx08LXxdWJDZq1vuZnH/fxrPdStccRraXfxoDEWp4hKG+3YVW/btnhNAGDoyqklH
Sij3QBvPh4/WAOAUuZsHpzhGOBR5g1Owyywr2aoxi1tP60VVKO1fFaaXFelkGvggJwaKykWCdLV8
R68L7R4hVny/URbVprl5cjD3HwRL0Ay82EcuqyFXf77FhKQL2za1vzaeH8mcSu1PcRA6B0AZN4xt
L7I/07gT7xVOppJclXg33OwSXFnZc8EqZC5xJ8N2VHGM9x3W6hy69euZvO2HBXPQxMdWrGqwLBGM
DfpufW4kzBmTmESZXjUilBFxhxcxy9CxQyHzV0xMpZBn6JPPGN+1aWmAbp8UvboG25oTmoCuIpdX
gkI5qKyNdPjbWgwza6yQ5oqVY5oNieqBL8fAYWMeIj7GY3NHHig7dqUv4aGAqa2FKR+u5xIrktuz
Q3dxZaxJtgYsFz9l/sbPni2quLVGySAG6jfyFmwk8boZ4c6bpQuDDJp9p7SnuRuJA5S/X02//rMI
wRSCjRBVHZskKd7QxP9qbabVZE1D9meMtfIFIlBGIOCSZn4wTyB5lDXrbsmjzIrlQzDKyRkftu5q
3nQIvYOgH/aSH7L+utLk1ihWqFBPaffxAgOAtfq2if0qI2CMtcrvKQQpcVVD/3pBmANhT5tPEB88
kRYR1DHab0QHJg1z/1UHAi6qoBUXi8wGx39CHas1C3Xw1F3Gz1/bsvu232dx+JLnBLcdQU9jfDiK
LOTEsBI58c4OBUXYXl7zvCkinfQIh4P9IIWdhseq6BNv29PYVGuMEpeMg5dhc4uAxHoKX9jcb36/
gCrCH/4U3S1e6lsPQ8xXJr7ca2AxcGkOkbrU8T4Ch4twQ5o6hI8wojnp7DTtz4H17xdmklOq2GDh
SWUBDxJ8St3HWCokPThZ6Gs1W5MQ41nlNNZ/fShlLyUvLHu0otMcm3D8ZLmsT9MRxdm36RoZZZoC
l+HCGBqAkM7g9Ik15EFfAFUI/NIrA0ao9LFFF+nSaOZFAlXYMgzyeeaHGIfGAWgKnHkyeS9kRCDQ
gMV2DIUWVsWSj4rj2rQFn++gxcquR+OtrsektiPllDsKLViwBWXDDDNVIR1jT+pmWhtZ2LI5qa+0
wiITCXKNiscDWcFjxAyuzcxktgccqf7VS6fbWW3wJvltdryELAkAaGrEUuhZnASBTIWdS9sXQYRi
nG2gXLS4TBpNV7JkgjW8PKG6ZvBP2riQHsafBwGwamWWCy+6wAweYGT93phOzyWJp9oamlWR1vXc
kiBpKIfye/8IFznTo+QoXWbCYDRyTB8OpZz3oSVjE9WvOY2XwZNrGZI4LPlHd0uTocVNyjKv4jX8
yt7hIUq+NOoBGajtKQ9rwq+bm0EgIk0KUsNFrqwtlDKXVXwGhRZPaDYMJ5K0js3TrI4ChbdsL3Da
Sfly7uxRIVTC4ApF9Dlx328Ty/X1+o4nmd0xMcsHsq1pnud1Nxweh0MYXGR2ZR71WkwUmiuIw6kZ
f/DSf5Awa1UR37L/U7jJsgKYDf8fmmzoi2NI2lVpTqyCFA9INKbBn3A6cRQ5G0nqIhzUv4Jnh7tG
Ad2blkiG+fsZuvXZL76LVSXOp+7UPyOUE0qHv5xSQ2ZezPPuZykoxOMh00rOCS6qIK8WwLbJkIMZ
a5W21UJq0FlUJBtysHAtSbJvwKcv3F7kJxrAdDrOT46Po9KdMM8KSyuhufulyrs+3g8mGRS3RKLa
85yFnfZIXM9e3Q1yIT1wN3fGO2tMrliN8ZW0/PqjMdabYOTwtUZrtB7B3PghQIw18s8l8bJreIud
VXiupLTGIuLe2v8WdilwEYyDjQhXwP1iM7sI/1duNRN2kcwL8eHOEq0mjiKcndeMMi46kdbzILtA
WdF2xiGYWKnCaL7XZtGiC1ztK+D9J3oRBr/KiZpbjwrPw2by26ZGKEGbLf7cNu6WKsJ66ukXjIX+
9jSXXbgdmCn4X7wMgfAW/KnI76tUxVVSsWdnSGgrzAiMlBblT5qh3oulkn6tG694I3WZQ8iBUE/z
hXaeqqNOFIaTyKJpSxhed1hfLMg8RU8NKZNRzbpsp+pKBdv5QvFUx4/bGeF7JDUorR3zkQB7nJWe
pFGXHSmCGXc4FgpV4sIcPkS6vvwJY5XEP9ungnIfPxOj6MSRC1bN8gFe4kcSJWpykfGVLzR4Z7Xm
WXFEtWuFBXxcR22ZsBpvRh5MWqV0SJ+5wRzfKkrhFOI7hzpZU550oVj99f1BVimhlUpRUGtwfDbL
t/OyjEtGhDJx5mlkDdXDXut295e1ufbkmea6ixY9YoHEiizk7in/xwCT9FVtiWaxRTzFjFT3yqau
CdE2yqq4WZDxOHmc1y7m/xtRhOvx3pSYLWvXmQpUlmA+vxc9LdVQIrCht5K3PvladKrayEuk/FNQ
BtWC88d5U1tUOOHk1hPkd9L1of4FwfKmgm1Msn7Ojmo0cL55Q4rPuXy1xLLNPM1M+GvE/K52XBbP
7UNcMuMvq1lyFA6Wkq4S3TwiFsABT7hOtytS9EqGlimjNVRhvlE0CxQclfESE9O3mCVcGVOr/y9W
IgMNkTqfmyYkPlcmLMRY3lJPnnbweJJrQOIv0uFyk0EF1mNDDUt6s0LRMRpK+syMXx9cGIFv/UQB
n6Cl868sx/hXQX9ZI+gPPJw8wlKkXlVWZdqNP9Kjr0ujCGEUL0gbTVXfIsd4WtCPoRE2UtcBVx9i
UcRWGEzmHj83ambJHRh8t40AQcpdaf0hY2mudQwpgPR52Ny9HTX7OE/Qze0tlgtD1rb+lXj2F1FA
as4pmpDP3IjgGZa+5bSF9zoqU79p3Z92+DlAP/WxACUs6YYSvuC50HWZPuamCVtqpmr1FD165kNH
pUDxe51eguq62FwPbCsweW1U8k9D8GKZ2P8x9L6wjSckJWJX7sR6hJDMw3y3irxhq4HsMcBfUq70
3GXOLlE9ERa8O8WqRRQuEogTJ/aBZk/92KPmC80bLg1KfS0VWWOu93AgEyOuiahQvyHTZ4CdBVGe
jdyjFLosM5d5DdXEWd/cGelOKjHnWFiokfg5y/zg3soQuaVdn0Eo+H2n4Ch3B9dsZuiA/mI8Kg8H
/tCFENPPbd93C6B4g3k24hYDOTjWfyXkAIZdn8vAFsI9TJuuqv5RfT0FcZDBb0NMEKTHDyJnSerl
ebEpkpetG+6rcUuCg2DtzsPqd2LMKyhCA5wa4MPdoaTDheHulcX78/H05di2DmotdI6PXW3NDUGi
FKGaVcIpC/Va1+Kk1HOjlDWVHFzFGsGqqGJpwIyULNuAug4lNiAhR6GWy86a+xUy8gyt8GAKgwQg
m1/1h/xRyPcSMDTtT7aWmry541RT8/vf/DQuNjkgH/7lRHpeTqHSCmxVOJ9FTZIqkdKs5RJN/Q7R
UuRBoKrJcDxIi3WEsdtdqCP5TBdlekdDk8sfteN/1E0P0BjWLBinqvnKAKTYDfqaMI8SUytRdMNk
TTOgpqwJaLTi1EgaqLNtVG949TensMTFUEbpnVHfSjR0r6c+MncY2wajf40cz7GeBsLiHHepbxu5
fdsiAdr6dSbWwPEDiwTUf1T6UTjER+mfJqg6xHHUIdsyZpqBY+TNtUyQsqp2RROUcRVzHv/AEXeq
Fi2IdlfAMiuvlalp5+XABwnZ5bdnjPE85vPDzkhbRujKPClqHITJ70QcKFBaX359oKC8pkL7icRs
BZ+860gIIVxhz9vXmuxlb0mSTkF/jZogq0fPeZBaqje0rlo3EMDxSD9Q03NWLVkzunPbpXUpIRaV
SQKdiNmCvNHEflRTeLIUj2ysyRMoIFHBrVYNkrZuF3Al2+GREmb+5IOU5hcMX7sihy4rrdl4lOeh
plRtrW+H74uzvZL0YYNhOP10dES+2qCZYdmOe25R4g9vxFEMnlEeugoZl+shFq5NA1JWAfhfa9aR
TjdZG/RDvoAupskoORW1cfsc7KRtF9kH8zbd3wcvWSnA7e2n3zizaKXy7kit9mkIS/UL6xHFUOvG
z7lLPnxe0dEyu0BjxWL3FShkk++fD0/wFy2/bHh8wsetHikiFktSnl9JtYr6eNslGerrW4lj1vFq
HG0xO+bknVe4gganSlhZRiRgGcMoH1mH7OlGjZru3iDZZ3rZOeJ+f6PMxmqNpp5K0nAiVo+qWo8s
Z8bhHSwERDD6+EWWH2uzLYR34OodHAFHakkFxptuMfsqsXMbLkCdZJ56tYC6ykhe9nV7TLO2OA4I
DXwRddzHDxT5oqzToGWyJRsmfZC04m2ZxTqAhSiF/57VVIps66VV2Hvq3Z/RpHJKRe5PFKr/hX0e
pw/CG6cpMTS2GdMSZj1yONvNacCS3r4uNkI/DUrO90o6i4sPX15xFls9Tli8Tcb7SQOGU5ze/YQS
2Uw2pqwUaomiNy3OLaC21i7rkmVhhoBniip7SyeZcsIaAIPhG2ijrWe9NWTtAT/4dbpOiH9Bodoo
a0Z8vxoQaGc81c6WwUty3Kfe4No7sKUpUlTjwABC/cgROJwWwqDO4yNe+wyrBVM5W6sLsSaB6YlR
kag4ASCks3sCWbPnBCUUaIvATNrhgq8Kvc3e46/nKdzGITL2078/a5SO7/DeuLn8/zpTSH7IRzuh
WPw0V3tRQMY19HKzdeMF6/TzgnbfxOYS13qULoMyJbe7skNctpR5ia0/TZGRF56IZBVfDlYAYC+p
rUjCJhz7HEf5PuL5RC6/qqQOl4SJMYrfgAXTE2PmU2p5eHXBJG+WeJfsnkfHXx/bEFXoExpfVWOt
7Mv/wg9Z4oTB8pM9ERljZmWvySKdTWPKNeFlHeFArH5G+u2TftGwDgTzd27XyMwY5lNPgdA93iWr
94rMmmQLNaZFrNqkyuGUOUOK5ABhd4xvR9qPTV9NHSQnD+09Urso9sK002QqpCPhd43hyuoWTpw/
escuey5fOFpT0wNX0O8D5sgz7MHJMJDHugsFt08jFt0D7t3xYsxNAZGRdr+rU6QRbSnSR7tX9/92
ugZyA5kFhbt4WSOMW2znqQJXxXdABfmdMiW6IitAQ1fBUQDidTLJRqAzNwrcw156pOHcO/vxqaSN
JW1YsOzLHj5JQ6YvpIYF7qRs/ssjw0KE8O8zPxEz4OjF8hoq5PYQUHFQn5ie1FQUQk/h7M0GvOYe
JYS5BdJVtftW7nGD2cXawlKKwlMh9BaVD6lyOOvtnBv6JB5joDYaFEakevJ6M9Audp41ttESCkzd
NdaQqB7RYU0kZ0KXHYvKeGrhJqeA5Lta5sMZidmubiyVguJ3veSTsPHOoKWPfU8mXwGjl2iDnoD8
+6wUUPdHgCkBbZMz8OmwScjy2+/qYlC8iJiEl1olcBrh5Hbo6E4WD2RTbQYYSMHpz/anTPcCYBbq
Xdj+g30ACzraZ1InDrfwdnoGu9J+IumNmRkdIrMt1+q/SYAt30Ob/3h6NMlEMqFtuxxWA1GriIgc
UlguIpZYS0Vpa95LPJHgdpbUHSY2P+jSGFBkbygr6L7xec/X2XO9LlLv9hq3YF6UG9GPt8rsJc8y
J5bCKLDDijD62Oj8yXcixy94Mv6Ubl1qPHLavKVE6880bcRr14yOytkaNWYRVO15ZMlKULXbqY9H
pqY562LkQ/dvry8AM4rDp8qNICcxhONdJMQ3FqXg87ekyWaMs748nlqnx+0GHhULAvIh2e3DUGLK
QlQYomV5H1d5YAVxcP/KKd4L6lQTEH+VibLm34Epn3QIQIBAFT5AIK6NytpVCFefzRif/kGADS5G
v86A6PzAcoJn1iFMWXxfQI8EccP3o7sVrhVk6lpTpRdCbTaVY8MbO0Z3GG3rKSUq7Zqtjp1hCBQA
EnfGWrv9Zry7UkhAoGBFPP1CjcNDYcV0CaiJKFxmDOuexLdsFnR1x+eRDfkr7rUWkKairYN+cfpI
dvE92ieHQ6KasOk5SQUFtP1iQEi861LCd2KAEFta1uZwNgJB2jaaieKbLUZ0LiwB434G9lBQl1So
Au733nkWQt8XUp7YhL6jTpbYp56lbYF8NfMQDumBM7+OxlGRvv9uNpl3xllNZjHyVv1dn4G3L45v
5IJDTfpzIaVrbtG8IYwJlRkmCJ/5FdWCG7mi+M/q1yAUhIACkvNiVNE0uxP3J1mVerV9wxu/nfOV
zqA+gpd3RXJ8QbBJCtP67ae5yN+AKVBhJ4skl0q7f3oL9mgf7JZEvc9gxJHWlN+o8NKy/I52Zr9q
Tlu8kDIdXwpnTOOzkIgnwPtBF4+y0LLNF+j/fVNEBKgUl3cSNgdLBgvOMDzMCJHD9jmZFuQVfbEw
5t6uzga/LCSuU5Iq0gfyK0iexwjhDA+N9CEjylxmGB66T/B1vHhsCvZoefX25m7SJn9oZK/nlSoL
wn5kN9kLqVws4+bbyEG2qZwOSZsOiRKVFsSOKFe5IvqU7EBbBjmlaUqJJTzPVlIcmLBDuzIt2yu6
mmYwbBbBxPDFDGI2puWWstU/xO6pjCG+Kp940FSwggVPQFS7OGVg1P2nDh7HJ15uOdVBg/bwQkUG
dplyX7YdAUrz7rgQR3HBttMCgT1dpeMNbKFZA+JzQf97ejQWzh94eqG+xAlhG/Mn6dizoOTeMldq
GqAD0mQf07OTVMFfVe9V9tNcx/ztxSwp6B5APtlKH0F7Ntq2vnyvPkn8pw5Nt8oCabHfiS/3NLsN
kKCT1wQ+RMPMblw5PtrFGtwpTGM8NLNWQwjLTswQ/Yp/mkv6zZvfhCwo51cpvppizKeFGcBRoxVK
P8+1L1HKoAlKk3dzEJ6Otlw8yAdyWRdG7WMWOnC7b2xlclqoJxy0eB9hQrHuomMz/t+BngXCGlHO
9pboaYfvFi2hqL1Q8pkIyJ/qQNBw5+YUBniGGdwYaEm1lp14cryK4iCPUuSrq/f7DbWR3IlEWt6X
A8BnlpPNeAFQ8sFnkPUxKJXfpZ22Mv57d+Ar2yT1bGQSrWLiUxxPqG0RqBrKjmWy2UXw8kObwq2T
vwRp2HP1vJS4bwMMsl6QKhrBpJ0+69eyQyN87wv12iRrUTYktgHpMvrMsxmzNJ4P9r0majVnuQHq
1d5MlmB6TTuD5IVYgf0Q/Zgh2PotJMnbGJG16wRMVCv3bQvGllxUN2gjI5O3J0nW88OMgZM6tPiC
Iw4dYy2UY4zVUoRcGOKSIYIi4k1TeuYskE7URVBvoSQeO01vGp5Q/9N06th7JkSKgJdVR52sbaxU
Rd1hctfzyQj9LkFveGPoGfMvah0HOhUWsn5j/uVy8GmO9SBMDIKKCOXFILNa1d1KYDZesnud4iKh
WSGXYT9oZrHXz94dxkVzjRdlqYsxC9McE6VnwrM6aJw8OgpTYz41978BpZzwZAzQs3JMi9bbgnJa
VKNYBtWq7J3glZinfUyT7dokP6FHWQvMsaB6UD4BcQ7KvZOMiBCQZ2g+W3/hm24CZaLK5awHwm6X
mJj0CX7WzIGW8TbbhM5ngGeBaodn3f/VqQJWdsCrSkMHQMfHNo/qwLQmev3hFyGwtt6Lx7q29t9A
SuBag5RWyPF+mVis9THEe7z6oeSgySPlskc9ECa0s2/5NqdBBheygyAJL7HkgSHffUjMdOwkBMcH
Eqvbxy+i79me3/G0qvZAKxzXF+jxjlAsB+evp6kBtYiwW+jNe474mvbDV+MbExAA5EhlaFue3WTB
OE2gSUqqhO7u8JVGBmSrVGaOmCn7IBBVgizVVgMbcVtyK/qwcuIhULjc1U15Nbd1QGyOb3TKAqZN
ucvmzyk5KyG/FYqp/JKtEurAfx9FEZRG5ZheVlpAlqcIv0XbY7UesHQT29bUwbdWRJYsKHGV2iYo
FsBmtp5P1B4cnPcto2Enu5L7rln1Bef3FaHKHlI/kBZ8/9kyGms5e8qElLnEOFKFLDrrKiLuIeXS
GTZeuJcR08jbjlpUq1SBQY46a+lO5NPkWrgJxal1HEbsJFvwqJ1gqoZiZ94/xCons9L39IO53aGx
lxHhC4Qt05ML8og79F5imaMWBVirfIK2E++MNXSJa3Xggi+Te797jgPuBjZa1mARz2Rs4pgWifhu
yTI1VIh2FZAcgwSrJmVH09ei9Kwsx4Qja5ROdK5AuTALzTUWky7czr2AudwzZqBPA5NMhfwOEIPW
6pnRmuYQJ2jPAWM+K7FCYO2KooQBGUyKR0gVqyPrt+KEfeRbjyBGUENcpXrRwOskW8n11CexjuWg
g+PYZR5aqFu0QGF2FKU2f+T/UMyoAokCtT/lg6twNvB/44lmmreqtjiQKlutESDUcPJ2qtws3iup
ZKkwcAkQalh6eIu8CRI6q5qVBMkjCbjA/oFU0vEe0VsxXGytwJRg72vogzwzBfAxVBjGCBMfjc3Q
yLj3B0CJENETJJJjWS7YlAEaQukosYxAefsWNQNKRDZXtwSPKJxrEndOCMwm4MT4vORHEwkMTG5W
CdjkAQkKoA3Hnx+lI4hULgo/CkwIdBtZigvVIMHCAC96JcKiWXkt0MW6xyR8/IjLDyiqpkn6uK+s
rAfGtCn/y/2uJYJB6M0znXKtwg2uQVYFMNleNSTsmZiOlyPwEFneHYmsI4EAD2T7AnhLarDmc+VQ
uYP/qsPoq2l2mJCD9ML4P0J54Jb/EWzvwXtb3TCgJB8IAXWL79Cqn0QvK8ndY22AEpLtdAXX/VN8
ZPEQAY+KUCtTHdPTQxxa4/ivnl78lJq5WydxHLQv0b7h4fJJ0aAlqEHfCZjIo2J+yKXdKrQpKT14
f94MVXqC5c0lIV4IQBUHyCsHEN5CkV6/+r8OAFxpfTr7SBQJoks7+olj3Rjw9jfR/fEI3rPoCIYo
yP7B/rmgwJ9+uetAz0bQnEAev4gHgRWHJmmG2aNwo8XFbPG/3rAOXOUxDvNMUBAmaMGDJw2LCJZu
FsXBGXdxcUwFRWcEHvWxRj/bTZtVbEvUm++yMz29MaQWqurNZzQw51DeiY9SDrljN3e9waC4SNQL
kSGkTb+F9WTpPTNCLWySeRZiYPe9LglV9WSw3WIAfG83u27HUfSh6gLbjXfstIBbizGHO6sEi1ra
70vCuPVQzBhWwdmElYqUko+KvBYjEAXz0ZouNYPDMduzzYlUoIxbqSABYMbBmlEYuguy5/Y1MgE0
M2wB5C+tybNp52buubwAwXlapKCuOPGBtCkpD15AaN+1fv89XuAN8QEoikhw7WVxvyshweyuf8V6
Ibqcr77bxgZCUW51Rrbzhs6ucdGnMkNJqgxv2JZgZEsFgCak3+TC+kNSvV9D43FkfA/NvgCHbOuU
vgUFqzyfKhhre25fkmH9/AORmxtViXVXzJzqi26TBfLwIY4RM+ke29FgID10lCFZ/fPmwffnlMGw
rTAwx8vWPAquqoOUUZjJBh/tdqhyQ4YVXOhI+TFdN4SC9EniAwIxdWKx8BbX0X1YDSevaDy/5rLm
ZFE6BcAhliKderAoADF4cozL1PgrTRHVfdEGYl3avI60uViE/SK8446QxqX5Rp33EU2ZXBKynOmI
6GLv8wmBId06frjYfqGjNqF9RnHWtcU65k6ZyFUPsy7f57hQHJXcRv+XqxB766fKVRS7p9RJgzty
84fcZsd60YFj2YR1GQjk2sqnv2GkZOeSzHLC0avAHTiUpTGvqTfCupeqkmDid1h9FjqWztu8QVdy
sWV+XVAEpahRzRBhSJvZ8V535Pn842Q8pXwzsY2uJVhfQAK4h8wv3noYfpXwLqQkHugj4oZ1DNEL
ThTDh7nJkmB4gH47kgT6Vt3/02BcNrmADXpaoWXIMpSvyJBwg4KcCefSepy1JN5CmMYULR0uss7f
VW9M8+k0BiWllTVPvC1q1Me3VO9snxv4Kpr/9Grfue8rEW3ZgfPY8DgtVs0o6mSrcY0sUlDiIoAk
K04t6sloGCb9tEIX5CI8JfF1kFcHYjndQ5t6JfUGX1XnwBYArWQ0DXNtaCILlz6Cq8URkDy9PDFi
fa4wpje/YN9HvgYmaENMxEjuokX/164bZFaKufj1Ycc8xDTsCk/dXvV3CcRoSBaSffTIa2CXyHZ8
GKlMUN75EN5/dpa0VcqeImkTkrfg5YKClrYIFHi+c8IT+5+fTuEeCMIV+jU7opCPULZdXZhOVMb7
z876OMJ52534AnZALd4I8fiulleDjmuzRHTVff/ixbnNHbTF/ji4M+kJNWqTW1IzT/20eDsnmy4d
cqs/pIH2vLrTi8KpVqfc7L1FbUWk6dh7ntfgtBayCClWPQ6Skk4t7r6ugRkfIhVzBa63t0owST4b
CygHbopedCNVzoLx4/MJpkK2ZkRh45aNgOK0r/bOliPd9ytVujTiuQwH1FfFmQVb86ytshBxPcMQ
UUjJXy0+HJIIgE46NHNj3J+A+jQSewjd9kW8K8ejslhkyXqFRyhbWg5NJqOoWhvELK4TbJm574Xx
Yul7+PrIOL+E3O4Ixl7+H0LC6b7oWjA7MXLsAFPBU4o9svcKizQPuG3/VQaPT8zRYvxPa8p9P+pQ
wkkuE4MEW70zlC8toUBlrQlg5qXHIfjcpeQB8XNaU0AH6oAE8aSysPh6j7utW9PU5XEfJSNAnwym
gvrCvmPTkCXkuWRAod61QZBKIiAOIy74V3XOA+gSGzEFiTM16cawpC619Kxuo09d6iNIcBT41/Ik
EkDO+wCkhSyQ47/TtW0cnyWQ4XVwwGm0X00NNoh9gN9cp2PVd2V/wMaTUXKgTACmQ0xpzq2aqk/C
XX6cYgabTHp0WzjdgFvctVtWDDuJrC/jP7uqxUwAsGevD5fz5Q7MqkpsrJO0qEDaphZA5kh3vWPA
2i4d7yULJhihR91NSetdoZGraW3X+NAJgIzxopb+JjN/n1yJsxP9wWYCWQtQCMg4tOs1EhC1H9GU
S4jdBRa98nvkDfaNLy/MwTDyVgjlBsC7CnIA7uqTIL0IXnCYx04x1KDh1vVcypSY+CXA7kPbh7jk
/lFTXgX43omRBi5kM4rzUFvJ8MwJC5k0UbbdGgAnYLurA/fjUfn3pJzXvfGJMhY3Yxx8uR0jcWxq
nKQLhkrWp5wFFr5O3/1Trman4vAniVNMC4/tV2fubNetTE49HVfEZw4/mJzjNf79CmYKe9TRkCcZ
oiqYocIuL0j9eVxpDXKXSTqQkO97E7VJV20wKVsWXik0NH/M0dVRbCY6LRjB8PDQ6Huud2SKhWWT
QBT6Z2bnqvBf4L/sNZP9weNG1A5jDpWL0DOtGH1chAof1wZb5/1D3YLnhn7wWAW4PlR6Wf42oN6q
oNWx54Y6MrhHZ9tKDr3dk1j3M4uReokx45AboB2883B7vV31IK6O62PjK1fiFEWD7FQP9a/RU+IC
CmgYoYl95tpeDhwrRNp6qDTC2xjKD/CFRCPb+4gAUbvn8rzs4JkuR956+XAY/iMR7PGOCLjOM+tc
4zQ5f56yAEEqyTIKLCqJWYHB+h7RO/PP6ucSmPQ8ohixvYF+n0kvDtWgKanBYUq23yIWzMYpIvpm
kqkB8XWHdL87G9x3gQAAd4RCMhpp+bQo0CgAHmPYtp7SVteWi6UL63k69RqN8vEJFk7JVUNwFj5m
fNhQmTwR1c4pxGjtnNeUCBKi+vWjIIgJUcG789O+UdS5lj2IiCutCidQW9SRmPhrF0C3wlt3Uzfi
psf9BY7HmQkjs4Bc4PHhMA8WuFo3bkp60LPzlY4XdDNimq5J5CVwbcEPufOI8Q6L4SBBI4XGD/NP
ghWq5YcklgXNsX/7z4opFgPopc5oalA2KQPfSqcWi2JMKpmfRLtdNPxVXQhrX8ka0t5w4+jlfYhN
K3KiM/6oJ9Tmj+6f7Pf0JaFAfcDuGXpC/tEslJcioyGLKxy3uPoyjEEO1+AA4gPUZn3DFw8iBjFt
6vmpeyMwbPJPMRC+qusIALdT1QOoZnv5pXcWzCweWuAa4UDKy4hLbizt0XLeP2VTranSoSC/08Fv
nmm94MiK6LMwwTzuqEq/lkVRkZo8WS2mAeG5nEsVFBFwIghYeEl+lUMqyMU3U2l/yIU/mrEBD+p3
XluwZdzyfnvSHXJiBuFGjcIQmTxE0tQ4L+eGz/W8Vps/xKxRasDeCXMxhScGrGC4a2DL0+5rv/pe
m32AhWbz07aHlN2LGAn5eu4Um0LAEfcfyRgORMvdQL0O+Xr6onXwHVW5gIOt96VMOn8TxVVOdmxL
Z9VomlOVgkE6CPyFAnmlgnmRTq6Mb44+jTREN7SaN4wAPeTTC79BfRntFUl/jnJK39ZUz7DvvzLv
BJa+xGNOeLSLG93I1GliLoMrZ9eYGlDxEyOzCvkYWulLj1K4r+3lVFtJl2YDzc8F1E0b7osBa0j/
/T7fmKpYBBpXbae1gw1dh/O8A8xsSgSAZimjmZVAfVCw1pRoKkWlrR6HYpB7ys4wHMk6Unf4nqVc
Ff2StW7uyOfuqAVWg/r+MuqYV/TTE5QVtiF8YA2231ogBQCf5zlXu5ouR7nIMYtg5S67DN5rC/Jy
mi9Fuo1AKqGHZSVTzAweDkkLIwj/B4XRO9l9CU6oQxGEFXSXvyr+m/IeY+8OLqLVM1ClJEsoAj7r
zK4Wc4Vjul9DMAgY+hqPpU/YRzJgzKgbO77pkarGw0QEq8H3lBOs+VCv5o83UVofZaTQUMzqjUh/
HbLWd/SxKLJhaea0gLRZO81CU1uNUgAfXiGj1YK74wkf5whSJNltT8MK+i2NEW2iArVI8bnsfluM
anQONnR5M0YPjheRcAeN0fYYmy2oCe60AN7rOBhibNVJK7mnxd5bI8Zcz+S5+/PWMbST8+e27DQb
MoptAz9CJh8mlY1uL29sUEkQUJAtwDOZATk7Y1KRqx/MMI/TnJNHIju7SwYDJq6duK2lA6il6PFz
ZlrnoTf6+erqT5W3bNP3je3pEpS6cOhi5W0epXFNDut1WfA/2eK1vpXvamyEl2+w18JEJuEp8unk
KVxclpD2Pen2wpUskiqLvIoicd/5OuExrTjZx7gHIV943HoBy+1wUGKYJ8W6IAZHOxOmgXchQHa9
kGqsoIf8DRayXp60x7BAt4FbOoLWg0o+An5W2iISrA7v+7BW+9k+jZpzRz52oRvgr0stjaM5oDQ6
oByA6ntD0hoEGR26nUUwY+QX7DXKMXPjgBzVflAnQN/SLbdMfW/EbuINTQgSRCZZ+QH67XIzcU9+
5YQXAwfna1WLWiY9HRTY3AGthlITBoftvpi33n77HeypM6hc+h1DzWQPQg4OzhauVncz/sibtPe1
wXUmTGpOsXh0FUujsd2Ljj3PiHHxzARl0hTCCv0BjklRPsYJ4Z1DcZQLuqtibZjfIlbxd1I3F6nc
ByWe5MjyCdXB77POeT43sj6oJwxm+wM4OIphPAro1nebYANBhwRtjspv6Ind3Y5i18KDOsjpyd+k
m+lcHXfRytVUi0lXxs0rhz+jz4moOg2yhfZmRnnAOTzILWkTwzfYpz5oVO/QF7Sk6U7LCcxp/9Rq
46V7tOkwPQOWcC8rWTz9UXO6MrLwSVOS4k3LL/L2waaanl30DC4qGfF5FnPkjYyvod0VXPz6FpLD
FknPE5HxvMWQg8opU5d6Pe37ugOtLMivv9SobFEVwq7EVl48TtX3pZFUX6M7qYojYj8MTakMt+6B
zlRHtjqK5FCogZD7bsoxRLEja14k/+N0acnU/0bP/aBMdCCkRw2fU28FdtfjfCp/fOyol7hcLubV
g1qX7bK3oMcDYb7dmO/CFVjkRwn8t7+7qp2DP3XKmHMe2F4cgwmrHPJis8DJtisO6pVxDLHO4C0X
mrw2vL2OU3h+YXFnBjCFIhrqDc6Rlik6XINXj+e+8eTYWeefP+I3ZODp01zqtLe2+y28nncn30fb
32iBaxqLLgD+ZyZ7f/L1lRCP8utw/8g/moauOq5txOcISPYofotpaen00YkSFoqsPEUbyq3nwFnd
b3OlPCepC+VJBsXAfhiPqwtSyiJpTwrGJxRX859HdlsmM/kd7B3mfmFWA0y5x3BO6/zhd1qqojh4
O1D54a0UJfukA7YILrN0q63Jltq73aBN3Pnc/Wg+JkXTNGHxbXYvxfclomKoG1Q2m1egBHmH3/2V
KpKrePYjcdJ9noLTpIS3Uf6vMF3qBPeE1ZbjPQ/tmBk3ZtRGXI9r+jd57nhp5sS/yWS0b5zm42D8
IFRtmGbXhwUxVXg8ythUyE/yvvDjGscDTJHMkbgNBD1MNaiinqOItuyjaXVUoYyJmlGSGpU+0gRF
LxTvtfuPpy+Sbr+iUI3DRLREbopsatXyjLvLujVsXQ1zOOJguTqM1U0IwiCK8VcAKMgPxurCZRxm
MHiQEgam778DhInHVPkc92sah1Tj9siyrv3RrDhMBsvL8zTm0f2NZtNNWP3U2DWOs4GOBeDTTrMF
KqiwiPL8MuKnFTJmc3WhIqB46pJ5SyTMjnH0+6A+UtIV3vtVyZC2XgNK8ra7rrWAbytWD3lIXijo
iA+s4s++YZGFb6Ftq+nuBq6Kvoon3+7N5Von4rnUlbxi81d0DoZXIUlbWcerqIAn/drXE2g1pJ1V
ysc/g0xBiOCI0cVfzPpcn719mT22cDfQQI/bsXRspJNPDZdQhxaqsRmOOBkvYnFpb1wyFYnA4GkU
0HEwkCZKinBnIf0jPuM4uSkm1j8BvVncIkEDczn4QnpNXon84ziMcecDQCtMy01cZwZ1SlfwYYE/
DkAjdKc1drn09Q8JEA68GOIdafQZoQxgDm5qq+hBsBXmc43UYpn5LuXyEYBVmZJoDED4kl2zw61V
WHGZA/DZEYSUt9kxl5dUDp6/zisogKEVefNOTebeZEUnS1IltpvP+6Ot7YFr9t9E+h7EVatTHk0U
tqKSCN9ZoQ3ue2QVOHyqOzkM74b5c03C7RG3oIhPR7T/DgBWWIE2hqwAzr4i05qTG9I8UXPARUDa
2juPMGtDenTRnpHZ2K5Wgjycv1RQIxlmqKQL+bP56eWPgUvpyOmV4sUp2voLtEYQZ87UiTo+I/Sr
9jya+ZeDIcY3+lSeoIVrk72WEoTqB8SpiIsxa1IH9ykkEmlucGNFw2+VslHFk+sKHDWoHUxO/4U5
xRzFsVj6qdla8yKuUAeqK8SDYIps1X9uVy08sXjk7QBnmvM5pzwMz216JjGBM6oOmMPtsNbDKfjx
MYdoV9mByGvtM+vkT+GMpwM6IjI7npyqXLewjvms1RStGpIzA5lBGRCYqND80O3xi4Tiv3qqHalb
wkaDqMYmcTVoDmOwiXJ6PLLCqdMASMpGCUF2auR869qNmRw0HNQa98Arnwpr2OBJa+laJBsFk43N
gYBvORA7U3Ayk8+lTB5bxLPJxzzhSBxP0D2tD7CeiHt+s1pSxvWGZW8HRnWV5ACr+G1CoAep1IZf
gnKsT0jtcN71EPfQZs0YXil78+yJBMuA+xx65zw8CGDpHaQ49jw0UMrHu4557j/G8Py3EIvb5ukF
e1uPwfsnx2nvjMfQLLY/JzdRe4e1vyO/k5fzuC1eKjk3GRxsojukUk6Ja49RWE1EsHExLnhopA8Q
eZ0QL5Av7BavtkafgZeFoA0ABH6FRQRMhFGehRDL4pYMiRRL6aJfEmHelAt/SwHtaBNd8g0vS+Go
26S4CRrZmZxW7Ksy1ik/UXPOQRZEyL8kRGVoim2W+RETP0RyXktsh06FIl1JM25yUuJOSKRvBhk/
aMQNkM2dgLVa9hlg6zwPbOozUQX0gagaaVEa1s87YvrOk3fdRgDvuMXnqBKfZOH75tikeza3yKmt
DsB/NvnZ3Zdc5sb9/20axe6O4sCTWChG6NlgreiOtV4ISjfSA3MBJ28b8bgNUaWLnkZOUeowW1ce
TZLwwP+2Q/tEyT57fq61asI6ZZiTXFT8sxa1y93XA3kU5KRo49wwxEqNNdGaiT6wdkaf1oANosc3
/8UtPIXKc5pbwNYEStuenWES4mUEPm2V7+KcZRIkeDmozrH6gquHYGwoWEFdSbC0zN2e+p3e9gqV
LFobaiiAaEUmbvNIzvxIkEXMi6GYZWECvr0oeNrobOIdFB4YIQKil+4OuCC94hqDjq7PbkFKP06y
bLW7IcqCfCRfyW2hAVCww5Bt02UwT+BS7l/X6oX/ChwhI6hsJ2nH/ktgA/PCZkUeQSy9lcyhdy96
hhJll3HUme8pXrX5sZ+BHrCuqTANiIvpYt7SmwGGATUEIRbTwQev6Evn5HbVbQhxFJnaDswbsEt5
b/ufwJ0gj+TgJ28IZi27lQHE2nvFBlWVVtWWsbItK6HhPzN9umPz++vdHu3xAIpK5J/4XEAqokWF
5uNtLYUpzCtMRvmkAUkIi2X8+irrfLUohU+lN1NKlfeNCCJ0GRYLds6ROyX3KrtG0YgCv8Ah1uNa
f+cL6OK4JbgrZeLMN0kEUQ0won7x1k15XEk4jmeoyVBc63TxrhHuNRugLsrXgix0l64VTA2Dq+dL
kWU0aKCQpurkyCs6CBOm3daYgeyaq7CRFdCnEDOGp2Ek8Aua9Pmcqesf/cqRIC+CJ99veYA0K1JR
5cs+8oIRZsMepS1quZRC59B7SQ9LlirKdN7/OL0TZtLnOTr7g9WyfAMQ7za2ApgfLimeJm9/B68O
DmjD/pl49Kq8LIlzhBqU+pKPsBlMtXiSEFjONV65z7nulO1IaGUs8tCYzH3aiv9ieUaFKd9K5XsK
n0ebmyA4JEa9PG+i3aG9BuG9f++AcTKvc5U9Hh8SdQNo0OQaSvhJNfVVDs1Lmra45wPqxzHKKT+K
iGxgEMs/o/K3A7AD82Zp5PBEXHWWRxF18qkuh8MAV+tdNSVdbqydZYcL0+2vj8+OeqLu2GoScnZp
vid/xfQRUOPilLTDUDhVbVj0UMis4Tt9z8XApN+1nY4Wiy9KKTsiH/JL+jhPR5wZ/4ehv1xMQGPl
icGkVkkp1DbUWqhWyY/XlfulDmk6e+aRXBElPk/yeevI1OLWZwNUhsmkWkP2VkZNr2sIFguMImD1
m7v5IED6ea8kw0nQbfWL6OmdjVrjIX9JtJEf9ZlfYToFkHoDwbZs107AaTOM4J5AAy5w+9XV+bzg
MDx+chuCVyTefEC9GWr4TkYnsJFm5Tbrci9k2kMqC0RZV5bido2jgtK8OWvjeX93ltI9JaFjl1JS
ffxGmqYWQpFvgZPQIKx2Tuhw+MBtcv9a62kH758nN2V5bMHVzbyf5BfdFF3hQW9M01i7VEXGm4cT
5HhUObv0D+FmzfN1Dz0hl/smms/2SOQFE8lbMv/5P+Ki2dpaF1pW6kKplbyzgrmVRSHN9xMxzafX
Ib0IrzGTIvunNayYni93VXYSOO+3TLVnyIBChgET/ePQB2uc8VDAM+yqLQwarW0F14hGeEMtggV7
28M8KAk8vos6EllbMmwHmS+sQdmP9FNOE/2nYn+Ln0gn2WZVE0djyuA4QCqsQfwTzVgHTk1Qc1J4
vaJPGtytEL/sB9b6DessuuIrxkWQeVJa9lMvtDqQMA+vGQ/8EUq2wPL5AHFTrNXV6LmKmaeVev+o
FP+szwhR/fiXH/Uo4e1m8ILjIbVCXnh0mrkw5qeyAFIVOIerpmRRC7ylZpfP6YT+YM0+/MgWgkTj
4+/2ZUiLbB9NfVfKPWBdaTkbZgrpH6CJdG2Ye8G0GIMdXbEA/bKZBtEZxqXOjGsYUxC/IxxFQixt
8YINvcQmDCLrATHAGqts0RclSJcY0q+k1AbzYMYEdmEDSrTKCTtYdTg6/2iv8JGeUMnuQ0+mtMJW
0wdMCYl2eyR2qak7J231sv4pkqGTa0maUtVoH7OaZd1REKB4YCkoAZzmdwFW0b1RcTUa8BTmkAlg
+ohpokUWywAbYSvbK9tiLXcL2muI4t0/iHOiI9UBK3fYzgFKjGsTeu66OWdOnatWJfVYgSHmtcav
x/ee2qYgnXvOviCiX54Hh+A5lQkYIQ8RFlVnRT6iXCaRfUz2D5oSQXQlQ7VL0I/Hxpt7vL1qpFg5
81KI3Y3B959WWyDqt44N6ngB0u/OBloT0XWD4jo7mH6v55Os75pspKE+mBb1znPF7+nt0Eg75iRj
lQyOSGqdCNU6ZCKgCeGP/Cap2/90RQVzd/A71yhR/KirJCyRttZJuDxDj5HnImPh/qG+anPKOoGL
fyOtjtC5XUuOk8eGSromDNoVg2YTkR9TVG00QLJ9GMfxYzxRf+Kirte/buHuRuS7uH+M0fOB/U2R
dCB560rJoteOAOn03R8iniY4zIOfEalFRdj/aQyysmrK9BAdlxlZEuCLFSncRFDJw8dUkJzQZkuS
Nq4GPz3qJ9BZ6Z1qWuihmJ7DjSGwk9v38sQRYthKKV9dNlAHZAhNZ+R0ofqLdEYKUqnUIxM3ZEaN
Chqf3g3tltN+DvlnzEYrrNQgE81vI9Qrk6stmPopPBu5cgzqn3LyWzCqwZ1cJQu+BGAiM2Wed0c6
kwrmfL8n0/OJ/isyOXhisiQhWix85mMEzxM125przD+foxOeUJ8U1h0v89/PIbs/DYwzHwIHb2hx
CZZ3tG4lSq5wuXNF8sFqcGOtQJQJw4xsDcP9ZT8lIAZ6TmQ21FKLVaO2Ws4wbuaktx0QkRGgStXV
oWEkbOHTKYJcMAzuGWk+d1xxpumDI1QkzwM6gCCQkT46txWy7a39r2P1y4kuDfGR9abQ0Qfv8XxO
Q/ss+/K5PX1fXPIzyfLh5X/GUbuZdju5iNI3bv36thiwNdMyg/nRMe9NrMNSeEAcT3cs/W0q95qk
MBx+paJEXIkzgfOX2QezAvIxMwq+N8akxyc/WtQcfSh//kcwh/hWaYUqu6gwOx3VIwdeBHE/InUC
w7fzSdSvPnz8IUGUny2NFDEoZ1Cwwyf13BTvghSAKtwW0oJDffwkGkR9UE7hjqBiqY+nXgwN8ely
+8pFQyFpiu8O80VKafdFtGqeJuNwuJaOpPTgJXrkqcyzu9FFClJOcMgiNcgxSE/j0Mqtpf594Y9O
lULJbHfBSWo5jXDXzgGdGGVIn1ZU84aey02swX1+6OZ6U761Vj5r5ZV0MlxWiqof2ztXdXbee+s9
kpZRJuXBmrKQDFzarQNvYUGhKXN1Fi87jueOijv5/8bNDa839up2sL4uzbHLk7h6Me5xFVnPsyZd
wmBZkzHa8RqQLrN831S5GrBhdtQj23r6DamslHB7hJhspOoULxgg26sTVDsaRi5AT3w5vh4dTSh6
ved093EUyhpagE+yAu/wpedReW7pZoVoWKiPucC0lB+pmlP/RupgQB0cPxKOTh0xafBTJhB5Lbxx
Z+LoNmGLAUWOYSehSfugBdqgscSFDHCB95cGUaFnyIdiTL7chrU1AVwNpaf8x2dXVNcrwIa4F08d
/mjWBFlTLrL5VpBleh11JmpqfJODm79uuVLApMqRZV05wmeJfloWrd97vfb3rWMW0lZNpdBq5d3w
Qf+IR6qnHYQ0C7UB2WI5E942+6N47tJY/8Zki4KEGxq03ALp4yub8wasGl5n9/MoIvYnrs9PpnSL
7LD01QkdVRuA1MfC/7/HEmtgFLha9fVHdLRYFk8MTBv+u8/tnxrGXS8LrHo7Vl6bI6X3KaYPxGWD
HJFq+zp+0/HkY+pyA7jStydMgLLuow/wPklbKGKYtUkHpzbLptTnMHSbXqFJWkmoVuStgtrtdDaP
Gz35B8WiVQJXBKk0lpU4VWbL1FPVPWa1Vz6NDYPSFOkofP+CNj2U+Sp+sBWpGpQ/fqbzX0ne3QGP
t9WgGeI5XdMPvjljYZE2eGLa3uvQ5MCRyO84LUiN8GiLHrBPx10QZ1Y3PDTmS83hlvFYa4ersUXH
ON7hMEsnmooJYyQY1TegPKKeDKFvjP8w2XYgqBqLjjvkaX5BoJImnK6ZtUiubVhGwwCXQP2p9wEL
HT7r12i5KrewZ6AdAkP/Ehh7OosZLVZH0+cUjaC3cYUalnuuzdVXVVp35epqXxr8PHd52VGMad5I
+oWZArTSYsKAg4CSxUkVV3CD7Py21QIE7otSaVUwt1cTf2QmbfSDEcq0eFRL1FD3BEo/EQfwMgf5
Re3TfG0gcvgQGAzg0nfmDWaxF+AVUBSclG1Mb5rebavDxl9SKB3Z5giU0/xiT4KWcFyTr0qaAwKQ
wXcO1JLttXDA6U2Lgh0fxwfS2wLGjH1kPX7+teEqLY/Qf28HoqAf7ukaSaGMozOQri0XvUC2lLth
qXV9T0VEyyJJYhBNe6u4peG3UPpM5Silre6uar/+eMoZzR9m/IxvvpM9+9Klr1zXOnj534+R9IdA
rqB5SmD/+5WGdg5cJNbarOmb830SGQfxS+fNoGp0ISwnJpOSA9QqEAgYXgbSoiNHlVvTEHxtOXIf
6ltiR3zVpR0ovhN/WjGIxoOU7EJmShm+N1biXd3HtIKh6CH/d7bMNL2DM/j9QueCjHBxPQnH44hx
1fQLQFbPEq9lkBJE2KyonDwP5SkV79fet2nDpDgFvB9UFX8RL71PA1vfQhN6y92aOBlNAxqO0gEz
+QJf9rtdhGWkE/hotEnh/3taIaSV/wd6N7x+o6P72B1tT3sh6ZcFX3LQptVTpzUnkRZU6ZrOGoNJ
dhoLXB2tHCnk8FLoEhXTN8ouZmJyd9S0ZXZax6hDK5sjMJZ3yUOdQE7yUGcxpzhpDj3Uq2z8dQk2
b2n9SqAvUBKN9oL97w8btvzlzb2s2oatLSGYwjDAOanYiOKGbnLOR7YR/b76Z+x24KjQjC98M2Zr
iYT4YR9A1eWMAjJlGWcS4dwVDG3lrN49wvHM8tm2G9X4j9zs9GvXbNoMMleZQQ2G6m0za56ggi+X
FOItzHyOQoj3vPhdyO7f3ppAlWMaGGCmQf9ffF9HWa2XuOYO35vhEYjqFhKusGLrHG9q8AeAZaNo
oQubqdsYSt+y7Iyq8UeuYRWyL+9Ze1kICzP2NUCZAdhUXw362IdCZELi9XF9evw978OlODpGUEtG
SzfcNGJR/YvljKKnvSUE2Q4wSoQdhUgnVt7q4n4f7AU4CWT92kzs6U3QutgFZDAVmXNw7cN3BhI7
biAHOlhT0cBa+c7MtinMDbSh0Rqib7TLsPJY+myJ7B8CY/uQlBthQHoYkJQFzBFO0XcxrZ4zFz47
FT/5ArfTSac1eD5vI3lafAf/q7rSUAGX49Y3iKJG5HoHYLT7hNm+RfYY8U4vIxkwacgJHljL6FT0
XYjNMeR9rNeALjEpBhdnDbu2pmP4iVHLxiY8rXnc5EmuhWy076FcuOdtNF8l/u3K+LWXtpxvGy7M
0KbNRJEO21yBYpNzpW5widpArGzT+m1tSSUB1l5PxHUpaXrzgQ8SxXInU88PNlOxhV2Y1lz7fWSR
5vnIzZiQdHGmMokoBLvv51O5/edAPTLBr0uProvbW2EINBhuckI40XH4cc0F5ErSwj76EqSwSDDO
81g0XzSh8RyxDL3JFwA9mNLAgTOGLwRJVu+4GNqXyrpTfXmJh97/QaPHJ2Q+8Jkjn35AHM+yc/qI
37fd67Fq4yU4ywrnuHwDFEDlIJVMoYZNM0RFEuvECykFWpiSK7X2tbHa5R/AiTA5lwqgpppvll1P
J/unTJAnC97aMXeybT3hjvCEhBTwXlDOs7m39Lt08XIce5fvuwB3IrRN4HopWnmVz1h0YvsZkA8u
mGHjJU7iosbyv9TeBYjK+i0RU2uP1rpHzhr/a/urS7Tca8jsJFUFD7A8R8gzdQseCFreHVym1Aq6
fjrYn6a2T6gAounP6dJ5DD0aXpEov5/shXfYOSeHU2eacbqfYuLLhDB+7JYla/+4mPa7GBQpm20z
4XkRPyvU0gijTb0mscmM5Jgepa3FpCjkFyDkt2X8KmFXhPksrxfPLGp6DhndOP3CHAWfBV4G7rcF
JHl9qaQXM1UONuu6aBvHLgCBgZg+p7ZIT3tNySik1xbaKTkXBO7rykKPfg/FAgLC3riQe8q91eoQ
fV9Se/QdJ96gQd71csFTEZ6osgJXFnCKQWxQPWp6XnYCilTRSgQokHtIzEv8rR1Ajoo3Kt6GJe6Y
F/ZvV9PcGveAMmbvfwW87jiHgs06i7E6yDmdv/VolHLIL1CQA+E1Fs48B+jX4r6hKi7t6zX2Pzj8
8CRfgdW8QxuhrHwmW+niA5aFMSNknYSqoZoxOQfu20FVSSFo97Xj7j66f3dodLO3h1dmm4qF0IdA
TmaUtBIjJxPSk+SXwz15QnlL1cwe+THa6DGrGDCaGVMs4ESmQ8AgHeEdkR7pshshPNH3GIcvTYvc
Ma1kGAooBVyPPfljJnwm3lFYPtz90dZ/O+1dlk1kHOxKSa1jRk+EydshEdRKrcOYM0sqZkQ3n9ZV
ZTmfZpabFgFFochWocu+FCKP7kJ7RtiDcIG70SgEhxBe2BjuJG4zescKI9gmsE1BZtyRAouh25KA
qSyWYGJEexH6a/x9rtcI/pzO8BSPOwYOhCViWVo+GTR7UUzePIDFSsJ3UaBsP0ylc3u1R4pwYsEr
p3zKFHob3uURqXSfR6BierU0s4l9HFpkCzLiMxAzpA4ftkmoHGF3VU+tn3A7HrF05CtZr56JoRRe
rfYLxhi7nbmbcW+Q4TqPDg5Ip1jB6OIUltd7UjoYhsEFLLIaTneDksutoBHK01frZshf9pHslD20
VWKZq7UzuJ4cbFKiv+qhA3JNqUXYZv6iM++b5EvzLSFsdCR3gISR7zHXlBGgkxQtwV4lauJrZdVI
pdL1U7cxz2inUyNgFcUtDaX+VgnQiV0ihUd+W+4bN3X5DGEVel5B/17eUeuWGlR5nOvTaLfmXFbX
09Quz93uOXm2+6kpE++uDmiCO1XXNVSm+EtOTWv1bgpLUzUoL1wWA0CF0XmUVwXtAfPgRl8qLQcN
L3G895djsaC3HmmwxiG52Zj68isfXG9DrzmjU1V9UXHiEBBqSI4XJ6x3djsBHJx3GrD1TeUIF9Fe
GGcDboipPej2IlKJigmhnuXuvG6b7FjB+QF5qQfJ4sR2IJZP482RaqPwVjp4S8pBLUrpFcKb587I
yqjrU95B6ro34v6B08im2fUmeU3pAIiymhAsCl1260Cv29s1dZLPs4sJj5sL1VJrJAKazOpMugcj
Gi6mFtL5PLf8dCXe5hQ+0Cof4Y28Zqw27PSzYl7lP7JzJ12QrEn1qDpKOw2hUEWQOWVpBUp/u9PJ
UWG4UJ/Ju0LFJdCkfmBl8PPj1XSo8Ooax/46Nh8vrEryMNRpvIxdJXvUNkq1wcJj39wzQz9j1XoZ
l2s7gwuOpurl+DM4JS5MzjKMEWiG2smR0kph6IqOf2ezL4QOL5jMzDz1v0ShhbEMw9lcmEO5JPdx
UTRvUWa5AuWnZ8d+z/17LCvIev0tth0si+oZr9P0RA21DeZdigPnneFiJMRGP08pvLSHUIygDS99
diJbbPi4NzZwzqIMfzif3/1qsTuEhzO8KXzDVKJdVqgAQWXk0/2PEoHnoHm+4a7xSOt9KkPq0y8c
To9hH97wFrEczkC7IrhYIBJSVBOLLUdglYZ3wjp2o0wV4Uia96qr+hvDV+x69YsrE+02aqC6y5/0
+yp7JZn9J5YVKcostX4InkgidhjYCfLhhUcr4n+Zkbl7mNZO645/yFswxrpxjUzKPsPu0q+Y5eIt
FI75SpiFPXvKl5AiRanGSUikhnVB7fFBEdH6Z81vxhnBdh+ECQe+hj3D56zQ2GpPOnobl3wdDmVw
D1XnfSs1BvijxGwXX8v+CqmDis63R1e45VRR4JriNAtDViOkuCYZZkK8oF+yb6D8pGjVv9VD/tCs
JlyRfpmq/UdlLPPa/e3J2zt+SS/s7H2QVV/1H3NgUYBQTUrZ+y9+DV1shIrBGnVfsRpWOUul9hZx
rfWcq/v3sDgC0+DORCUc2Gv2wtz6jR7YAGVtsALd0m5wTVoI85Urw2jqKvZ2Y2kuCqugmipdR8U5
o+qI5N/I2WLYIUdUuq7vBA2vnqwvvNj/8foUhmML2B1Hx9ZTqIBVezqCNSJY5BDBD+j6ztANCZCD
Y73RnsUrR5zucyHHAGwIT2it4Vit7CzmCbxHePGqu8mAR3Q5bJOTbt2Llv4flAF3F52KwQoJ3UbO
oYDFYv5h2KizaShaUgja8hTeUvIASxcYw0jvBuG1Rqf9b2HVRd8mXzy/g1yYKQq//Wjbm4tHmCc1
LHU20Zh8lCCz7jVEt16r2Z+8JL2SQd1k5iu5+RT8L6q4lCu6F0MNB8t5fj8doiLuEoqwuQw30hNT
noI+GhE2s2Kjdiw0xcUYRLuWE+WXacKOi7jyDcKhDL76IrA0c4vo/D8r+lt1ido/4XRpigquwmDj
6OWI9/O6OZahL7YEWaOoK+3kK/sW+OGBYcdD5GI/YwKHUZ0ckUXSeGlLo59XqoBFup1o70jW60Ks
R3JwRZx1uGcixGjYXKIu/HSMFtmR+f49EChoxH7gI7BX2upcazqvYeSOmriV4ZmxMRTL8OOrSXkN
4uObb0o3+PcIJ61TTW6gziQS+RPcb9xlyD2MY/E2nRNikgGtnBLKGXFKAC7yLpE8SW2ATYh6+udF
sqSjg/dUf/U/ac1r9Zwljb5fx7BtWz+YST82HJCG79bv13XVOCJX81MpLGyQEpiu1An+aNTuDxJ0
Id1zoLHvwzeG5RA1M7Y4eMlvBDnN5ko7Z+oE1OI2ibKGQgItt9W2dxhJVETjVTo6PqSLaJFZKFTE
NIVUZwfvQDAUe7YgCeoEw/MlQH0Wo/J2W/kShNJIYoDPII+vO3ZAhrBxVWm26Y6utZvXETMx0yLI
Pwfqblkl2oGiCWJ+XY21uvBTiIUJsjE10sCowGgfKFrYPVEWvvyspBcNnC4w5peczAOBiTsBQGGp
6MGKfXWy4aqRx8lafep44gx4Ptj5hyQtuDkf1Rz8gb5PbAOVZ/t0yHuMuA+NMrdo1Ci2FSZxI9Sm
umTiWHx77tJ97pUZX7Zmdjiidc8pEKHID+j+IO3m6tFRCm/se8nIlveMMaVpFl8R3Mc7dzyIcX6G
pdjPlCNOeOYG6dMJCfPqFJkfNsoZI6tpBOL7ziLridNgJHE7Nl8c55IQtfe1dRbPjWmFwJXJfGoO
tQYttHAfn5/H2q7RFxOrmPlU/irFf/dhn55kHPnuIbAlx6mjF1Wd3tBrYVlRkWZQXyWzR03SgTeD
xKjfcWL/XKp1t4hIiquRJ2ERN5g17h1LR4uHv8MkptSe3fLyQmFpqnKtV3Aqg7iBnUcQmuiP+5v7
n04JqYTmqzbBb+ZcbO5emiW950kUXAbT09qhpGjuGFNi8FFcP0ofUxLBt44PmFI91KG6RsIiZTaB
0X6DIpfdkm3bUDzLswmZXegzrZZOptfx/KmTNMFdrez/aLzk5N1e1uwVqUhql/XBUC3ZkdbpIhDJ
a27YyMyeqigiEyO16W7amk3MV6UASiB/p6nSr3bLkNg1xTgMl7HyZnVlwyUvUkWKIZ19M+cecKrr
6QJDGJkjGxdNxGzHWcirVgB4ULhscdxaKLEI3cBBwfm0sTZ6YKa1gfwYqpPVy+ww4v4NKO44sg7u
4yvljlkeTE7/pMhSmOhUOnh+XfoyeSnwzJcKTaVCILPKBz99SX9l1VLGe+4STcgUpGn6u/QDxwyT
K1ncp3ePkM5NHr9+wJyT9Xo7a0bqJcTZWZ0TCkJAg8gtVjy36yXyd8R3/5XuzhEtrzkCnCuWBMUu
WjjC0Hh54pUBJJoYqqX2ic8Q7dKCy1daDlzTnASdUGrl5w7e6u04X7uvSqCMjVe10T9Z6qU3KbbL
j6qlj11m5+uV57p9WOGrFQs8ldR/XrbKAbwt/YX4riyr/T8Us7rYqvKoMvjtnta2QWU0onvzZV1v
3186n6oAa9j84caH0zzcUvVpUht/CDqLC8RNRelO/OEFpoPopr5e1dk8WFmVbUnYuWxdzMlzW3gZ
xZqPz5qg7A1WXQ7eAzNCBUOaapAmVejlQMcv8aaXXO1WrBBlK0kvkVrUcCOvoH5Uzx8yommoYyYd
xUmtcxnuQzch/gJo200kt97Ue9AIqxf0roOARGslj7LtjrJ0gukQ3bL6FHKODkAAu1Pr5Z4RdKjP
EyA68+Y28NPl9gwiceUVN7znmUGZUT8aVe7FzVcWgv+3/fkb9nrOTzMmMureHUSRRklwnw+f/XJ1
5VQQ06JlHclDHjkUgxjeaVXf/PclxTlXlKUGYd70fbf7sCJHtERP3a8MZt+tdyl8tcDnC0Y3tnDs
z3+doeGXVBBwDZGoNG8txXfLm1MqGBdsuIuNTvV8cR+gHMxkT6LifCxy5dmDl1D+G0JclfRYCUdS
3ZY4rYT2yFUBsogcLhnZZaLPeom4rM+xoW1jPEoMQTXEPuOtIVfNRGsXphARjwJhoD53FpAYIB42
8t2pBo6ktK+jxv0KB2p5RyHek7nn5N02jOIT71lHqIOkhcHhmonUdN5YjcXH6sclPHFhY3WqUQbu
NYyDFGvH/+XqX31OAO2E/DPZvGV9szhUiUWxxuwB93Rv3jf+h5TxqCdHfVIrF5zCAHfUMMPkh1Lh
/BrQgTWoqoD/s+ZmDX1mXUDHaTa8bhoBXsNwAjnH5gvxs30iN02GrX0ti3qnCpVa0em5SxLguSu0
gpFHrUTMeiNIefxsTY05WkeB+mf8ke9UgtIIupf+u/2Okp4DBfGwmRPjEMvD9XCmGvATjp4iWP6D
h1BiiOcu3nXnXdBwVM3l5Ox4AvTnLmjkNWzO9HZgLbmpXSl05B0wR/1kZ7VTcPV0FKGgD38bSMFZ
IAqj3nyqZ0o2dMnCvtNlhLLXJXbCZC+r/OXA1bBPno4ht2Sh79PCqH3DiTOBa6tZXQB/YcNQigD0
LLiRNHTcUd9EOiH0ROf7QaPrHwMiue3FVqKn06Chu8b6ZbP8blfCDSMreQAsf0i5QOr0Wx/hueNX
ca9GPi+UjX8NWjO5Udf3GzIlJHOucRGnR4ccFlfcl9euMznpiyvh4gyThXKA7RSR6nkQ/d/LI3Hw
eEdM4N3wq9lPmPoZLMReK32NrC4GWIDF0+NVUjF5djA9zTpjJTx+BSBVjMjW8JI7tOPSnnOVFiU7
TCu2elYhXy5I0Kv5f62zBNwbQx46dHr91VMEzLTk3+kYJ0oHuS7YpL7kSZZHIZWHrSTyI1YyX2Xr
VuXe5tOARsWqPAXel5VL6aii3kv1XdH4uvczaRYaJfndrif0KJliS9TKL4z7QtU9jt0mN12I0O+m
4WVO104MnARVA1TxcGPavQA9Z7C57LJvbbpaYRwJoUlOQe/hLX6gb5NOULvSKQpEQkuSBvA+0Ac2
Dtp64mr6mL7gGTXzFv8ibazTHIedp6GDeTaG2NqPptTsH0BPcr9FjFQ3yHHI+xwJImfEJg/UnICM
NzGFJQACTAeKV3HTeQJYe/Ljb9WCkxWQFdRGTEhmUexak2AdBmpC1ARoy3nHSD2w61NHrWlvRirP
wPcuFJJJGn8qPLOhc91Csayt/6zcBoAHzQs8SQy6aSlzIXshntGUqXxwZewU9efIx+GvS+BNNfso
aVozSu/MO70uV2Yk2z2d5rL90boN/kIQ5nfn7M8UTm/nHwfFtM+7O2c1ssNEtXQOVahVIrps6QLe
LeGH1LjoyIdLajdqOR88nGM0lDSn1YftDSMSyvWy4AQnOm9nGsxTWoiR3wnI/0ZcRx8tMJqPeBsm
ziJ5/u4E+xO0hIVehpGm41fjYuDL+eqZwj4baN1A0y1lrSACTjFKq8ldrKxaE1Q4CBDrwmwFPHzw
09ucRtD+R8Zqtc7cDqS3tC24IQESTWGHE0gMXlRvPSPL3f1n005CaTzK4O6S5HVC1LvoLMO7fpwd
uRTt8gewV1v6EpUT0uZCvQH6j73MCLv5Tp3qZca89wVGNZnQ2bIiNZ5YdsiE00ReEpPUTn+OpkwC
2cRS5TleTAba4Jo8NG1tuOy6aCHcWmlVQKZjgmZYeim2FJ4GGiYqzkObz0qxGEvmwDLbIEFcH1FV
NyCMj0lQ13HE06sWSqGSMMoFaYX7PAuPGTwa4hg77l/6UUKiKIDfSomaOnedGxZSZFSJQ6/8CHZs
Si9bFRNnCx+tx8WiLbv7k7YArz8fHYgH6vk8YkcTY37pzPm65JUZtMbU+57LhHCtfRlnttsQAjmf
EJvszGpfXmQjgnGwS/63JfltBA2zfdi5GcSvALeeR+syyfOkKA+FMwBwQAjHjSj0XjsvVcaomAtI
6SzfhxY6UJ5u1qPX1nkRONcOdkUsDvZSz04eR0Kpw2nHz9cEZlriL7H3PigPuSlI1b60nvk89Ups
aecVOPW/GVr0sCYlV1/w976fNYI/GUifuUhtqn3OrRtNMZnFGSv+2b8YvyoPjwF/QeRyUM8YS54P
KwzF2G2FAsRjzlj72JuvCGfkoaJ+7ThnSGyQZ9NKkP4ra6uo0XS2PeJVcV4zGUErdlbcgBRbyz65
FIeW3izhC6SpVcZfkXOFB6YIIPAIj13hDnuTUhpodYyISLkGq+YjijFxkmHaGnZgN15yHrvLHDJk
ef/2ZhkAR4i25jva3ZrDRgqqsJjvwOHOOqcZ+UjojgA4x4BocmwRJ6WyMTodJCWk62PoIxikRCUf
CWekkYTAI2N08KWcjq980A24i7yEo7//SshU83+n6jkcPL159yKUf9Jj+g4RW0YZoRVQOTqB2p1F
uT5ETJkcyUMqnitNUhE6X/IDmJVSWLo5mV+AnYZTvE+Bc989SM2ssCay27KyjTOeZ2d7iyKRJV3/
IRVn3vEhPC6zQ90r4hafgYsLQLuRE3G9WUgFGy9MN8wnT8O/GHRh79iwubo2IIZUh6rg036wj3dT
dIKd+N6d9Kz7eKwoRLZbP5Tuq+PH2r3A/HoaDXSX/C0lop9pKPuKnz02li+1i6axMe5abeDcBvqm
7fhmWyv9WPoP06SsKTOyVBnBZiuqMGUyUUy9OyRiAFs9ZwXcBPEoGSuwb/2AVTz7BSU7RYYR6s0A
xTy2y1RTNDw0cvnVdbY37hFIDflNP2te7Q/UZrhPYYKcM8eQpqBi7mi+yjjq/NTc4wg4sgd41zpZ
qOp+mcm40C5qQ06NNisvr0Bg7laEmxzEQg9PP4VPTbiGcg9C14YluVL+15xDAJ+YAxISHuSTK7iA
0Yke2jCB5Uk8GXVE77AiMK9AxnEWamwkm9uUT7xYB2BCu4g3/KiEPudFFhCQgdx7/AVynWdFvvPK
PTeFijfqLgmYaMcnFcJutJq7zCBdnq3Cufv1PpwgRvr4jGcKfVNPriZL5a1w+orhyEpbYp0Bwj0V
z4/U4vmBZTrv5AjqK34rKsNvfLSAv1JDUZm7DnuEJQW9bxg8WAElCkv+8Gv7i2YEgkXsYXJg1mDh
CzX+TQzoMc54/lRdVAW8aci0s4u1aODvEpYm0Bwwrs/YuTdbWZ3KcNk8HZRXayIpt78RUEjhiGuD
F+NHENE8zvoRByXC6viI2h+uwrmNY/p79t8CJvbSMrMZJUxokaIOwt6dLcfT/g98ocg3FEjARVaG
Sa8hGQSaEp+tf5JwFQkwTsNCj48H3fEMjU9leeWC3qcuXYFSSH6C0LDCVeYNHqMOsUfSSt0gCigh
9J7jE4885E1SOj6eipGtfJF45/ADABPtxul2uyhfnPZXrDJYJ20JBNKYh76hG3nSCtRse6N27m8n
3vyj6+fUg6ZkM7OYOPH+yT4kwAJOpUCl6cLsQxCG+dbp5ZbuFQ6LS+RkkVwz+4hU5wwNqHFBfhF6
Ri93Adj7Px4GWUB9fvPooF4xAgqXq78b4DSge/ofVtZSN4cbSxEgYSr6uxQsgSZrG/BK9vwEdU/u
SQAaagS28NIYYLTXEioo7r28G9iFseiNSP5lDST4mYvDKwWHO8NHqgidxK1HO4utBfnj2pINs/Jz
1HBf6MERQWJ8agOhWEbFH1dD//FsUrDz95J6ZA0B4UOB+SJA4KCRMzoijEQh1v7yLEFQLJn34ISd
X6qKVytDmMjeTjUWiQflzxXxM/odMi7pXqTMPy6QLvUVr1WKsMwLfa6Jy81xRcll0Vc8GpxywVcm
T8BtShcHu+/Od5u8EUMfmVqLQNPN021f6f8/gJ3qdyDq9wXEd7Y4a+A5pFeCRJBmVYdI17UAWo85
2l+frf8gVvDXyR8Ku7NOBMoyu4qBss0ZHgr+qPaVSyphdEjTLLBFtkuPzTbYu6YUGnE4vS0pPphZ
Ewxt4xsw/thfx7cgWlsl8agDvqCe6rAHk9hBo1x6DyYF3ltHKd3Wxqr876haQJi62nJGF1zSjxNF
k+5aGzvyFADxEZpha+I2cMTXG5xjZRewI1yGLG8aK8kYy5mw9PzccZaKl3LjXlfhKwXeHdFa1aNI
hOAKeJddxPFugd7pQlnJJYyg7DUk3MxaEU9OGE7RM+XkPjppaT4o/FN0PztJgGBUmbT2O6V6JOHt
K/hb5bSgqKORbJ+vOUdg2+iilkhJMKGAZhYMI+Yb4ltNfYFFjLpdIXqnfNDFRueaBUw5ZLSKspnA
cUXpWoNx6cfYyQ7CFKUPYSismbCy3h3V/ZCogoXjgd12pFGhl+onRHb+K1Pf0YD5uYjSdMI//p0K
54hBhivAMLD3bD/yrjGC7UrC33Iu2vTOHmaskASmlJ13C9chQxUHZt99jp7oQS0sHNV0dCIEKhl/
SRZPelyitIkCXp2gpJHHzB7RbZT39oDj3zK+4yZVLpzaHaqChc5gIkIwYpuuP09nHq1x5h0Clo2x
IWMn5Z8TwWjSmH5t31yCg+DrOYK5p5hB7L7FQmxuFdK4l2H2wg0Oo9ulcCD9W6hN2zgt/B47SADJ
ShkdsvoEE9r+5nlYCDiz9Gk+XYKRU6JcRNsaFNZVh1P1yxbwKeIP20jzDkLWcOijlSRrcGieulTC
xndC12a33aC+hX1yazwEwTQAgLrvH4mqdwTYmckdD2PlBkPBqxUidGWqk29ZTqp39bNfynW7yLXw
qxUfLD/6i0e7L24AsrmDmwYHoqJQf+wwD5LJvwA4GTgN6Xo3MYeOHd0atNWhHmd/z2n63BfbxvSg
fpKrvA3n1Oa7aNhr9zXBfzMiMFWb+5ExFNW2vzq+UUhyKwp/fLEEnG6XFzH/mVhr0cFUrOvQMkRd
6NOpf35qTAIqL4jb38d2+9/bulany2DltMGxKPalXKfP0Bmo8oL3nfuuR9jpfrA4vT4EpOib0OBC
CBgMFJ1AR20OWdBSqeL/L64mi5ZdETlCVEfFhqDEClmP0RE8MiODB1Sm4EI83OsA2rstlpreYLcT
lPnmYEse5IFtfEfR+lrMoSma86lKqEyj1oBwTwngb8H7a6ryg8R9yN2Onr20gFbtBV512dPsGeD/
I0HvZBkxv59eQ8ujPQEyuDTfuXDf1MHvLmKaxyCabsWHn3gNm9Z1zcNuh9cOChTaYjM8kHZmbut7
9wUjFCeCuDTcKWmlfOmdHSumIi6CyQMnfDfh2dE/dDOYCRk9m2knmd6ptBlnKfPszjNHov8fTlX+
z22pGXv7i+k6q/Hozl4mTmOzf+v+eD7Q8tBMFolvgWeXTsZA5ySj/WFxw5UKMjIK3l+OhEhSCL7s
An0cbUidub2rRDw7eFfI/YfSmAMWHRbQ759ihYXwsNbmf84T4I172KlqHUXGQT+UgQKECXZxvH/i
c6sIwVgprTrmjJWFRb3iEP/2AaZwJ3oh1WJsFCf50zDXfs6Dh2oJ9sbxzQp8vB37tAsnO6oqi3FF
GipDoAsCfCaWO+1sqSe54izMwkXBGqoI0uZToVtTST8hZn1oQLgkjBX5+5WXNfaURsd9GPWpRoKa
tnHwNZWD1cvaFJ6xZ9Vfx5Z//H98RtgTcsnNQ5bDHKct4PMJDI5tysHObr7LZTiizr+I142R+/zm
lpQ7UvUwoeV6ocSpnpYW068VnVo8EAOr+0h62EIzxFYJv6R2hwaEy6sfPru1Y8bKW5lLYmhg3PSM
MfHlGrkcndmHfsFYOKSLthjezcYE7aVVscz9bmOT9gBZSaV2oo9RrlCIBzWmmt//JD6NaqKnxWmz
OxsnU7516dxE7avHzl0UnAvo/6jxXKk2jF1xdHDDrt50wKR280nTKyREuZA63GK/02nzL643wjuz
p4VXKksetruRAV4IqPr2h0tMmZkGXWgJ3nQVip6UCNrXu2NntxQ6C5zKDo0ULROFPA8pewODt/ck
NtBKNQdFHopD2y3AUR8Tuqsr9uZzirW9VRvBdVSBwyhuZaGWiqfXi5yMpwedanspiGwqmpkfCdrD
1DVmSvlDj086oSpJ/ry6vDcEHrarhp82TrjpYm5NnTCSuY5J2C+RClZThkT0evKfXmW3sXkW4pgx
BTgHoeXUvaeazfcfFnOi9zKSjJDuQcyeyzS1HaaU6FZ0jtU9vwjnk5zUY6ksZm+idQNA5fyhsjvA
XjstK6IvcJ4UngSATzdk7qfQGkzGRAPd59zxoy7FLxscrv1pFj7BO0fwdc50ljNakQ1pbcBKIuxW
zfPkz8DMlkUyeYy9G8Wo1Z4nLWuVZ4qQnb7FSY+iwOTQfYenRg5kA0coK0lGtxseqY5oo9xEryme
Ib373th0vz8zJIl2kb7I4HoMBQ85BqMiNjn1NrkOFImfCP084XBLH5D2iZMBewDwOlohlR9JFxWd
14kusCuRWTp7foWsp6UJIPEQEqQFGggZGB0kdCZuMWafys9+BDnQuaKuDk2gtEe0U9yyEEpTAaNL
siufqhsCLEMAD9k/128mG/KPi8QESNQsU1LTv73mXb+Sw6hKyGIua70IufYpNiUN5NsY4VjGFSli
B0Tp7j78ne0nXvfixzO6Y3aFDNMNYwGUcRdbqzRkoj9AadfN3lOK6Z8jFAw/2+/hy3Q2pVSzPKvr
OISpg61vsgCRGjpvQKpzPoB9vcA+Sb32+49q6EuQ0HzmCO7N+GBDRuHf92+H+7RoLac09eIHtapD
fq7VYfzlNJ+b+iX8MS7HHS/SMUarGRqG2I5fvJ5pIFnOf9yk62OVA/acr13sMPMJqBkEjB/g9tAF
89twO2KzQe0OVPTwR9vIimO7lDlrloUOSjsrtGr1NI79F6twabEhLWzMs6IzyGjxM0MvmOW0ccBG
qsvDBosxYwb3EQ7mD6aBhRGmJaOGOBzW94SmJDJiJLR1OwX0nnazeul3BWW8QvLs29Khl+uP5nMd
JFKKGMc8cs/t7duBFy3brti9LLdqtYRU5XorQtwhaz5kbBGyqco/n1LIdHQ2+QIqYKXMjpki40xe
E0gWZ/5+JhjrNsaIOH5u26q+F/YzXsJtkAY7C8SvNrKKmr/1wBROSBRE6ldZb7VQjDe/p6V4SH+W
IIRQzjT6X3y+yJN2dyNa5RU2EY2+83AiooMIgetDH9cmtB60kj623MrHVYMcoUT/ynyNQkeMP7uo
2jkYRRkKyOxZP2aFOi09Vp1eHjSUOtJPXB5K5nZHRnNp8vpDztjglarpWOojBKLnvyHSwVo4STbA
JytGf24vHaY3DPcpfIDJ+uc3u9pZtzIvkV5txBHYuqoT/TtRd3H5o+DFAr7av566nityJxV7xWb+
TvPyfgAV9WwAZNkeaR+i/vyun8sUBqeh8BoS34x+Up8awLsBmVBQuUeE3tJVboy43LZfs0CEeuZF
iXi+/2TVcKTNP+syd/1WQSKWnbXHEddN6ax9dMOcgX170j5GVtOYLjWeErf0lJC6GqhIUNTG9HVZ
w4w/14t7bAYlgcwu15uXC2fuCyUHIJAj1pHwDzyyWI1AqDaBC+xt5vMYJvcVpL1diZPXNOgs94Ht
CIto7Gv5TsbaXJs51gSSNWhdQBAKkp96La7vawrqt036+Fpkmz5p8AJCvCiBfoLbHM24UX1PaONw
HC+YfsRtInSNU+oNwkwVCKD9Hw0gE9onRkpXfM4UnbCp4E4DIeaUwpK1eJ+0M21VgX0/LNN3mo23
esbIK/V8uuxszBBQVNKosNXdvYwFyQjfygfLeWStF2lSuz8n6bxrxGRg9z3TwhijJ0cRg4nLAWhf
xvcoZdj/4BfgGPEOJ1DouQWLOF1xiLfmIgBVmlRK62l26yFQB10yt+zkgNeZ6aq6chq/rScjATMc
00f0oVw4wY/5n3+S6O6OQt8joQab5PKOCtgjEdvqfIJhdBA7VXsTOkgVv0o1o4qlXRJquoQ3X5pV
a8OdMrkcZNZLOkK361uUTKmIaffvsJKgChgkG9APXUmXqm4B8ltuBjnHV0osIb0tadYGifhe9phJ
up4pgTQqU3uDDj/gg4XeoBZVeiLn5Gv8evhGIekHoOGNFWgMxLpl+dbF8cwVwmmZfTrI/5FDy5nf
DlCFWzQ6SllCv5HjVAgWiMf7wUylGkveiP7LUad1nDJmZ2hnKINM5EWoc3x/tSG+jOfmpR92JMyW
EuZN3YjkQd5fKYTF88+XOYHgzAhHECQCsikJyUPXMfO/yClSGlm8kQ/P5Mrxe9ws1NYL8bThtY3l
rYsAB9goR2VpCI7RoxJXHoA79oMqvgjVvS9KzmGOyX5vy0sqFux4p8QiGOfs1aw6FiAiqoI8dTy8
ZHpChUfqooZ2ChNjNpvEPOr5InU/ktdIixvcSEcABYtE+nJn8IYdh75LTvihKF2PUu1E5+j6Y1Lx
jJnLP/PZdxB3LqqY3PxLegVHlF5jWefiGv/NHXW3iOMC9PwfmXQkxs9UePpfz4EQC5K2O8sANe2M
8/2VU4t2Jws/vKUx5EL1sW34MJiQGO7dubQsu3EUUA0zW1KrtXzxzKrAU98zw9C0+789JaxrDW51
2ip07Q3tNFbIAGhZ+8knJ+tWYnhveSvlvYJjCsL5f8iqGxz42nhR7OGJs6FJmolP+7VIZ7Cz/yNw
O3ZJPHzaW8SXnxPSfY4jucqrQU8RWX232oM+njhPmL6IvzJUxfodyL/0VQrpaPgH0hoYpj7vpwdu
M5jeIlir0GRV1eRuMNj3cx993wlnW6sFi34Q/lD3AtD4r61pGlQl9hISc2LMdU9pr2T/gRHE7cYs
b1IoavOjHNNlTdEAfP5lBtyWN5E0FLEdGRF+w/Sgd7Thfvtf5GJXOFaOjNV55wudh1I9Q9vjH03v
ZyTiGm2sCgNcKin4nbl0yUWOQpQ6Ql833G0Ea2/IC7Fjs1iNd4CWjjA0LccVPrFhOfYouqWrHWBA
iai3lL/sI059O9AYoumGJeFphWQL7VmduREv9hXG5+IgIfnIcOGC8A4N8cfX4j5fCXqxkN7jY1Y6
Fe0AwBfB08mQdkPKQEs9EYahSfRUDltCjI/b+FRQpquzwGne4qC8WjZBTCAXh8aXcEjalYObcty8
9deUCiBUz/w8LRSThjO84dE7uDU6JiqKwGKfQwWwslCfmPAGKU8T6QY3v2n28LAfs3z2UvR+pjh3
nr3kzE9vKEsYBeGJXdkmcjFpHIkDI/A2Pb5jlhwEmLw7jtOSeRcgFX3WCZfgkGfg2/cLiVdctEFv
K4KRqr3R+ErIIPnhBcN6xrd/OMfqIn+JHqD3chtft6qsNDDo9QZmc8hCRqaK9NelX077pCH5cDWf
EtP/lFzhu+aMjDtCzbfo7yGe5oh0axZOtGYZb+75eXvO+FJhvOwQIplhbHI0WKRta46YKAJnzChs
8irT7itIX9KwGZe+crBVJKgOtKEBZO1JxKPCEGPLdvlTH8VBv/lRu7oWLgQX+D4Swze6dpIusmus
1yYGi14S8gSyf7eLjnqKvZeGe+nfCse6Z6BSyqzc+/+NaIb3phwfGC7T+TOpmJtHCGkVpaxGIBgm
1xEIV/qzVnvRjsCsnpUtKXLwSgjMO+Rl6uk8l5AdIkLiT/VLmL3N92bbpe6QF+dOFqS5KE2gGysQ
BQyJ7Q+9HNqTt3LV7CB7bjGso8JOUzBIir2z4pyWOjSge+f4gVFaG4wSFElpKn55s84m9A3z9K4M
+eUPZ6HwaeTbdqh9ymbFqxPWYrytaAXnFvQDfz7hFCou/gmnbNgBE+hh/mWj1vLRvMhXxy6peNKi
zNrI4pmp89ZUCvUG/LAlbnnyBsDcWPPa/aX6+DzvsFtavZZMyNgXpZJFxXnV2SBx9CwIuJA/OLQb
kxlBmghnM88s7xYPpZFVDa9ib9ZSp5oWL4PsAkwn54jPLnk5eruKwah0moODbqpnb/QpOXwRtSAP
9rkmM1W2z1M4IzvNjVzdEKv/D+h5wjOEkGKqHpJW6N92CPr5sqt20TOR3WlIIL8hejyvnFkNr+QI
5I3jEimjj7GuGqfnsXnNTLITQMPVoxAYeqvspUM/ffKfKQzYvI8RdXB93GKAVfXR4/WRRR0AfFE2
Ssfbf+Brx7SD6l4uVE+Mwn67npqfrVpk2bky9Di+mrq8ICXtcwbKBZeD7n0nAKeQjiJoUhAHjOa/
Cki+J9kIOohx799RUumUY/KJQHEGFAzoKb1u56oCwS+PbBo13TrOV4U3EOQUQlltlfId/U3G2k/X
/S4ZAguiNzxrikJ/lc298pqC87PAhrMVZrbAjEbahK4hE7fbMiwjzNPnw7PU6OzlT162xHhepj0T
hJVkU9JXOT5gzMkAnBTGblXkA6Og/WsWh6t+qi6zzEae25dI4xdEea2A5x2PylHg/d0JSnGgnQ9U
m5WbWC1T4SlgHpvUJYUq/iLRx20iU8/jc+j377lsBwGppCCzO8ygH5uxRIS3R3+6fethVMF4Yrbe
wXWeYnzLhZFSiZn8MTbs8rkDl8rpxEKyN65Ti2erNKdvHLu4XDtAwTkEND5QaXlSJuA4BZUOZ/Oj
fGL2WmDagzqy7erdlPr4gLuY3eoQvRslkJzosh+juqDln/kvhX95PwFocBSPUl8v1AX+VwKeyrSB
DYdWdaIxBKYhQrKsXoKpOecuFIRszsDt9S17qlFaBozBkVGlhX4C6COxeL2QuKFaOCegxJWOQVBM
h3P2VNCDE+tTXcMj41TQrJzz5Qx/6pyIoRPTZlO6dQsDAcML7ckUZK7h1lqBzBvGMLe2eSkFGBSf
PG4Rb8FoIxLrUX1oZGcoD9rYm406tY756l9deB2gAmUqZr8tU1BhvfX0qFA1ec0FrJqxn8vGzKex
0t+EQhTLHRenkRUy1IKpslGVKeaqWF3U1/6a6/aDHbakyMbG6DXQqquXs3c/Csu4rZW9+4B1vbSK
A/uz/dr8zDB7AYUmeHaKWM1JojNp3brM+JKoV+isjCU9fKV2GO7N5818Vze1WIbIj8WhOgWX9uwy
lxGtoqGWbUXiy3jJ0RG2/bXp4ClrPSVy20a9uznp34+Q3Pa+IbBYgvP2iasPKlaJTeBurXr8zV+f
kUj7GU4Ru1btcKDcBS9jE4mwF7v70oUdwMqMDgLSNRRwiYvQH184KpY5/yOrcmYOhUP4bzLe9/2r
v3Bc1fy9Gle/Ii9IfeAaviFQPUZX2LqX9Au9ZiEbXBejRlfBJtNuSvTs7URKLP9A4JjBgX++ALy5
jHXXyoFq2zSuGzcdmYZAfwHl4TEFXyD+jr8a7Mv099UvSojFJfQJjdrlrnekR8igc+5iplByhFVA
VbWb3ZP4rAAwVSxT2x3MD6+yM2ZdOEVWBVvfEowU96CyzCANDSw3OFnPn/DoSfjUuxarORmTvJxX
eFVAO9EVkLLDR9sY9MkF/3/MrY9VYNsUjFALFARX9Y/NmZDEGsGAZZ9HYa0c2MeJMeOMhbNQZ2Xu
Ol359yMrjJd7mKURx5iQMBtUwPT+SQ9yBTrK0C86o9m95sqOn+dkLTvIsTifKdZZ5qTYxNrZeqmO
/XbW/hMBF2zMo+5lE/gmQB19vOBllcOAu361icG1p7Q4cFv4lHA6ZOLWZ+7Ty4CXcgfTC2c95QOG
V8lYqwRnpiXBjt5bc60CN9mJC0Coxk5Rw746a1BwLpzMg/KqhF9Dq1TKxgcRZQKuowMoYrO1mWyD
hayeuw/UpAgPic3IEcAoTACpR0eTDUQ9Gs+mK9ojcKfcq1SluRiPnIyAMbGX1uqgTSqVu3EatWHv
m1HUMDDRdN6fl3+kdhYLZO5mq2U8JGAdsZaa2PKhQXBz+nnqKx/nWHbd1TPZa7BcIXtqxKwfsbOO
QcWyvsEHJp5zV1sSVz+zLj8ONVa/AK5qwqPvV0jVpAI7SDf1G7TtsH58hgU7U9Kd7KG8p04vczCn
mp1bppsCV2+/x9JoYtDcygICZpKMVlmrvd29mLLvto6U6Li5f+Y9Wrsrtkpdo+wNRL5sFOOZG4Zv
arsTwmOZ4AVQ8T1n9UV7kk5Iq1wu+TYsQuMt5RuhZQ0BwcIuvsmIeQVof1lV59RQOjpiv5a7lZ/M
Lh2HHHIoPqeyPE0OFM5CF9XobcpKyTFMs3UBgNNaDtLXKfT5TRFRQ4cDl0laay0DKdjiB9i+Zr7F
dmxPg7MmNhCRRVx6DXkVv4miv+iun0nkpIdsAUVn0R0pbgKFqXFf/GBVGQtA+V5sYezn3kcd3rku
vmL74rL+4ej/UxL4U8IdwCOau9Xf6sOZkN46je1mgYgfnHxKGMFK4rPAjS/6ETZo4r/1Fsrum4Y/
ICYsRLr9cL9ewqkuAnBjQ3ud3lw0qjeDjOgyRa2MLrlqvNl/R8jzXQjRXCWa/sdbRzMWIB7HbXQv
NiuYYVSeDBG+g/KmiEuy8XmjaqSD87IlW21Xm08D+fghjK37Hu+aZdSfXPUKoS/y5kUQSV7ahEwX
cLwGqDD1kUzjzoMSTEewqtW4LBkvwz+uFEX0kxNsPDTUEA7+GSmCWRZacaL51UA1trdR9HGnc7tK
WjIajXzN4FAmfm/N4kPNCzwFOh6zJ33+m6oL9Qd2syGLmnoHDyE7MInf2Rwq7qOpg9Q8qUuzY4Ao
ZHmhyt4tdE9NsOKNx0PxEmXQ6w+cVeCWNW2zHpTkBN82CDtaUezUrwhaUXVSLfyVL/cfLhvWuavJ
OGOan0rj2aq32JQrHlFmyw74QW7IJUavebdBEikWFqgoU8TL0JYqYTEaKsyOMKWgzJ1/KSr5Hd+4
rkTI+oFEyV9CxWVbZLAFZ/KzerleWnliBpk50tGbmZfrhoruF6DK/v/DX9DK0URmfPiuJkYwY1XE
VzH0t2Nsp8NsZIoBmdcpL/d7Ut9LpYuI66DAkOvo5SUKdhrI0wcBV4N/x4X8/6henDNQwsEto1Ry
0tGzLyZaMd98X8Rpbr7KVo1biH8a6VdOp9KP188f14I853E3em+MZxUYsP2qQXc25GahpLL4h9vO
xnxAjnO3hjJVLnKUu5B1TSqLBi7wsDLHjkiUgU6ztG8f/XtLa0gw8cKvSz9JoDoGdhRU4UAv4itN
vzCiVabOV54nXxcHWyHxPszeRYdz5OCTWGrgMN3PkJMgGh995iYtbpeQt64QnRsI78jDPdkGmNET
tkasK51b6ESkD/A7LNMeVIbRu0L/RTNjmCAaZarRq6EOu3TB8qL2u2/wxsUNLHGhpOBa39zNpyfO
DcYl7Ih5Ewsy/KwrFEv7Q1SSqrK5hEpdQnWe/L3yJmKYf1tS1UCELeBhclF77MWultrJzL7p5tDD
WFwKPvt01XlZxnw0ZvtNkfgzJG9Lm2mu499IS87JmFdZEmX9M9SMlYz3wuiIhxPFWvqdVrQGwrup
JEqaX5omt12Wmnk9wEe0+t3F7eUs+KhJ8sBijw6VMSW4/hAIKdzaOUDnSnO66tzY9Z7T2kiksmzX
iq2UuZPHnvN0WYIc6kFMT4TABVgBXhogWpcNmr1SPI+/cBZ+A/gC6Uu32AfYcyZEMhnaZhR8i7GV
g7c55Boj7xG4UlyGVHTuRhVU5AetwoynFDZBf9zHYpfwS+OlBkcq8hYx/gT48lBmYtiNuRBNnqKQ
ner20g4wgQyoEUwzSASr2AJzOpWzqDBAePLdVj9dmZ10tbs6Q4359KqS74zlbG4aI652P0hcBa4a
xAHCI/auoE8N5QfJ58+9WgvGIMw8GxUbO/Fc66hbplX8f6+jqcLWS33FECKUFyyrNQJRKlv/wfas
11fnY82NcxN5e4xKxF+ILkPzt2xjkybJJrwL/U7GfGu5Ms2OV8IdR2EG5n+rrtFElvp1cpoIcn1a
P1T2OnjPTm8NHI1IDp/zI13I/HyiQKY8hs+cySnJCluHv8cA43ihprOMTJgvrshvWV3a3gxBFuPs
kmAFNmaUI0TSjC3p6qB+xXm2kgB24jzJJMhgFJqQKXsZy/GIBXFhkVDK+fF+n2fcZIJEfz9z1Qlo
hMUyA31UkJfLCy271WDDTU9ahT6qKVALXBMEGir79QxpswUJlQ9HLOefJKG05/rw6Aw+ERgL7lcK
tl7lI2KT7xuKoj3p1YGH/Nu4QR4tYSNqS6AiPiaU7m7kLrOvU7DR23jRa6TDxWrajZUNA/5FNS7Y
xEgE8p9V4yBX9myQqKxotglXsGyMl0T87qcA69qg9UEcxR87ova1RDoNK7zDWd3sIkYLh1BaUYBL
3Kkw7iPiVFzz62Fcn27a1bsbaEu+CEtkjuhMo5UwocJQqONnuokP003qVqX6nSSRDCR3xqd/4vwq
7F8vL14U4EVovSJ+epHMxvBDp9AfT7WMTVMRFEJMv0TmczaAkb7x2Gry3lhSe2HGVbNxDWzPyqhG
90DSyTAO1ggkOpRFY3xflr6OUc0ny0Eb0SIB0YDWZJonWYwvSe2hz+RoFbkX9gPtIJvmmwSiZsnS
c5K+M2yvBdnByIW4sKgiJoIN0kozhunQJRGvHaXuFru3CXqto7exOkkjr9UMFWOdR3JoRq1kih/k
TSzjDpArXVdK6wz8frlVIT4OOVocrhCeAcCyMk2y9k9fUZcU5MPJ0YpIf3kqHih81tvg/LZ/L+9A
xgRbnqlL2XqgCuYpZJItsCKpduFF1r3v3+mHkl1lO798kuwqUgkxAp5AVQZ+M3Ais/T/GSyz2qMo
6hE8LU5AOjWFDkpP+2T6yiX8BsNT4HZ0tnEDiY9YZiz0itHjLCH4i14Erp7jTSG8lwUQtBFFtOmd
CMtfnF9fSHv4wwlJ9agSzFUF7DB/LewB259Lgcsb7E9qjBx4Ob5yPyFoRmgsSyDwrJxRHIo+LmL6
TG325PJvtvNdji76fKNz8yR+qLTKPwxelcJ8rzgXIy1wBlhelXXTssKsFDF//mpNjTSVK446pOxr
iVY268rwlbMLuWKZQCTf27AgJsKA5np8pUw4WHVmmqNu6iLo/zLDKk96M9gprHAkW9smzhFPnLr7
S6gmzENxBJrHLiZObX3WDjqoDxSiwb6MQLyXeqJcAVhVpOIdyUlJyy9A6ob8WQQy4l6ZLAUKc3IH
ApjXsTnRiJMdPQdquWac3fkzmIri1hfwlXD6gXHoGC9mk7bhLeMk4y21Mzu8G9pkArHgV+JYoLF6
0krkMfeEE2gopHZ76zOmZgQQaFjup0YXFz/T3n1BwDyMxVv2KEt8VbrHbvp+SlypdVrvAxikvXX7
y7pGXo9PszPNgAQ7lDxwl7XtBtENYIuw7zUyWC91Y4cn1dQoMgflS7qYr96IFDMx02x/cg7ut230
XzUTSRcDlfEj3rnymsbm927jFFp8Ft+ogVhOlmtZCbxKAfkUVAXgmMrS6BzyuZpdlR2Qk8Unh6Cr
enrGkWU8l4nllluhXtljU5+4IX3q/3NV/uIzknlXnQZHzuP8KadskLSooZo2ZYwoCDz8jGDRtQXT
7AIlY6NAz26KDJyH5j80sMS596VNNpRSe5MLasZ74H60rWdtszkDD6XD7biSQ/U9L13NCVgkTEQI
NR174uGH1ryi3YFO3fG3XgCuIbtkX+xy4MYV8goeGbkIpZ4EF5ePcTbgWQdmnWeqZ/vId2f+BNIp
WOiS84HspuHMGp21FSoOqYYoQmd/ZBum3O35XhyCnqmHPaTRB+hOuE6YB6cwQ/XKIUQ93lxW7U94
5Lwiog0Bdm+5opGghpZa0oPIL0xulv/05rNuC+Oh8xxlwLkTR0YCZ7SOJ7f5Xr0K9iKgl31T3b5U
mvXhLgY0KlsTf3N0e2sUS+29hwMBgfOmQA0ydk7dnSNYAvc5URw7ncNZi59rbvTgNhGpZlEeUSkb
cnEsQj+ICfBngvR8HHhx6DyZRKaBkz0s4+sfB3mLmwXSoepJY5+VSHX4D9eKyQ44EInLEtCZhRcB
bESR7IwIz+Ub2Bku66ZaM5DQ7vt9NbeYkayWdulDuJrVVmvpIXFLoz37LXvygSjdFzayzeM44sBU
CJVS5R75O1PevzXM1mheday73W7zH/0bRb5pPvRSUAhtkUxOnIRUrFFZAaUwooqZOMUIlTOcP1nc
b4sVaJumsm1BDbD0BGgFmpvycyXiqUul2TA4XDEXWtAWuu5kzAIoQQ+uOJugXaNutbvvbtvHsZ69
vClYhNmgAego9AtT3BUf5w7keONWWxOvrMZba7OVtdJTwlVqWzT3oPRi6ZuFlQpFU3wD2Jbi6ITU
6Dtw5BsgsAHWpm9VyR1/KRYo038RKAWJBvTJgVarOAh9di5wUwytF2oMjiZXgDe14XJqgOi+QvvM
DmGYsU6wTR26SxfvMNb6f1TTppJDtN7Z2TYK/VU8tdyYBiNP253NKeS3Lk2V9twEx5h0pVrNzflE
f2n1WYHae0hIqzP0p/DyITX3SYIjqoX+118zHLM1ywTafdzr1lBp0zy0diglA6QbT4KFqooXWRNX
nb3mWViIhGU0ZHBT8bMkU3KsKnlOIeb7rszcQbd0fpzGbktxyb7x/mg6AXRO/XceQbRMY2Ldg/FU
EzKAX5/r7+FdD6BrDgLkuKWjKeP2RS1GBqpe/1PW9aCstx6ntdzRDNTQCvOeL4aHRsMaApPPR2nq
4K8KBT7r5xJ7kFQkuYh4lUS6/5y/0P6L1U30QInjs4o6tHH1O7SHVlsflhGKOL8KRCvrh9EtULdO
AvuRzT7KuOX2Gg3nZ0uQ66lx95aJHiePzp8A7LgeYkhcIa35+8ZgcgnQLIYeOGhOEkhqCNldV9AJ
i73D5boOQBKW7GNPEKYFNmZRJIuFaApE7ajMoawJ5XTnwRZaL+mggM+X4L9CM/B8FB+ckk6He/JZ
sCd4RalL9nnsjibijchMGsryDF8BHLWZmVj8EMMzJEcrg9A4PXf06SQ9Abnby7IfQEPw9sSQhd+I
W67qpWsnkM+ooouByFtwdswdA+q6JRy1gAX+ent4MR3fkXWU7n+99SyOjcFaq41H2QKT++LHsxSp
W0mwgq/BqMaBrHq30kmc2EulYQXaVbOWha2xUohL9WAZ9/PiTX6h8E/v617R7i0wg5ifEjNJg82o
Ubh3IIN1zVK40t6NRnW2yISri3pz7UR4ivR7Ozfo7RK2KUUzV+Ayh744udHkkfy+n7gonBRJgRdd
OKadQ+GyEwUb150teI3LiUFva/UJqrPCuAH59qVAujgw83lv+igFpbw0qbrMJprbD7tu60A//RDn
KPDKNaQF0/B9uslzoQM05QKnx1ohbddJQnXzYJgp+IvfKZh75UVOUqLJoEO+XiVAaQpQL8eOBfGJ
p7glo5AYf9IAkd+h7nA6h7md4JWOdTbBdjnIqDc8/d3Nf9wiFYr7zkF/6zoEzk5zhmhezXAceEJb
fizCfHOrd1vDAA8NVNIN/aryKrqxwUr0eXW3ticcsR3PlwsXAJ6FxrubPpRHusJJburz/Z4ucqR9
rmLg4DTXRXvrDHNXRWYdBjoJtqhi+5k/awqlMK9H0v6x0g/Xssoa5Y/9Gqjk9OBQrtroZ47Pe2Ln
R0gldUnpd3qXTrftsOO5qb0Cxog5R9LJiXzgB6eUYyTNnexrz0R3vgWWwZ9EYkC4vpZll+xFVQBH
5mHIPAEm7MANnOUL0u5OHEsfowlmLvnqj9WAi1iRYO7v9Teb7xqXSdKHC4aDThjlwnyke4q5DDyL
35o/Z6OuM7FT5Suv+H3MAuuCUDNzP/lDGL63moI0jiydYhG799CYSGQl4XlI7f/Xb4RjAgz1mYCb
YGuOVmoGOKCgevPudibaEgXTeF+kGJhowFW1gErZYu7FRBO/MlHe3zCeMbZO+Q9zoqCGwZy+6qAx
/QAo/bjp9idwEZw8m4CLJ2J0Wy0gvYylIVwSp+voB8E5On/K05zQvLrKSeTydBzwNCR/J8IaTUXo
scbixwsjEkwtGwLnMzuU+3DFdvH3vsQrIC8g0XpyY+TjDjEJp3EftRqCWc7nri3sR01+1PXjq5GR
+bSJp3OjGVmBNdU17DOHm5ecJhTcHwIO7RWv6kEhk+bq5L5Ir74+D4KuHr7wUcjC4aAmKhOHJu2o
8bLOec+KRcgfYKXj0W1wOxGfrn1/g4ET3Y71yukJS4TknQkKDZQazYx045XVPu+18uJvoNo/1+Yd
7u1F8LHuCzBt3HFE1ctjQ38/kzakxIGRlQ/LaIobMJBgtB/dGX7a5Yyb/65Za77WptnBaY+EKzQI
SdWCkMolS7uUS+aUdDlr/Zp119VeApL6IFVHYJb13GxDdUtkVAY5Tk28A24trfZq29myKLLNMS+q
l+XTlyMvjlGLttD3yGYmVy3cplrRHF9qZAXm1SqipzdxlmtlAg4B1gniVzOPdtljGR5pyhslDBPj
qqKRCcTBEjk75dqmmxeVNZC1dITzcQyGlEOYGQQxKW8ZwzDL6wJLrW25idJeBC9oe5jvq1kwTqmW
woKlKqDE9bltAK5+1eEslbvWI2s1UXx41WilXC37U/71C7WD1sFjeXEfDkRHiMu/wwxDqTxgdvAL
hXCGNFVSiopm2uu/6rh26qmgcVKnj+168J+xayuKfxUm60d1e0hV24YUScAq3dbnJ9wMQO9BPKwn
cX5cKbFl8+qbkSLXgHzSEk8K0S2LJTVan5L734ZqtqweHO/alM/Uz1qqVb3nHPi60QVsPdrL5D8s
WJJVTM//1wZTdbo/fLQAoC0fUHRXu/+PuvC03gDP4Sho8x6iI6a11VykfuhugJO62+pwp6nzYOe3
wWSSVXZjlbWddlSn5bPXQcPrxg9jxWvpDuL0F3UixgTkNyaqbCfumbe/0wK369LrbJNG3MfEcWCU
cf1WQb9sL+cJt+rQMgZh3SgAxa4DE5uO4Bd0YEphKJBngiwSKGs5/kXOaifn9DXt6I4tfMXrbh0J
OoYekBducxelkHFcp25nc81jlGU/L9bkbMrEkm+U5g/iL9n8FVys4ASf3RXr4qJw4mp7Lqw6a255
Vyh1pSytxjyV0JYDJ4u5UlumthM4704e4QMJWWQRUp8F4Qx/MadNyee/oB3lOHXP3uCMJIZgGJn/
+Ldgv8nax8zyBkfuuOzvENLe9A/TIXjmxL+/hOymeRxhbUjnoh1xjRDDiIvCVtZFFI0UBhSnPxXn
NLm3SRFpl0pEqpA0AoW3L/+yaidxdiyJKuLqs/YZ5MaZJI1JQeo1clmesyZiYbgl6OumY9WMOCsO
jaFTN1sPNuvHsBZ07W5SaaRs3qXfKnHzr4kqC9whsVUK6DLowdggujfjKTq00U8ro7jdeZsKZMSM
pSHfnsWFqu4c8ca5g9F+9ZIa1grilTNyjzIua3mJ21IahBogvAO4qhIg9lb4lkfGAYmg/fzHFxEU
xYM2v/SJjFcdr3aLYJ1KreLCQzRr79plb6GFjOzJnIrAl41fKoMjrWZB0EJAlhFpAREClyZ0bNF+
00m5htNOU1eGp6Wx0Kr6fBPh6qVoL1WH51U+aMrr+lXa30pQYu1/FmRPdGVArLM8GBkpcjshwaV+
jX1gXrj+5z40ABYqxQ6s0Aec3aoSzwguwO6lfENREzLx2erD8UCLetaUJBMRxlRWKRhzfv38u5sh
IRJVOqz6q4YXJz5lKIRKXF8YT60Mn46B+xgSC2k4hNwBgpK41kI9+JxdzSHFft11/IKNTQMBx0aU
f6C4r2sbpyttais0CWjmZJgd8O8oQ6GqnHdC/j8OIO371b7IQnTIILaJUQ9NsEM7qfphn9Ef1R1L
hm9AOL2Do97s9SaeedkR5lS29EBmnuKHvd7DPIGG9EVtFyLOr7xyypuRmyLTER7QMeKbx5rCEYFj
0FnGz7Znoi8xfjlojmBZlJIYe8+/AlldL16IJVBlI6MSC3QQ59Svi2fOc9hSbI9poKX9g6Wxx6sU
/FtkplJN0vjpMoRs8o9d7CWMXoqEBWvu15Eg2IP6hfc5QW/qmPqkgtAW9rculsLcrcALbQxql324
/5bLw9rLTzRf7+0wlohdRVJzpy+Mu4IXvFcBlfV4detikOY15yXsQ8G1filc7dVEp4DuErWOQIZ6
ktq+DDqcM06WvG1ckj7YF4P6QnTtCY6UjmY/QUKIcp2mpG2ySsUrwu1YoWqL6etIIO/RLztc3HqE
sSrbUkebE+uUayWQPkNX5hVuul5sWLo12grBWzg6h8MNX3ONWZRKAbRsdR+MLZhzaz+uZwMBLgPk
lRPJW2r/UyeOvgEHAsBXRaPWcDPQ/5yRhZwHLru6d19Q1v4bTb7wr+jxx3x/m8ewSOxwfo34Z3+k
h2yfTBoPKh2Rain2GsQrXB1upHSzSCjOqiiWiEX3CCEUIaYrEUvOqoXwNjhPP/qBsQ2M2kKSJrZJ
ffLXkQn7X07bwC4cf2K766BtMoMEq//T5G0j5aKoDOVfBdGLQtPTkNNOxZcpx4hMrBvL0j28Db8g
nwT5RDm3OhC8LI7uwOzyOAputMwf7IgWr7rE8G7O3d6YbT5i8hUfup9DVGBQVttoh5XFwembilfN
GRNCzoQMBbOkjetP6EHxT0zlLm85YWeTteHVh2AI7WaT5lvd9XU/DcruoYGAIqZPRW6L2blkNEG/
LZA36SeZa46QABAW53o3hcv7HDWttcuFg8LVNbDv6LFZLWekMx/Zr5WsP8+Dry2MFd0eTVlb2n5e
nCpJMwuONBxgHuzHCPUf6vYD1NcvzsdtHKRXAqDmYJX1a/06yL8k+jyBUi+AQacjFqmE+ATcY1/Q
RZEpAH7rgVMne8LINQIjqGovl2IVy3vPNhziNroxpbiOSo4d6UjiiePGnKR5RGcUsiEA5fa4dw58
0AGk1xzco+FuIF8UxIC59yeW5+RTG7q6yQwXxe+UHKkZ9yOdxD6/xiWJBJGuWgIMCZCqQeX+2m0G
iMH5OW6Joo2d4Mob/ud111+f0KIVKr3GLf7e4tkRA9g2bvNQ79VB5MRuRfwed+jWHPwXNnHw629B
YZmttotaBbhRfO5Pf5S7ZBG8/gjHH6yw4LzBSbpPq76T6ibZjgM1NljC6BNhhFoI+YfYffsT2Ecs
JOqeNPc8FmoWhoh5TXxTOArM8iv+mgrkwEMkIjoQZkWM0jPWAlyG5kbx7hXG+7zDjoAyNc1liVRe
n7R9gARttv07RsD6HbKhYm/E4P0ExxOaMYm+OS6irK8WDcqgwOGICrY8CLw6RS280B7yFLogXewm
g75SC0bP9ZnyoMwGTeXzZ9TQBjrgxFybGpM6TDnJRssgjNWTS/k/ujFxS/n3BTZwQXH5ngvqnNnA
chHpEwi25nn4WkO2i+SGH6DoWpoce0DqVzHKcZhipSPXBvaIQrof7u+7PZMOvJgtpRXQXnTNjUZ1
1MD4ys6QoASdP0cmno9gVM8dtsuvsGxz8vXpGBYE2b1taWnk5WADCiJxbr2VehlskgvIULhrC0bi
nOYa9KxzCJaDOcB5YhmxpPDiPC0COqWRBOG1udRL5GBFdAB8gOgBRMRoV6oZDZkfZyivQEAQwhLs
CU1lLR+2abKeoepSHH/9N3fcRO/7nrvQnH8Ym8J90twr2j3HEaZOiXgvll1NYga8PNd/f3trw5Cw
tZ3lgkps4R7fy/3CiD+IoeMfFEyrS0LyQXPleB2t/LK3q8ha3R1e/g3SvXc44MQJZob2o7PQDLBV
MeMm6Hmz8NtIZz5yY4AKsVAMGar49/905X9WpwiKnjzI7oBo9jEHW6lWSDc0z45YL1YrHic58mZD
uJOBE+kX/LNspUNdSSo82jHPdTlG82LupuKvXw1oLZaae5IEcmYymQ+fSRRNH3Z5J4lqzwCiywjc
9DkIegAtdta17xlfwJq2O/TwkudpFmgy3lz04PpdIFAKvx0UjIsRODhd8H0Y1YC0BoFq4JfVPqaW
iu99FUhl9V5xTLIIdifnxqTxvDdim3yN7wvXSv0tmdT2Hv4GzN55XUtV9wWHMZAs0sXwY+WPOrWn
LuRE5DJavvxS0AwTnmrPhZ2g6Ko+Epoyq3Rr2rKsQeH43dDLHi7x4x6VpNSRzdhqU8xWmGXbrE6P
lc8UkdQCqOOxpDLDdLmgPUenW3g2yi/Ez0zgj5K79IrWFqCUeXDQmUPL1aZurINmUHusNi1f0qPV
ykV416wc/+8C5k7L0iq/mk+BVHrGISdrWO/oGaS9++LcdrN791UHY/tbuuveGpTz7gNrgR+3wo5g
TFQRGNRVUCFxY/PVv2zYtotDC7MG2PyWVewxd8y9aApme/hArl6tawyxsbsgK8BeawZIy0hslZjk
99T9H9m7PF8aji97QOnejtTXUPG/5hNx7uap5Oj+fWhFd/7D1CUVbVsRtPjPxQSoXC2uBQWsOzvc
VOb6pArveO6OgFEctUWeqjcvrp2PkXPEKBxU9xM2r0YgpaD3nXUhn54ca02+tOyL2YyTMseqv6dy
9mWEPdOSTr9wFEVFxFSEklfOVL0StxZ2Uj/s1NALkNjmrQVKpHNZ2aPJaUxzFwnmjmBDTqExZly1
Kqqf9QPZq3xQTISxPHVfgn+5WOtAdCJ1c+SF/5g/ujpp9BpJdsfRolowS/KzkoKGiwFXm/Mx46/E
knv2iVVllxIQb6Q19/s92CWB22WriCGLq0Pyw570tiNruRRjP9GYGi8OkpR6u+tRzaRdQp/vLzcJ
qzykvhMGP9Iu41udshkLUUa0Sdc/IrdBVsen/+nucVHIfOdndvgQEVruWaLDdRpFaNmCo6AiCvOE
PVP/QpIDhKDKj/pEm1tS1MLJVS/z+xLWbaw0UPOSOFwvpqsSzRTU5C5fb8i0WDAjrmS/v+VaUOI+
oJlNrWQQlXVHiq1gx6fHGKayvIWt3hJTiiSqz5ONMTxPjyOb78URdEvmWSypafXYBVhxlE56OHQf
wh6HA0QRmaGiBNap77coxxtPNEkCcdzvdb0vdOtTyt1kJcMevTSTmfH001g9TrexnDff8SShKC1y
LyxmRuEN6HVrKls/mVVuR77DMHJgduZ7nwMxb54dDn974A7SIR+s11a5knF/rCm9+IqsB3n/4y+T
3BkqYy6PmvgTZ1jmE3wiBgqNuhVqpwz7JHPv7wzwa9Fds0wzURRqPnHBXZ63JAB0D+o+7p9dRMVb
Mw/Acejb/CEzMjD8DjcUeXNCHU7r+3ygVGUN1a71bVHJ84z3GNj5gdbxSNpK5AYt/DwWkMbGcjmz
iAN63a3Y0mfErnLbd95UldOhNeUXg1nBF0PJVnN2YjAjxYLKxu4CiL6DKww8pUY5Ihg5yeo6nco0
VjIRBm/BOYUZ02H5CMv6OQhtRQ06IlzpuFbO3k+q+iRGcSZFGsSVz54upiieB1nhIddwHji+di9w
niqgyIzfWzYtKgcnTTmrcCxv/BCfqsPY6GQOaQhYqU7m5H/RmO9DrDDAmrObFDRdgBxycBBVDqXQ
wZfvaJuN705JJWvYZI3fvCxlAO49+K6wmPcQVecFuSxQnTndVw5gqrBCw/OYpYt//g0n884Kv/Oi
pN53gNsgd835JaXr7pFUswj7HaeFeGc2YqbrwYeaoQc0/Va1issFFqXwts/Kgrt6cS7mIyCPmx86
nurZlmxXqDtia/BxjTzXg6JCQfBu5hhgcHzvuGO1lpiRbIIIcaQc6CFVQa+1XMRfCrqC6pMItqNs
/FGUF8R47e6tpbulZ+crJ7IrWQDtY63MPmfPRSqQiBPFqof86QPgUQndypGq9u+vp1kplvE0hhQP
qOuKrt+HWtgIq502ZaTrvJUFelG3RMyz4xEBLXOpcOgjXXl5fN9UgFR9P7M5LoSuQDs2/3tARhpT
q5sHLWGikvr1yy8RB2awMeB2mrRUhAo27ky+7zmgboeBNG3QgVyGp5Zcl47FdVgVpFrV+1Ai5cXx
68SLYdfeGTtCq+aLPtjxaEiYRtrhpkFp+jVmT2hPSeyHGtKcChRUHuHsLtiQeuDhDp7aYNf2k2g0
UmEBD3J2x91CQrmm7oiabVjbIuBawzJQKNPkOX3P363jxb2YDWNDR8zYOjOBxWwJRUqFE8CBDRj4
qzcr8MeDqX4t6AAv5hWhVRKpkCpP7x6Ri4ja/yESscwwJauXDyKQpdGGkcoDfSnXd5E40FNoYArX
q1+G/bR4HvMBmzmtWC3RIYDFZ/cexcGnyO57BMmbBUBhb/H6WcJD2O7XiaPrAgDtnvuF20nbUll/
Tq0/7kbeCzY3Jdu5yP0MDpqlxwJ6T8jOu9nM4XPKe21PnUS/Kt7Wn/1Shygk4rbXIiceVR9z9fIA
XH5KZkzOSa2fIo8qNauW7NTj5Y8darUB1ksFadRUi8Mv7zoqTXWEQhYWXPff41sa1L1lf7lnzG1B
6/IUAQF2DVF2PUaq8si6b4hq9XvNA5DxlRYBJpOSiryeY1+Wq1pRCFwMlid9Jh/KHRnNJ4uzlo4Q
wOfWkwdARY9wOeP2e9gPzH/ghkR/pu8+7Vv6fMryJH8HgNgUZM/28sbv5SDyocWkLej1jS8eF3o3
voV1j8c0/Q6a6DftiUNvbFq3hyA6VTd1uhlDpsuifQnz6szCJ4OXJ5sFcHXoZswxF0Op0R8ZRzgg
yr6+u8ne/x/RUG3CcWmWLQqPHHGhb54fmU5i+fI6vWQHVVa5aHZ1GgFy3zTeUSNC+vexYwD9lOtF
j1bVWx8Hc2K2cMMnCIz5s12zuFLW3fPv3MzE20vzmNdDRyCaew6/p33vIgcenMRZDC7j7gHXKnl8
QxhngRA8lOAT9Uu8NQmlYIkdUUZlPTyiX8CW8MH3LTbXX1HwJELBIq0XlYVEtl1N+duAFOnJKRHU
WGIX4RYVvYJZMauGn1/4xDXAShWfwvDBpOSVOTlHuHdvjKLeSV3ylBRSR+Mbrt8R1dH0PknpQWN7
ucCnyxkNSf9OeT4yOSfeN5Vn+5x3jAvgOEmG6IBPBdTOLKRLLfBcRanEK4oQTOtJRMBlYGs48Qdo
vnuvc++hGpInKeTsRw80Dxoql3YX5+S39Mw3/RaD0vM4iVA8C0QcCun8MWkZpr1wjk9yNKB1ouJZ
mWkY00Lb/pnui0+JIXbv5vjNGZAeB6anptNSI7Utz9Gx6zhDiMZSOf9venAd+67zPrcm61mIQS5R
qRDwrYK4lTCUV4X4lM3sC8ZDZMTdZeLoCO/lPbibkyr/E6nYCg5XQTTIkQU6pGc519SGkMKaNxEs
PbWBjkrFvlNm7DDHQZVnxIWTft3vRffjLOxBQLxsA03brqohYfMh6OO2lO2400U6T5A9sP4HU6u/
7uyMjbmNjz0JrpW+GlztK4U95qDE+13w9/Rqnds/xlKy/I28dy6mzZnfBfna5U8b+JC5vnHU6hbI
/C9vK5XRAJ+z9O0nN7Q3t5SvERiiHRqXSjPsMSYcizSUJO5z68Q3n7313UhavZJX0fNAc3tqMB+K
thAUXro75DiS5mwAlOKyHpk9bh8lGsHqouPDHJlhvbnQ+y8Y8RJetPi5P5iLWeIDoxVQGgD/9I5n
qsasxBjgtZEnvxkgtOvwBj56638Oa4Eh5ty8xb9Xe1/Q7ElpLepqz6AEdjPnfLMjAWl1YXIh7/tR
Nq2xG+8jzg2kJ1LVFmY4YgtS7xbYjDoSI0tijFgu64emD/Ibx+98XOQ0y9BJEQCxiru2fE00ueIF
m8aT7T9jr6S3bbmpPCyOYSbWXzDmAW4SRz5+Qdki9eNwp8v9A/16yn07NX2TxkxiewmnMP1BODzp
we+4PGmxISvGDTexXDmpXO6SjGR5a9ojt4izpqcyJ2r7UCIDz0d37AmhwvXN/whLX1bqv029WZsh
AqBEzR/4T5vOShB+Gn//SPduJkqG+HiR08PaOA8aI+DldDnJ+A+7f3dj23DD+B3sD7Qpkpi18eBC
Anz0ymMbsEGjYxjRDpzQgHgxkTHHPm3+iM4fBLTND5rvPYldJreNLuWb0ViRegGbh90f0nOqH3cD
z/ZytjsvEmp0j4tsAKPEIyAu6s94ZVeGdm2eEK5ZWxHv3fBl/Un27E72QTW41U6aiAfhRJ9eW7Iz
xAXUbEnK7b2XtOasFdhCnJ1IJjW2AKw/9+TNBxJ5WOZkiTTc06uymXOSUp8iD6clehuPbMtEl3M8
5ytTAdt7VqNrQ4oj0jzGY4pTT191GsmaTyiTusd2wfvYBUkE6dI434mmgZePRwBAR1RzY5wFhwPl
AYRx1J5PmhqFsF1xv2CI0M5T3lZRBIjR2TBT5b4yGbXfUiCTy/H9xo2g4rkvxR6hTk8Fv/miWliS
PMWXpPu5MTvpc4mxkSpE5eIHeGhCIxZZsRnZ3Cq8lELwVNksxOdafMObnpgmXkkHXlSCkmUIJWAs
U2Pyi/P0yj7cCQY0EuFp9kM29KHxEFS1ydPizLT5/GoyVm7PIoOcYb4NtX0UzVtqy4/6qc2gsJxG
dZerh6e8k/JAZbbL2Bb2D8V+PMonTvo6iCJgdYc2L56DDoKbM8tuVAAL+rFl6wBAGjmCkh025mVI
/+0kKiJHytkVC482YzpBYoOlvwihdVkyt6mjxqcf1ZcrDqkiqDzS+kEY4JmpKi6YlL7jO299Fk3V
x+K2q+bU0IRG5Hoh5KbUGr6AEd6YIsfUXkQKzYji/YC21ozE8hqXBllaBGjYYefXuCRoMSSlJyWk
kSUsTVUkNf2Xzv026J9Q5mKWZk1/bTafZM6riaYrtyZskNYCVcYrTBhqYNUpnANJjPy2gB0w9BcY
Fi2IyFtOs3btdfXVvWksOBOqCUlIrqX/tIpWQM0UoEBAHJEwb91ogIy3Jf2WVq+kdQbdPkxkNlJb
EFzAF150myEdKdhcvXhKv4iI0e7liJfrwtAGEn0jnxWfCp4Rrsklly6fXlNB2dk+Y7Vr1QwmAQf6
bxW2ZJ9Q1UE+XQcLyUlIJOyRR98Jo2NUpmPRMysBB9p876ie6SXcLQEe8rR/N7D4OUW52VDhOH8s
s5Jd71G5XCHsCfnKV9TKwlN1lHzc7Tb9Mi4FAazbaiKxuBySjsRLL5Kh8povzNYAizZG1HPfH2YV
fsV88GLkAY6p007Jo/Uj5EqlkmDs47lwcnix+zkGvuLp5Mv4RmD69l4WLlxgznxYB8awXC6yxScO
RzPe/n1vzpnuhr0UtdKskdwPXH5meiQcWN9cwzzo5i1nHvWyP33jN25oCIiILU5OM+sdyKUAXLZ7
CY5wQNj+qfBpXuB6eB7csp3kZ7x394qvrtQj6OzLwtE9hZHSsAGunTrlc2LE31S8ULAhoBmjf19v
2xvLnDN1Aw/qAMd75wEFge6nlEyWGBZ80jXI3xnErGGUgEI2NwjRoY1HdRuREoT4yb2eLEqiLOZD
m7V5NK+Z8soC85UqMjmU9zxhI9ZKgawhVtJ59lD+pL5PonOhACI5agBpt7IcuUCsFQKDGFlbLHsU
WO9l3Cd3qHWmvJNzzoNg27Ggn7zk4Q16f4ZMLRBZXt5tqjT/wgi4qew9M36DxRtIaXW/txvZZy8W
DsBT/vTsZubDsBnLN+gfqO5E4mDFNfrWHBsCgGzn/PtScFT070JSNuL0Ze8NULXe9rTPi8b/cuUP
Dv+jMp/lJLSokhDVGqz4n6gsIGD5GirEyj3/kWFDC7hY8hP+bCjplxmAZg6R0UqlU3HptcQYGcSI
OguiwLxuurWxj+LhvC6qg83ukO5IJLI62RHKXHBpwCHkQlZqYGZgnOF+3alArxCaDlfTaxxIfplb
jBUGHWt+hnm5Tk6U/BS0FTUsFbCw7NwvmLVyYDQg1MQPoY2NTQO3/rCbc6piFGHbDoYmJjD12Egm
NM6OvuD/GmEBPC8k9cJEVNK3MQQ1hqrFmiDJ4kHXVoBLAQwWi9LNRza16XPLT1nqzSZsmZewcUMr
yXXk0xWb7FTfMbFx4Bli2Esikp2p/oFjE/4E4llF5Uu2Cl7Ny4PtRuGKSawHxGfFozBYJFiV69Xa
QJ/NcAXXX3w3eIdcGmmn/tgAXhHco+1mJVrSnl4CdayG3GrTG6suhEefNXS468DB7/sKDu4C8YfA
5LAkHV99OV5E5pQUlllwnyWF2KzoTvXBPe7tgiwsIqxMusAYzpv3KO+UGSYTWOd9e03VD2fV9/m1
fbUpnjKpXlBiszC00Xe/39cgajXQizsPhSHsUJKafrfhp326KZreWW3GxHpRh+RkaQrA7OymGPyC
R1fJon9WW8cfH9ppu1L5hhqRadKrlPDzAynJX3jWoydF5mTbVeHa8cZnMoHWdeLsC43184ZkorjD
NLFzo/GhIEhl7vYCBJ64EFOzIpvUgW4zxBW1FNAjFGcM2fS1VoPoeWf4cixqDJxns2TOYCGrHo1L
yvypGespPQo13m1/jJ2zUNE1Paqep1MYp+zLdHXyRIWkBvT0tcjjVjFAhY2Gn98Nhel71YT2jZ7y
NLeg4J74Uq53eLxYlPnY58zG2Ez1o/c0UdpA6XfGMEBU5/1FygnXBb24GWe626g2kImu3Au6JRM2
krQM1Qvmy6E2Z96Vo9uOTDglWzImOALio8q4ppTxXVBblV7QFBupmEE8LsCPnrN/K7GbvMflgW3E
R1mMldihbSOhIqpIp4VNPfXk5WPRDTEEv1iBFDcEQJosK9Z2vd6vP4qyX4O+7wsDeSIMLcMw06YI
MYlUpdPcduYYA7Gdu39O5Q7+kGTZEecaQCNPyEGCNryyhMWgPj6eM4DD/9lsaxMgxxPFKbEoORfM
bLunuAFko71rjOK4aB6ZV1W+U7PiKgIdRjAsc+nU368D11K6fT5gh7s6AGWc9Rzr2jiWeWHHSDZB
mQlHMtSX7d1jNpCZu6g0z1y2vatdV58bZ8mGBsAq554bZ0VfeYAQIhg3rJrZtl3NJye41fMvuiMA
VKRsL/s30rGdt0A/H8qNAojJaxCdPDFfhEFzQIsk214bWJy+SFkf2nHOAnmy1VaXM8srm9oUvAWl
7f+SmgIkQO52lUOaxFZrufCKJ3x+E3trJf1dtNF8EnAyxhysy7cyd9b53Vv9HWTyrZgZgQI2lz3y
2+FcHN8h65TCW7bXb6Qe4OI+t94uMNDVH6nDwrn2w6vD57jLNXzSVnEDstfGWoLe1fk4vZcJEjXx
g5u6IH1d1ItiAAM2uLwc9vuAIkZzUnJawkwm0AbBlr4YvnF6+CuUypAuD3ohW9sRUAOM6i676avD
bXh8tyYQIrDhWt54cZOB5TDQMraIq0w+eAodGd6Ok5pmLbsj6U3VVafDvtOEefVsFf3xj4uzd/V9
gFAwqwMR4YySq85OVdho8jjwotO8Z3a0fqI4i4SK9VgiOqMYklCPgbLyLUJGbbc6ZdhVX6+E8KzY
Iole9M+x5DZFtr3xrBedDK98P7qitUwFlEgLWQwwQyj0yMoKQQnXKshIVHFDT7JR+36xU9cFNFP7
GOzCwDfn17T1dHlpslW8MFv4/YXOigMKJ3kPb0aNfcESuZ75va4JgwfJ3hiATH8Q2XnoopA1F43b
G6+1QiLofEIfF2ci8zNe+uUrFDXOS2xUgK8yN0mzFSQwnZA5KUCb2WDc2aF53jZW8sWFgowxoKSP
q2ZRRBpY89503h6RIGFgb+OrX+IzaehW3gMUA3Q3xfnb9Ui77zXgXM6Uyow2otmk1RK4+Qv12N6l
wliYEV9Qqq+PVdZ0SOnOZswoMF6ZHeK4XpEXQS2ULJwfAlozQmWZqeH8GysekhsjRCJjfbe4dh9T
qF/p3Yyr68cfIPwu0qBec+dq+zUok/wkWEwtBKwy8eTXAueB4UOsUaLDv+rpRjtRXknr+w+/mqUK
YFtreA/TkZUgBcSlUwABh6ce1Jk1kZmAa5QaFoEhw/P+fyMocNQGXJj55T+V7WSOKDaV/eURI6+x
dwqyY6FTMPuY7lzH2u0wgMZoAoHJXMOvKPw9TjSIAaB2ZRn2aOmolCtCLrsfx0FvqpFLNWQN/zhb
JLLgpZYVP7hHdXZxYic4nWsbki411awdHyew4b50A9Z8sFy5+FPo4fl7EL2ImjcbWclMmKObeFGT
rXB3VgRwD3VW8V5gnjSj/WZkpu5KZJAuY4oU6X4RMr0yr6tNkZdIthtKAw5o1uQdX9EII8ZnX+/g
Ae309lXQTNGwfo9jNZVr09zdmtSYdd3w3r6WhrkiJptMwD9slOfRcG8xLy2c/ULuU3Vsj+jei/3u
crq8eNyHUWSJhikUaUOGzD68XPdIyPSFfC7X9kpTHEzSqrzNRemDfFQrNt/a/adXBdusgJwoH2rJ
kOloZn2ExmmwOiksPK+FYoArhbHFbN0jh58GL45S0W/bf04wvpcsqENVpP4b/gaDd2mQGZQIDJbK
5pI+bJVUQODimVIOZzKyYVy43duiosU8EDn/TLKHACaZZMBOerF5xNmX99XD34A8RwZTcMy19+HR
SLkgxrYX1iI2tjCFFecilr3/5GAq62OVWt0QBYhIUDNwstecZNaIWmJGUMaFCnYO892JMDBbt+we
5gQsvEVfXI5hNT6tnYkBE7DoICONMKR6ilOfzo4raJH4mf4JtQC1cLmeCZH6WxIrlbpYZmFN4E5K
Jr9/KR16uHEDmWf8cf+rcdABVo1Y5Ht4fsX+HYExhO7tZjihvwnkcOmXZOUACxXVWHXxtrpcbDYB
4SliMvVUujkcriS/nEsmje6Wvnu+fUpk+71FqoPBFk7tiynPIVJwW9kLRUMvlE6vfPys1Ac8QdjK
ahxKzSUOKnqdCnuDmDE6lpQ30+5Z/mV48mVMLUyIWyBKgmvuLu/iSO7GtoJS3Ep9ilTGqgvQvY/i
SZMdn/5IUlfWl0BCRG/CkIryap09L65EfpKBSEhp6ZW1aqUMUG/HC0ChLfHhhQdX2xvNm7y6Y8GH
i0NtqXvbUaUSYe6VIZXoBvEevnumTaI7xT4H2oB3ERg1R6DCgzV/snw510zNfg//KpDWNK6GcCFl
bCGInkTXNJAnGTWUGir+/iG0tN5EXad8d8EoZk1jPEcNAIAAzJDlYANyeFSvQkHYMGG+mMru0RzX
9sLD0m8AxQpDj8AqUIs3ylYwz7cdbpGze83Q31g+Me8E0S0JkxrpZPsOd29XTU74vYxVpbFa3Hdl
lKsfE0Vk51MSfsUwBRTVldvOvbhRKYlj+RkTwHGUh7nirapejWh5KOhpvReNtGbWz3OU6vUipb7M
I+TxDlMEBM3P42D3xzOVvlxU21vJKp232BzwzWSKa7IPsESV7l0lkHW1CqD+P5+wmCJVRNmEdJyx
Dv7Jb2+1BBUCwtXI9ulWqCSdfhRYD7jOcKTd/Xug/OVlv/6fyEKI4Be79NiZ7K3KYlXiqXSJXXf6
G/9QBvNQp4CPd6fS/je3j4hTWzow/A+R5aT7g19SL3AEJTmvSlZXWxH2zTYwyZ30Tu/Q5cndtlgX
p/9CbMQwLWTtAI/pFuBW5WfMEZYk6kJ+wksM1+GkzSPu7zK76xYWakp8FKMpd322LBAQCLCXikxI
kHrsj9Lk9KFvXUlZ2geTz7TwnLxF2XuK5r1nOoT7MmAce1yIgJm/+348hWQNsUAbbzijgeddE8Wv
k1tIhcRK4t5HHzl3uZfd7RpXOutcyooNopGLVaAQfXaLKgeL+L+e7coGeMxb90f12VZ+4tFMi6rJ
xyV+UMmCkzNCVwkUS2ab1nSH+XlJVavPdNKPXDHCnyTLwJzar4/lsXymBwKIehsVcVm3xGhIJmds
gwelVkgkByW9n274Ibainjltq0oYjt4uoB6YQVRTjX/NysAiXlZi8VE3y8S4K+L1Mv9GDeeYwIKW
TJfKAQRIR+oWSaFShMmDoCiZChYOtMSZZFWMk6OZZx7Gj3ifLcO+1Sr0zPeENeXOddj2haoH6aK+
bnfe7Nvll08ZurFJxTfUF200w7TDtEOaKLhX412QnMe3++EO2jxEyfe0yqlBZl8ZpQMsKTZ1Hpt9
rnSdroxdFVKTKJZkvqGalx1GUxwGCDNmLXfa68qZpBD/u37khgg4JqdJBUnPQHxXvCM5xD/yySRX
zp8aAYPf+2Sewft6jTFU2DuJYUUkHFI4+cozfXqfpM1sJJdPGoySUXKWCpDMF6evv10kAXbbYpVu
2Ob6StGg0iZnXWjStZVljI61MTv2qujuTdJJ8HwPNy+DjdZldSNVbbvnRi3hcWfPwPlXtGCavSkj
PCSvtWT4/CqZfTLPeY/hcf8EhWVqgHfW4gnSFWefJdkTLMxHIfIUYJIqKIZeUPlHTEZlbQLAG7SG
v+dDP7SeNsBDiq4Kbpg9ngEA4JTWYu9Bu9LJ1B0g2atDg/hVSDOP8ac3aCh03Mf2egj744qxSOiS
1kB3YtGTKZrZYqIEHu0uE69Dk8IXAAnO2kLXVlKE8sE8Zl+4dVItn3XZpB/PCexEmqqDFANcArFL
xaiS4Ijri92PONn9SJweAZABJkNEbMpyY9hHuNKetOzrhg1X1wgIoiyy+Uluv7t3TN3FRaf9YMcU
xp78ffzp2JjNHCzBy8gE1SqG/AFgM2AfHx2EyBq4/O/VwNWRkEzeEY4ynW6D0EbvMlvcgBuLNVes
ojs4z64IiwoNfDfh8KWQdVeHGZ7IMWbXLsuPB1gGoeRf2uslCuMnrlsFltITJSzqY9Rwtw2zPNXI
dJQkEvKjEMklYBBZhHxOo0B9xQfouSXagUUyJOeyjZrgQmzCDjnrueKfq/aLnBKtInX7zVKwdEyH
TM8cv3/ORU0pp1ZXrEMF21V+3Otw6CHemfLsfi+MAPIpR8cPHBbl5vda7MAyvhF9Zwq8WO4uXg5Z
05V6KJN63U0AJQ+7MIKMfIy0MYDg3I1EDdl1Dko53hFvmazhbrmcXawqVUQyjzzKhqEgLTBK7FIZ
Zbiesn8eSxMSm52kByBLcHwPKTo7CvJjRhTdoZqi9eJM/AaCzfvqkEusR2xhnA9gF6wJbhNunrxa
9F0OpX2vMyXYkE+uqVMipOP7XmVR66LpHQFye5/IB5+exi/V97clhYJBf7xWDmO0f1QZEAXb9+mp
ZX/vcj6Uu3HwAkhaVsACUkhVmmVP3U7crICU/BOUD8QceuIX9topANH6RPgs1xJzd2e49ENQqXcn
1616E/fbPQo5Hwsz1oD9GHuE3JhJcVHcuLUfTGgUH0TqQ5EgO0Nc+hWJXhEChe3TcwdkT9x+H670
3a82sFK2B+9UBEh5FlxE5hi3BbhfuAztOkTR7iBSW2msEeRvzje3CMiyTPC7qVWTMvTEaU6ii6C7
FT9hrNOEQWm8S2O0asxYtaSi7fmHSaiXPVXCibKS0HxE+rRTIChi8Kb0gfOHGXsF8XZt/xfprSDy
QYc35S5kXNWlt5nPfiYUDjuC7mZVsbj2G3rWoToxEr6zzfkpXPit1DkiOkpDnj+7BSsMuQO9oujj
mx1t8KHL2pqGccpnA5C86HANQSvC/vcwq+6fJOuBedqyYLeAsUMltnizpHsy4GkKLXbtgwZbV66Z
JcneU7TVzsZU2I93dUrvZZfz9BuIyBPrw5N2qZ8tb5QFSDZPKgFQAycmeuN7Sql84jM+69ypv9nD
ulFWMpusu7eFJnvOkL9vCEG1I3kllRXefj9FQdE3U/I0jK8hnKXNtXsQ9NXe3AdtNbpN8+YnoZCP
/RVt0JJ+m9A/Xcn0htjFSAGLorSL6Tb9POobHGd3OmjhcvduprjXQABuUmGTyoE6UTmzMnAKk/rM
SXrULxiu1Di2TR/aySppeQ9Y1R1rWbtX2gXQN/Y5th4CdFhnG4iXEH/4fGGpLsUJhGL901cvKAy6
nMj9Gs94ent6p2uPen8Q10n9aoERWHfgFgva9fGNQHy3LPsZVcQpU43/1yIU81DkayavqsgTpVDm
PZXxC71y91tXNHvV+nvZhW4QKNEzeUexqM0q3bsE9w3ioxLCzFooEHCfxdUXodp/pOSNp6N12yL9
vwNZG1JaxhIBVppWl/Mv9gDMYxSZ77oNh1TlLiw/MxoeWMFq8ujsvHa7/jeyZTx1MJtGERGlCSTs
3ikozrZmkYE3O/QtvlGe/b7T7oAYtXQi+ABQNmH7UKn+7BxwMFhlFLXFwlKJrOx62gQbfV6CYue4
rggft3JTP9r8VxrMOIxQXGnkehJdu06UcFgig5FpiLi0YF1UCnt8ZLBrvN0nuegtNfgedS4fbChz
zwmn2JoDPUN4ljSXa1y+o5x93IgHVyF886D/+aNmMWJSlj6VHpPZVdWYZp0mPJxm3lWkyDByUKgn
/PBYxqdxBwIboT7TJfzwzkOF/78uWYDqVSnpNQHc3CPMsqkfHnG7nxGYHMoriuSjPSdRaAPDV+6v
3ZsED574uTYJlk9Gwq6iePyhH4OXTZ/KIS9DFAJljdfOQIeorhBlIETQypESU84SkAs4MFWElJj/
w6c2fIzkTkJe5/VvjxWfVeMskgvfx+A5Bdrnq+PCps0Je2Ubw8SU9dxFJCS0HQrN4rbiYJ42Tbv4
hYGfScQYcaaGahhH8zeS616f8RR9sAqXYtKwjHfxiVrnYQ5rsG6XFe6U58T5rhuzlXUi/2tkNFEx
DcC/r+bjkytj7niHQMSVEVIsqG3xaICpRllq/GYZobcEQSvAf8KI52Zmvy0p0KpBhuTyj8KGYo22
jbsJl2YZmo7PPKfsODdhLC1oF41h29fxOCZYXwM8iaIBCWu6Diro/gXWOrzvr6m+WEr2J1qAwxVT
LEyJDzZ1mDmZjzAmG7Q7JShFhiiQd+vmrXO11O9iDav1EhjY3BIVMXtDM9eymW5OSYsEpu7G9tbc
G2uS0sF8BeAk0+u8gg8hySYQ/xzhpKNvfzSQQkban1uSQiLH2bWEo3NtOlxqlaGTS9c68NBhua/Z
Ug+VZYOR28Hf4ryWK3Kr/UlQDjU4iRw6FGdl7bSQzNVysDVhj0R6oG44Za/aDu2YYFRnlxhfIalM
ErICHRI7xmWSX2bx+WyexHnYxh3BwQaPTHU/oRI08wX33EKLGhx4WQsQ4gLe4yVIo1pZPTcRKLVQ
Xd486aAaunOf040oZuQh3yh9mYXEyx/Y2qw8aUS09peWTSxQxhilGLzhzRVqs7MGq2F5QcqEYck1
/tDqd5TuogzetV/0Y8reGq2wOK38zbpqIz+FKcfYCl2LPiYFMq1G6euJPYWU+2ZnfGiFPxKGx7fL
VQJlJaTynLHl8aWFpOZuarmZKtyoBimdtxeQrUj1w4jTKp01KzYau3KZOnkYdYgAZaGM2XRO2+cO
mKk3FiCZ87kuc2+qXAsueVLFdHIcFDVVpPNld7U8D4sudbHucu7TtMfOerh+UQKj4XAcIsbnDO+q
cQGQ0wbmBqgb36lzIiRsqMWyRSgaoe/Suzat47maX44jR5HnQFslTFKLNUx6tlkO3FyIJolX0JOI
CswFNty5R4JmsBDE7STO+0KAKwzrjTHk35yUuKU1xrnUkF6HDSIFH4LGCKnS4Oo1N46QFL4kl9ir
ifMW1mc2NoSfOSdOtTLi/BpznNSwxS6IPOzClm8hlXQSRqvy/RfhO/lHUsPvK1fJAC6oSMz66ZGa
GeT+h82kXhTwN55KzGsx4eXTuXlIpZi4vHXu8BhNnjfCLjtTMGozj6BWOgRvNdiBeY+BmoJn3Vys
96G95F87kPEvQIJ3mEPwsKe51eaSobI3irY8RYGZ3VopAFEn95EjxODO+6pPatGv/34HLDw6PkFy
GdLdjKDzx5ddUPAenh7Mmi+tZDZMYob6EtiPBkElg+2KNX6+hnKYXGWNBxmLO0vJBZ7KxCDz4qpK
58IDTvkeC5kKJV4MNQYZZ2R87c74q95SP8CYlwEt2A+dDaEChNsU+3rdumB9J6UBhcKE9XPs3Gw3
+8sElpnlfPqKrckt7nuL7ma9VSy0gxA84R6DlC6LY13mFhintNUqLxWkNZVEx+rlnV6Cl/C+d/aZ
RKkd5MeReHQxSN2KtI8JrQ0EY+GQ485C0vLl8bRt4tnudSMEZtVmdK8KiTQIAAirnTXRdYVfo1g3
qiOYncNgwdQe1SxjYKq1hQmt1YZG7TVSnQ7AEQ0AEVLkLRcrMzyCNneHwAWxSFUPoNQVIVscbI9a
scikAwhvBI2UnkXIry2Lpmvw627/7ZI/4UORll7FuQpTQx98Z6RzJKoLHIpWJi/44Oi76bT71fCW
8pGYT60YWsZqZ1xAaWp/lB+6tRIZ6AdA+uR8VE/RerDT+A2Z2Cy38gpBcGRpwfruwhOBi2CGuFwB
l4L4lzEv5ot70kwkfzFqOn1c67QceALLgq+ASbEVD8O5JrRiLCFF5OLhrX+upHjAx3gQM25pnaII
gYmr6krV2jhkdUFQLBfEEu58J5gV9cKUed58B0rCVywnDZ4xIPzOop3M0P79DlJo5GGJvS6ys2q4
1hwfhbsXWAQ+iBIRRt0y8DtneBf7szWovQ2QmsUveuPO8PhJZZJzaCvZ6k+Ig8icWA10egTckZ4r
wcmc8pD3ucJydpjSOP6NCBRzuyaq6j03T+MJOseM9Z0rRPIedhNP3HMpRy2a9sziKcHdelzea2Rj
QgftQd0rtM6qygQgysua0Omo678ga5h+g8vyakDhlobnZQ0k5svkcaR7Or3R8av8MPNqkGnrWgjX
oKBX3sd2lb4ux+b27QChg3SY30Wp9TYlcs5VvIITCEVQo/qALpZ4kJla2E7APUEbayb6vupqARNf
O8QWAuzkRIl57gDmYBWNdwdTYki/+W2g0wlkg7LMASNrByFR3lhjtjj/lcrKM2hjcUdLSitcLZl4
3TDYUFPjib0/ievwWekGYuKJplDLuwxebnzGbyd3HvksSuQMM3UM28JZnyeU6bGGb+f0Ozqei456
YdNMEA039tMFbrKcRsBR3T86djQ56BSn8gg/phapUg8v0zLz478i4uAm6lPUsWzhHziLwOAJyUkq
cMoJQ5yDazClPuzt2CGfUq1G5y46B/6Lh/nAJIL7X9J1nFguyJ+3zEQNpThjb+4sJL+h9404NMJt
Rw1/6QB+WMV4eTERNsEWtuEKdS2kR/pExsf8vxG68IXazU1Jflx53fv1CBqwuKxb35wHmpxaN3wV
8qISpq82alVTv58ul4DLlSA/KiWT266AHDWsvNv1fyyjhG79TA97k+r5eD4skv85dj/qG1mdJM4U
jkkGgTFu8tet+d2KocBX2IhyoXbOCMt0LcW9VAVVGWJG7RtmjNz+XC8VYNM/BsGM13upOMi9Wfe4
wsJPBaYyvMkba3dJCOG7rahen/gb2/71XzrXXaEbLqNo81w9TTOTH5XI7+NCIeDGd4sIA/KSZXuH
G6Zc7to3PfYQ7iJeGPMiPb/PRkSA092F5FKN2/fcSQl8tA1FCo4ZmNmSB+P+X2OOcJGVGs9AMJFX
B5FoF31+JIeJhvQrFVe4jOw+iqYmbEc7OBgO4ABkrhC656XeP2tIQVDHbBTIH6UJ6Uz4SsuFOrL9
pgzIV8NLlYSPK7jcqVCJy1Qs7bGgYuCQcnEp9H6AoRUnQJ8BlcSViaocOA2gnxDzn+IdyBOSArSK
kaC/OhJQ4sO1boDewELNShppgkwuvchGjbuGccgKn9R9XwMRl66CvbRIBSq1dE5zY1iiNKbyIR87
IHl1NczpYrV2w9UXZMYRhTl6wUGYBBPPo9XOlu+M1qvt6aBzmZVcFBh7nwg3tMSRvG1+Ehv9D4w4
Hmga0s4DE1jmkkbFkGvTyOWBRmfO4mGT9VmHjxzG/N/WsdJkLNszBjxfoWcx8r27eItNLFqWtTsT
dHsCB9V2iznFLRN9BdrET8kn9Y0XIPc0Oa2MZ1k5trGwRi746nYHpNwHEhQpDgKBzn+GjEcbDxIH
lR1VyGvffvDw1+MVrXi7UnPIAjuG8jkVFH9iitqhpq2gZItBW5yXlky4ykobWLnmpgt6HCFarQSV
40I6gqIbOFKiOy1xAaHyNb2c9ZqkWAucdB40cJrPjK5RY/i5zuolZQ3eJL6aQI3bMRX9TSJpBnnN
FJpdKJtr9iIgzr8PQZGxulN99XalTKwac7n22hE9tUC7V6eb0wn/ozmDHu72M51nzA4JkhRUMhzb
ocO0reQC2kmf0loeJSZFM7rXvHb56F2jwAu/vNVdWNKandUs+DjhkkGtZc4mFBm92EmMTKv/tAUi
b8sXDe36ejoO1oI1lcIKLQPcTCvhUY39YRFfA3J1X8b9MSdkXdJTlBGrFpDkEbHHVTvY0hfTWB/c
7YuhTQ2P775hBL67WHABThKmtTGHQYFmOkNJmlaz5OHJ7K1qeVan5oCKFplwD6AWvLFl0IJSrPBU
Zlbqbaw97WS/MHoX8tGIvIJiPMZ+LAkA8yPtAsHs+CNuzDzOy8B/LkP6pjtyRxPC4JeaHaBOJpQ3
EHTrQ7vC6OPMCP5ZOTNEcAvSK4zC5fJTIptyJPPAVt8GgYjxGeAWsYnQfivbDQTLNxgs/E+vIEXR
SCVqGZUc+kxE0aJJ448tS1JonL3X/LvuH8ACQLmhg50EVjohxOVMBsxY9REmtVJdIIWHmRjasnnL
Cno9F8YmvYzoRiWUfLOKEd7ybkOOyJzwE1XKXKfpkyxJ7IpPP/G8si9vJWnG/a10Qq7COHGN549z
YNyHwpcGHzrV3m67JPpWaERtgTfHBb32B/jqBUSbH4vPQjtXKc33LWrJPhy1NcbuknUlECMOXICa
4TY/JwG5ez1ZuSVmIqT6uHHLF2Mu3mldtPU1M4+eJWj5ZFNu0AoSq2nzajmbfoLLFBXj2Gimm6S/
aUwYymIJYoY468/6F6c+zkq5rJgQzDBtc0vOEicRZfqhyepHYKTzCHpZGDB9ccM1K2e880D23O1A
TjXiX4czMvtwfaFLj/Tgl6aMh5BKLJGH/gbfc1ZUr9ymBKYmt8ql4HktWd5UMkRrSCqUN6pV5nVo
vuSzHLsm/PxCOLZGahSCQPxpfEkXTCXRDltZ0J1HMi0PgUIwfnJJTvJfmjwmmzKWCLFG2y/cZ4MA
pAHFNx8YsEuZL8ZxBJeV/OXHC2F5UY0cYCg3ODVkDaRjEJZIJPWpPbxD6uuLXuAh5jUeCfJ6CObR
WRD8LwTsOGZ28w2WBNy1BnJHtxhceFuJ3QsUoh2Uh0bhYGQ75H3jZ3PbxUShpPfFbmww5IZiwKDl
GC35zsVt2g0UOnHBuAXUoZ5Jqa34qVsw3dh07+dYVw1acvQbt22mPoCp9FJetEAvv+NsSo/O+Udz
/CRI2cI73VZhOPHloRUO1ozQVvVuTPCLVsMWCViEogo0aFvNiRjaa+d8dIk+YnrZNWV6YxuFQdCW
QpYcW20OmJFu/Sq+T52WRJpcjdMjvRtYv+aMdUb9en7a4jGqun0zYmya/xr1HMXpLV5mluqK3CMF
hnify21rOlLT3dgaSXWLd4xgxWjyvYdG4VxO7Evv7qWDX7bb0iyP1nOJKDOlwl8Pk5kZgn/6Bg+V
Cy0uALzOK0wYS6+hg4//7BTQtquhg694qhO2JgjP5NjIrl4TrMtCqAmrCEla/hhDEQG02LZIQmRh
52UwEDYMMYdhoPPb2KBRgz1EiTTbYEDjOX0OpI1pxrSAQm7Ex92EBX4qYrHni4k8m9RJvWggqA7T
dRHwtZQQPy0vfudT/fPGOOB9Sj6dJgpih+9pjlzupkGWpQyXI7ukfgs6865ukCRKoLfv/HbSZ0Ar
d3KTUOOYhqfKLd5fpidMdZjVs7kvO73VL7jZaLtpA1xykygbbHxNOuDobDBoSHoYHi+8jygATpfd
AXPHrOe5Fsr+IpxI+SRFCq/4A4onJi0JJ0In4r7HRs3uVSVBrrPuUkppgnyFL0irQQ8NUxdG0hn6
voro9Mb7Qo9C04RenXnfD5a4QaHRkM7OMZgM3zI2ojcCNYxVz0HfuiVraGuY0PCRQy7XG3RAODYf
0WDxMizwMDlHglKgGpk6Dp80wpIo2ayZKcESDNqcGwKsFnubb4UjLBXVUKRglCF4FsVSPsp3YU5Z
gjkIyjthV1qgD3aLVPUAammwpXTsICsBKB4rURks/kjlHBNR6ckP4hLL5kgtSiRpDtqdVC2qU1ex
LxHQqYEJutmteEu8R6K0ICYStwVxUMkkIp76AU6uYLIp9UaZ/nKj93YKaEGZ5mFpj3NDMV6/gqLt
hPei0+3j6ebaWAk52I6gVlkSelcD20nXPuk5uOs60vjxDD9CVgEoGUl/MEsvG5dgbl2JZRioL0D+
bYhzpF74ZMcWQC+3f6UcOg69hZwoxqERBpNn4J0YGDoJAMZsBm2omEEfGsAJLeAsGmQRrss3ROzU
Ufy7R7bijvbjwr+f/LNk/XeJu7zkCZsfH5XTZ6ZZIV2WY4pF154xpy2aQQfReZiA/3GqqtCKabtX
V1heUFF7Qczdh0J1KW/LWxKJhK6yvHddoDXZYn+Jo5j9nuVZ85uz8tNOxo/XJ/BEFRtj4N4lJpSY
UAis+EFptH87fSV1xnae0egHkg141jT/3SoNrzdnBuU7wAZNrktRDJkidjLTmA1E4WaR49So//tl
zr8fj/pcO6Dpz8i6x7HOpDCarV9yL5S+XX2kULvL+Au/3ywvlJeHYeh+6yfHi1fN5zPWS+SuwRl/
eIMI3sbcFmU3VtVwzwyUlrvbpVSL1WUsLDR0iYSTLKT/zHXD7NCzxNOEOQJaiwxE/66f46OVUTnx
0jQO32gdePaMXDGOfNYxRb4jkEMTWbqUhpqIENYRBDqRHJIrEoU4ljMa6XUEakatIhbqFE9l3wet
o3eyKrTYjT0gnY4+6TUyh0bukZ9ZU5BsCztAqApj+gJ/HmCA+x6R3uSu5/UyO9ZDbq8ayQz19l4y
dwSIX0XTVSyGeMRns896lHGMJsotOIFIkpkwTPqabqDZnhwjJAlkV0M8CmBhp0pkvGs28kuLa/xP
qXYRKa7FaRROCcF8CFDm6zUGQjhD37RuMmgZ3kbnhY1Dc91qmcFsuoTZwBOHDeBhp+ao6VOOsz9I
jHMQsFrBZW7dphg9uHQkHzt+RQb/9azbiqU8FVGuUFgwhNgpMe0Qd4vk4BW87uI0f6gxT6wPPbIu
QvEe5hPoH+cqzAp47YMkMSJmqmrgIf2D3yeo8V05DtkHoZqwgFRrcJM6Y6L7u/0g3B32ktvnYKLa
2tVsWbQFTBWIGBsx0uaJ9+RWjrbA4xVHH3UIxDcwe6jihsZAZEcN7vjbSdG/nIzM1qiMpT87dOxD
7ykiEZFFnly1qEAyW4PbrDbJow0lobjnpgSIpz7V/sQfMJuHbeHU3Z0tJ/wuAdSynETrn4XIZtl4
fs5MehqWFl6uB0mG4RGHESY/5aiI9iTS8Tu4MO9HFnyFxlV+B31Q+Q3mzOew6w9sLFLwJx/kQpeS
IsdSWWjXMOyjnvvy2dzMA1euaQKTy/VJuu+zXWJ1X0qHXU7VfUdBlNlpCuqXXud5G8QdZ5vtXvYi
FQTbltu7huK7sa2SWjC00S3OGzUrv+mp2BC6HSwAmHScqVF+GJnPkhPPw8jqUTud+Dx45jL8FP/Q
ebf7Z1FFs/I8maw93OiRwgxwtJDKHmPZbMi6NTCVWl9SHsbwhqkReCpW7i/oeM1MjVuXm/wCs5sx
01k9hqWHVxLdS5WHXcCFHjaB10TPbmrA5qNnwAxLrHj32hNbXK0uDjo+1IpYD1XGo+k2OiP4uiUo
JcyeDJDsUZPsVWXLgKnC03qZyYEwv+6ATjm1dcaFym6AK28+CT9MacZx+vzCsC4n0DCBiYCnFQl1
F4C7DzbKqi/vMIvWlRh59WzRK3U9qz1DKY2q5oB/wQ+05Oq6SlxFVpPiUBmmkAgDgrHa0Qg0dJaj
nyFh6AMka+OQBnVtrdO8ALqmRsRn+eYxfUlXlVehzZtszv6VqQFGhZs4E+trQwq2i81VUl9is0F+
ixagxCUSxeWKqA8r9ogxZhUAWse7JxzfsMJ5BuXC3zUfHLX/AxKrWt5RtznaY7y8jbUtL3zI3xjX
qm7QfpyhWV64BP/gq6O9Pdt2XG4PY/ZOeHbck0P2yjnkbqwKpjVVFT0RBB4zbpEeTgqVQarzsp6K
dT/ZZrXW6/wHaOhnQgD1RAYcmnqJX71vew4g0rt5OxQLwU87OUvtn7tSRYwin2SzyYhx62TalrCo
nTdmHNlwMJ8tZQ6whYYQ1OEwsuBcaqA05iSNZYhEBzR9hp14wV0lL2TS21qTfUh1ggFVXW6EFTB8
N861BwR5cF28H2yUqWNhGkXqoVEYfhTskbhv0c6tRa2oMdOi4vU/+LDyfy71KLy+FXxytmqoF5v1
Gj7FqDDnx6pjUuFtSAqi0fsdfl/dt4M2v2gDDQTrkl5TvvJmu4hAbqRQ7WRH4xuKp/AqzSj0P2Xm
Z7LnyXifRvDOTJudafdaii2ZGcqgJkOG7Mc3nixD3SMdn1E04ldwhDXkFA8RQnBCWALGB0b6VEb3
HawbkgtkZwX9NtOMrBw5xTrjxO1LAQ7/tgdxbCcYQuv0M17uQr2400s8GiPhOaWL9HQRbetRWiNi
8UAaWU51eoiZboGIo18iQ3JzhkBSUsZOLmq456zBTlvi9i7A4bOgtd1iNLPy83NN5TFPd2uAoMPr
iOUvVQtFbhbIJo00EpMkoGOXQsUljbFgOnuO2kg87z5ZS9FMQsWs8kFXXJwIzf/l4PPTgwGZ0XRJ
dSSEzA8+LrzdoR+F4YT9XqeUbyb/BfnI9psI4Z8JSrGM7TN+kl9BPKHRoIElSGknmvUDwT4Ms1LS
+J2zEY0H9g1+tMNAaciliW391os4+Z0aZ8n+b7RXgYjD8TkA4DJXVXQr9aPCBbP5Q4T60v8sKaLT
fNY5jPrb/3l5t70ubgeABQAVuCMa/N0/s0456tgW70THMNLnX38PnoMYVPl1p1e8UpT1w9MrSjlY
UHht5wPtvvnosgmjj6cU+AFUmFx8Fa16+dKJqWMUvYlTRBHYjDANZnlA+Cwz+8g4knYh7ux+nhNF
3wFmQX/Mnfd2MBhhrltlP988PpZfmVnqSrZ0nJh4ubnnua39mXNjlBvVHVh1hYMMdA20iUWAILHo
4suF3vVv2WPRXGTUJhda5C91F4zA3ApzS1CWmGglgeT5ctdOWeoafoCYVpXs2oskqnV3yPdhPcrJ
kU0y7BE7Bu1NcZYJ54LipQxElck200aZHIl6uzZo+3g1jpS/UNFyJdRQHdSdyRKg0H713rzlf5NV
N2Fk3yJZWJRSH1l8EUyc0jUgxmXC5YtXFhLGGjNer+Q5oX44jbiFqg0V9RNjX/cGdWSTIVEy9Fb8
Pza8Ge6fpW13W0TwpxnjPwAmLfF3UCq1kKxLZthOfwo/EuKr4qmyg8KY+KK34b8L54fSDj1GRQSB
zjg1JTuvH5jYUFY7yYYHoNhiRufD1ho42oQ66ZPDKuDO/FFMsmA7efr91i81+QoNLphlaTNRh4lV
eM6vO+o+xl68kFf1MZgDrDNYAMk9MAy6MJWwvK302YZwFrUrH8+DPKSbZegj/hU02v6IY2o8xBEi
qSJiFlrkRxZDeciTESFuhr6DC/ehGdpGYTPmc9aeQYRkP5/Us86hz4ya4wJLfvm60nkcAjatDMxu
qeDlSvfEZseV+0e7CXpWkzzl7d+Uv+a5b0frI/JiSgHxhRLdhW8Rli3l0Wl1ri4P3jdfI1dHbeAx
Kk5ZGeAz3cvbgYEO9eF0wixKMu8SGYIkNbEKxEsscK6lc/v+tj/NQXFR8SQH3k/LQ4PUF6h3O3KN
4bW//e66iaSdEzqOB5qXilK0WZ82agRhcp43rAcLbapbV96j/oE1tQBSTx6wIg+81nO9g1wrG415
pTalCkWpI5bkNfpL6JwdPJ6RHBZm2EyDli+y+TdlyNMcwxp++Wh9D15pkcHh3arg0jb/hfp5HZDR
0W0r9oHUAUibK9abjbtCHD8xe0Gsa04We1r91WAk0R2OjES/naaEjchOE3BYdY1Jp0VtZVv5/gRR
DWHCgrkk1AkCzBL2aU+KlMMRP73NEOGyQGl8DxsJWsIHWUIRaiWVTahM4eI4wA+U+jMSz+9RtN3Q
YOYThC1vj5XpkSgFrwIjJw5di9zeUi1gfPmFyVeozVLzkYEHJjU7SmX0i0bFf87I57ggrmuxy5+U
j4r2lfGrzMsz7MlHRwzeGUUmx2yPrz1htz0rwuLsasaIkpsig09RiNZZHr5rMi4YipclvBr7iSq7
Gu7Om0W8ZDlQ/2la1glZqMnRDYRTjW2jqT1HCMlkF5IIHGrJl17ptUZC07gnjjlnSL0gbxYnzsmc
xtKxK8SwZ2iya80CCyPP8xG+Z3wSI9N+KepIPcX3876g21+1bDWqcToAd4IGf4WvEDwdroSyPjMi
8aC2vsGlUxCfI/8aSHfAv6H2yiuj/ucfBWrUx3iyIZJKpQJbRjFWEhbA+wxTbwMSNykNcJrJmgN9
FQPcnKhIpuMjtneBoOJV1q6kT3jZXFRktgsO+XakM02OP29b/jO9xEA+8hLGn55B67GPAvdC2XeX
tVKmlX8w3BqCrBa7D+oUtq5pKgkLZtOmMm9rBEWO7+Xrnns2+w2EW6UWsTI/MjYY/nJedxnAhA7t
6yZCUG1zzYj6GrTUF1n78T93Q/9kG0w8S2MPTPMUDwTbR+m0ozI2XVC+G/3Siq+64j8NaQafwVgC
Upb09wiL221cHDyk8F6dS9+5fMMpxqMZXgy1O3sRhoWbqqh+va1PQgvTfIdXMzlizaxo+s4FvpN9
UO1BcJm7eMzgXS5KAbIwQMsmgK7nJGlHlafrefuETgZwtYZhMEME3o+hmw5uknKZjquO9IY47BWN
MWiL5E2mVZjm4GC8q82fMkU08cyo3qRdfbX6GASHDI05jtRI+gRwqsPazB6BHQt3VHh8PVseu4n6
ZmNZO6Racp3zKSorX5Zjr3iaylmjAEVtk/NKMsfF93mSLXH4sBGbwtZVD39cRPHFbi4SR9iayTf6
QWK+/nAIqzkJMdIIUyzw9Q81IROaooy5tqNufIHWdUzpZWMUzCVTlLK5eSFHewKaWcZ7fiZvV3xw
nlPo3qRxq/nyOQ19axe2bL/XPXfTkCuD43gxXVZPI4NkuDNIG35JySE7DFOvgfxnaIMcq4AFrjeq
1BZifm3ecSUvs6i9AnIaMXCTm4q49X8JrnXJEYo0K47tUhiAMQ1y7gBlbtxtkHGB6vvyHg6fKmdM
0l+WNGSnHfvDcM7W1r4LuoCMtm+PAuGZRoifFhazFo68+LY0LNnbGhvl8A3b7meS3XITv5nbP7Ea
8LWL2s/FsaBQCMbtZWiBVDXhNhUwnHgtZWEN3MPGMEwXGNRGIopmSuDyM6XgLo6dYqa0KzxymBxh
RdhBQ9HY1aLsppm8QIm2o9om/C/M3wNFsjGJ88FZGImxlddjSbxT9MOnQEv4bee3nTjnCInRMFWj
S/VAjX3vdaiuHMkg+1zjbCMCJKSlxodmk8ahLUXkZpN5jP3w67cKhv7QX6DCkyy6OlLncqn3Qj83
Q2MdPCjBrviwFs+MGG5vUImxzEfiYkqU69iidAeYQrDm97EgCaU6dzgOM15Gav5p+1iDFigMKru9
NrNXJ7NVa7lWAa+djhL77vnt1lCWjhGEN3LoeBDOlOebx/B4nH/hPlol+WSA/8HhZhAYB3Q2NeYo
ssAe3Akn2tly7Vb1RZCslyVmpQ+xsvGo49ZH3ziSSyUw6ObqohR78LcLdfAruvEAYfb9dpj2kiJ4
KKXX71F2qSi3FLi1G2AllXjTzvqebZim9Ed73+XBawgL++B/Ypdsn7d5Z+CyFiIohMRTBPlw9S/u
UMXMCvz1SBdgd4x81VE8Cr07HHlaGQw3jtLxo24ntzJ2D7CcyZyeEZzRWdXLvKee3y/BHLhKiFYh
R5N/Ps9EC+uwAUTTZxaSdEGdAGAfrtStAOnM4hYbxj5p3xrQx2jWV9db5hm/0+bexL/JbZH7nbTX
DiESVHLFj+MN+hvTCO0S9r/nMIq4hty5BMT4IsHh8mmFwCNR80DC8uTh+rACfgLNbZDF2gUJNhMt
K7FAVuxy6tQDFhAzBDemgCBKJTatfILTdD96DW9rM7aVrG2xgjnABUcfzPSrMtzDEXX3vGxc94tQ
aYuXhfZDdazvzZnqKyosuPsew8P/MyMl4egPCQ6dlp62mFtDwPv6Tzr6dBEteNHlV/8+i1wC+SNQ
LwZncLRXeny+fJ0VkIZBG+xZ+L6eocpkzD67Rufe9nG9xq7+ofGtP6K65HJ51FRZQDpRrTeKVtWk
Hz3pJHGiJw4A5gzQ/v1O+kHQe12rPwoTFAqJCLRpKKxMAGzYRqoN11+ABpO/lB+PJSfUr55NH8+Y
A0wXJvxgUhmIQu8OQLDnBJ4HKt9NO3KOm0883R/OFmXMhND9MEaqXD560Nvv6X2XGKCdTcI771Aq
YA2Ww/2xAlNzVhYj5DMOyH3BluSIGC/Ft2AGgbGLY3kNpPe9E7f2G64ab2sWlSEFhFJfetvK9uTS
k0pm/FPGNP48vI442lV3boYbyBbgpGSpBADozbu14ovLym39l2niKSvFnzB6xJqIafnBIku2I5Ze
jcYdSpJYkQTwijHYhiPP361i+2ocmB1E2eoGDjxd7pFWQ9iZ/AswPDAwyIiKqv9WHdTgXGYKSdvr
OzeI+CQJwinUMfXYl036kyC5x+tVT2lfPYs3sRTcQuy4DDO1a8mGSumneqiKPimLDEFY4HHkqsd2
qH6SqWMuBTEQ3VMUjzstPeqcik4d9eLCzcDmZ5uo8IJKyk7fZjvogKnSSxvK02MjrSCSRLgvzAGr
s7vdtboFCwcGZDPdZrnXhxvTi1zDDn8WiShxoewzbp+5v4Jn0Mv/T2wA1ePEylTnxxhWYwyz8c9/
fkbBIgHauGNVSFjBuVjSKjjDwTqveAAyDRqQByYgJbkSij9tIgfSaO/otNie7/HA5jLDgBLLWo5d
kQ69AfVXC5zKupaHWEW3hj1FeymlzralwgvKOyeY5n9O1ydiGK9Thz5jniKgQ1ts9pb27doOPwhX
IbbH7Xtm8DDCur4qpkHlWMYpxwtYfc2892lqtSOu8Y2xPIngrfsFtNCBI2iw0kCKaJq8+cuv1Myb
uK5HzcWLZVf1D4T5J37AcH9M6ughS4HCKG77PebAwvX9iYDHnJ0vMJwni0F5P4hjH3cTeFY/e+2r
rHhnD1qY4Ku8voP5t+VDlW7pLSlOMn4qabWSf6WO8OMFvYflp0CI3uVyzeLeepjhoN0FQ9Oq8XYW
bpgzblnvGCybaS7zCHCdp5TInat9BwlsBaUhubPPa1vH3ZZnvDMcG+dFVE808N/+RcQoNbfWbUZP
TYBb0DBYdOQUQbA3FzhX6AWKcs47e8UeneH1zSeej/IwmBexwDiWj6mxdVPntkbSA2iiZKQnXxe6
9xYdgqbUf2L4wPWWHJieg4tOAypVPrwwLbObPmVPQNRMuJl0fCInPZsdmCPucOn3VYrscXz88ppU
B4bIG5bD8KWTWSAVZx5aVbMPRxs6+ia38Vc2e5JSJevMMn+9rhTaMvnHtPlpMhuQZrNla4aBqcQt
5ZgG69dzUBy03ARoNWIN+RpqEawDdHyUIKZZ2TgqlmrDZqZXIiPtA5FCt+qOhHjdZ8JIVQngHt2+
CZXqzw5VwhMEDJvANFFz4gpQ6M2wDbcUHuzWu8/OreYd02tvw9cSYNFYSt37cQHvTgB/QIrfwzgZ
0jT3R+UA7omds3Pph/7fpOl8Fdmqs5VO7ZwoKwMeP0iQ08AVX3bp57Rc3rW8lEfzSONFXdambGPf
0Z1z1BHa2FtgMk++LNtx1wkx8WRUJCmpcCyLtTJbOSLMAj6d12v5TZvMbfEsXxO5nLIvleL471xk
KcBGrCdD8M8XENn67ZNR1IHqeTNjRAqYS/rh+z+lmtWeuOnP8qeE5HT8d5u80mqmYejIYRiVx07Z
Nsy/p5xqX3n1kv180/CYkP43uNCx39vUY5XZyqEtn4qpOVXYgkWEpLxwMKEV/P8CbzJ4PJn3g2/D
ShUWpnPZkVZbQfiR4Ku5WgpheOV8PxGJP9gxmejCqexjvQLs992Q74FK32IQej9gN67slursbuk2
gY9e2sF9Rkw4loGrl9fTFRSgDhIVj/Lx2YawXx+laKri8KiiQe22ENO2dChig1twUiJVKF7zGPxg
SChi8rdyZNUTI9A2crz13UVEI7lWB6v8QjmatdMkmfyEFOwFPuTpl1cNqnnZGLdTQpkXIDNyX63N
rHxa2OfE//tYh0kYmksk9mtV5i98hI+gvdB21PHIC935BrQo8ORTesP6TCUNJpKe8bj6aX5oGCIr
KOP6TJgyf2YcQBThEYa3ukG8pBrDC4BeY/ibixU4PgZNJ6x726LKodauIO1DGgXtcw00pVesYlmp
dtZXMmRAWTRBfNP6dGbi5C2ok0g21yrDGLOCaUTWQN4E8FayB9uLdJ0Syss98kKHP4bniTVPSLvs
GpxWPDExMjOK9QWbaU3349QqXazgAh95FSC3/LaLJMkWgNpO6Wj7Qi1uAjJ7QelnVUGEIayjxO1T
8vNROCr4Qg45k/SnE06iHDas4yPG4f6gFj2oTjaicFl1EUQvDD2VvqdQ10cjQZOoq4ZUcMFHi9sU
uukol+84tD1GvTqULEgdppDzB2JIL0Z9HU6JNl5OxQz633UmVaQ5bKqjDweeKs2r+y7YgIF+u6UZ
7ElAQe4sc5NRQhDWtTvY6L2wSgPfm5HLPT+vD/0mtdNYr73/YPJwEH0PlqU6ywloCV/G2I2uIMUL
CxH6h0hVH5/pxQ+WZQk7ExZhjkoOgUbUJ+Onf53kb0ePjSk+G3Q+tL/7qUdSyQk2iteCZL/EFH0U
fh5Z8H6AX+jAvFhp79GL1mWzQGwAQQS1JH4wbm8jC7MzcjB94uFtX3WAmLvXo4VAOidBX1cRNr/i
1w8Sp5jaIPT6adxxOIFI2t9PwCb+tjM+8zitiK+RUFuXHODN9CMmMO0XY4D6WddzrTCTlK76f2W7
geJHHY9FMwmtbyzwnvN9j7aNnBij/VwX84Km57CFqnRaFlQ+bZDmWPwwOxCSYvrbXewoefr/XbZG
CQpS7G2WQ0r7ozoIqMd1e9S7Ilc2PFGkdDxd9FeCdqFg8KKqFwTPTqxcGgrshk08E01UBod+FNgL
qcLg8zUY0Vidd4uLcb8ljnlYO5CYaUsItWzMyjR5ZyzalV4YsGQJ00yRPP/6XN+RQWLZeP99ooLp
dxr5Gf4FR4jM+MSr4IqUUWKhgU20kaCq4EjYnwavceoPzW+R2PdbRH8h3lPDrz6HTWuLYkz7E9My
6RBckEIl+j9V3rU1x0seeZA864dqhI1YJMSEtqV+Hc+Z/JuEupeu/gP/l+X+5e485OmhYlmInw2f
VBNYEw3PA9mNfiE5cxCxIwy+zByzt8EMwJiwVWT/Vxzz4FossmOyKMY0jXfD5F+zhfjKj2CHc5QC
L/KOJZqJxu/orv2Kat4sCQeQa76+LpCt60ocGa4ZMr4IVwRxrsd0o7pJN73tQNhQoU0WJYqoRkFE
dSyXWB/6Dl4ma4fiykPimJ/FZhAZDbK81C1+wHuzvt8Ddu7Ja545yWScrO2mm5jGfvngjcAl0A6Z
EqvBBcgSU6MsQIQgkmpudOVa3LqPrq8OACOjx44jF72Ag5Hw9rNNiVqhvlWTULpgq0lqaf/ruqYd
2uohG7cWi42LXDVYG8v8anwxB4gT/NN7b/CSSssul7ta2KKvMFst+YGbtaCVXDledjofJBuQbE+j
8VCUiDndr7UzHBzbdt94z8qWP3j8D5tJdiZb5pP9yE2TX1htj4H8ndXI5bsw8kN06cN/ZcY5kZrr
1ryZZLppto1Z8z9ELE/fN35pLD8SyiOtXEwM+UK4qrJf1dcWHp29xBUMK4EBffQQ+E6o90FiSe/a
7vpgT0aSxFBJBg7Jki1dInBq7JBS+yKzwcsRMZ0zS22dgtpZDFvKDOxqH1pqfuhlA6Lv56Jj3bXu
qkrtvwFlGiRSv8zWPWd+Ovxe0Sl65p4o15yV5QQnGMCZ+OxMrEXuCJlwW6A3ah5ouBd/LoS4Gv3d
typhEUYwsOhJynZnbUaf13z0orGuc+oU2fKg2ZkdnCoViTwU6AdNUhD7YZ6rgnAjtTmsik7mTqTp
aMsxxsm20HeubcXI+ygGphxcIgKChJPqDnCuGb6/0Ahpqqt6qjglO0ff2ovV6hM1/dt7OIMhAKsU
1Gzdu+tS1tS7zcZLsvE7qMKJyLScFnbg9+2pg6ZkWPE7MXj+fIsLnV/gOYcXLKg8+XeDKTCyqjOh
RNFwmghI6SQuibRYNIzuW4nL+yf1q9Cjd3Jdj4giFwrCvV87N/un2K5yTQdbNJdYxxcvjLMO+NqK
WPPWOFsoN+ZhXpmu5LUCodnOf8N0S9hnAHI7LlwVW8G+nvyeBq7bwON+fL5jOIjgLm6pmYaFDwxA
AeuQETePBIuTapUkjjNBXd2jSNRfsv0E9pSGJLt5yO9i02BO/ydja0+0uIyaUcpDZAwefJBOkmxX
r4VgfPxi2NNyC6PwePmz2q2b2REDp2Q3Tk8kQLg429sCjM64t45O4l+yJOgv+mzhHIXVBNkjwF9t
wOW54eySEs8kG8ABZB/gsTitRwk6wTGctQ97ysa0TTCaZgxzJnRaW8R9vxgf3986QIh6rrnVjK/l
U0jB8N/BwOgdKlTKeG4gg2qdXnLXUdl8umpqo5OGiVp4QEIYOnL7m4cFTQ8nCnQGL4PGfYTI3c8r
GsZRR2j3uRLw22ij01N/lgPzC7kX+jSfxmp3ynkbnPi8CV3K+TkDQVZ5VcCN4HDkveentCbSWBrd
fUbxQOur4qLXlU7bpAAewKBfYOyfbN+ikgvfoIayLokG2Af8XyBlaWnfNx+8p8cqsXZByJNecqDB
ofv00KJ+MrIbFqgbLFfgQ55w4El5pwkBkV6DetRF79fl5iKHKqBS1OQlUt4lqqY9skQly6XBWYiH
JAmFUUIRlVPXl7hmvAr+v+y9XK3UUaUeQ+uzks8TtOIpGKEuZFcn/dNUw0M5aFZeyYRX2qIcSesQ
eB0dtOnF3euEDtXhSWGDqaho/9U6NunkvGE2yw0NtBp/UsdYgEF+oQj2ParEAxAhjigNH6rc4w8J
0CYzk8jQeOogHZSspf5eXQjfoCQwEosfr7ZzOnKQMMLnX/LnACHvh66KiuZeLK+rGYlUmzfgkrxa
7vUpULosXQrG1r2/NEU1AMT8XrpEz7GFXQBDEZWicSYYZhMM09sP/+rmMvZ4SVrhdce6lUShsC7t
hgDeLdwCjhrlgcQbF3D+I1SWv6DgB01Wt5V+47WdLMmetIuFTdyEhoR/YMC4TMVeXGKKsx8lQsdM
4CBmRlWXj+PbhWqV2HPJOYZTj60imobkTa+4+sa7UkiqAquStgyHi2FUR49mNj5YlsoKtgDBjyoW
qvunBuJqNGttKCCMC6BqNpE+AMCzo2GQ6Nw8WsQlN0/GNLuiCSDnaycTQEkTmDfxDaCJY3hrqOl8
Tm7vmUkfxegROYJAbiU08obKjygYJQCSEIBw1Dpb4TIsCN31Ci2Jq8D7eT5RvF47EbyT7JFsqylv
KQyCnudR1L5P3rqz0AaLCjUSNK4spEUpel31St3NDqWyhaialOzxmwyE6sgdvhhxhnVQ5K23xJMu
/aT821RTH9RYqbE1CJlLXI6YvQzI4BqBh1D2ttN7/5QMrEetncK0Z+JCgMA5INr7MJ8TeWAfCZx4
jEqp6uja5DaUykB9tXhFLq68GNGJoWgHjKYWIv6eBhTkabGceVau3BWpFT8FYPJyCQ8L1KbUrV3m
qHIynjUZU5WgRVlPwC9o24TvDPYz53wY2Ukxc9RXZB7LVYI1oBo+MPfISejbboqLTSB/vIWrbfN4
4i4Z4OM5EMvBMtRwL9rwJOpq8xhzg2ojNGzojjFLhmk6fnjjtGT7wjO8No/BXfbm24rVAvtlgsDu
Z7+ilz4TCBIiQ4vgpWqHjjrLm7nsCAL3buy9GcoPyWSP7SXxKHj6gBAItemMYhG4noIYW8mgcNoD
8JPzL3KHDDXntXtRD+9DBnmULuDeBmiqFa/uPw0lKUTdzmRN4EfQd5X+4sn3ba2AjeCkNOk2kqpb
cehSVB71htj8sKFSROLlsziqo0FbEXm5awjVs7kn1dH61DhvyBkRN4rRFuuLRTyIAfMaTYDXRfDd
XWgussXgCLs74RlTneeW3p16BfNYJHemEcBIYcEu1gysXNNmPhAR8doXMhmuzxh1hGaydFgOocXF
s9OmaWlS3BkaYNYs4NrUUhVQQBB8YEM/dJHSMif5spBYpYmyK2HG1p03WE5g+V2pXhWHApFaFxZT
GFd9IJ4aHzaJQfb6yegpJsq7qDSNOV+MVukoZSKsVhpzmjrsihF6QeRVLlzsBcAPT5xBp+hb8pH0
clxlJvHaXjA/yxR+kFLkijg32If2GirG3ldDU0LHRjwMQ/WwaHBX+BmlfsTEDC4jJEGgbnrFEqFw
rO701iu/UyOwbmlqkk0Lv/37ZVUOnsDFYNI2g3K+z+gAYqJ0fQrndTjXSQRe1PWuaNweWg7DomyP
jGkURD8POrmhV8QoNVC7gGBCKlbEQ8X/5xsg3gQwE1gKxAdXRsm+3QXPiVZ6UkRp8nCmqJGCUE7Q
MavoSCAy8I3zSgUmyGHMMEydjD8MKzwILQvsg5LKGPl3wPU0mHPsJpH6YVxL7IGQT06KeMUHni/x
AXOEh7ma01u4L7Cn+ekBFy9x/LA15y6H3RC51qPtdlS0CCclWtVjt1TiIj9j+SseYPvzuVksQ4z5
3neiElA13wlY1tMP/om2J8/jLOHu1gjRqdQgtgmXu/3xAN2oglyjQ1b3yz1kCZ5QsU0/EPz0K+XB
sc1ixZNOfZ2z9XRzkog4x7Hxku6G23H3+mQGH+8sTaRf+Na8f/NQVNqGM5ZqORjv0cEgPtXB0QhV
GI44XCkFUdBSH9AKtb+zoeWrwt2yOCk99RxFrjC/dtoaqxnP5lDXw+Ma9UsBcEGD05xS3abSdBFJ
4d3zf/1LXLhh0qYKAkyvafqWl/pMIcF/nSs3vPehcgmVl7Qj7yGJeahA4ruoDPI3pmiTdmrKZcBf
Y15Gsye0b3CRtvg1lVG4weBV0gUGItx3D/DyCny63GfVXsia9po4eR0w8vT3o3Da0+oMrvSuPG5F
ASjGUOxgjwSu/K2Nz9Ls15JDmtepg7L6231NbVSIhU6qH5STos9HHz6Yox1JwLMXEUX6YVxoOYf9
TX/sJgNXQNwjODBc6ao36XfpvHrjfUuy4f8Otqx1FXHa/xn9Dl0wexSFkWBdCcRmkgs3R6BYh/ec
GeLte4hk4U+PiiEFHePfYrRRJBWEuotsjAuHBPVMWsrsqTiMhxdIbB8pu0ww0LjsrHY+COG/BbE2
RHYW6uVonWRJPCEF6P3vdHrNVzB5z0tC7Wo1iZ9O32uwDVkc7fwPUu8NpBD90c0ugw3lxHzq0KAS
+6LXhYkqYlEkyehgs6zUM2ySuaFUhFkmNHJWMTmB72d4wLwYKwUMdJbU2hJk18164W075fqdCr65
Hy80SYbYAa0fysf1ea00sP72cXXYlUfoJGqYzcupvhNv41lcD+3kJ6DPUO56xlluqwvr9OQlh3dU
UJPA+dz8NBFe6jaf/s1GXdyuB7a9wtTacmVBDbXvjaLPRyv6lF/7REL10VnABZqysPDKnsuW69+D
l342r1gm1pLJOHP71tKD6t7XeAsHf5yslQN+6CZ4fw0KCnuT1bPLpsZBUkuUirCCjY+jKdA8GaPt
G288URLt1IYksp6eFTWeS3ScT5X7AcMNqNnw+gfisUzvAVT/6gC7Ol+MhWmATg9P7gdovFuVMHHr
A3yHBlG5n+9Bh7H9WOiZBZiG1DP+gv54gr9y69T0zuNkOcUeSHMKE/ejS/mOZLKrRuuoi18uMtG6
b0/Z/y5yFRQSOanZ7xHQm0tkIhKaTFNUUjdX6iN3QEGrTqtaZfZIBJgP9VfMBndHZlekN+bjdjam
TIDqMfJHg7F6i9RLBmNrG9TajwUd2RtDT1r4SDVJs+gc8jlZMnom0qsH6TCA7vGI+YXutBFHr/qT
cgUwL4D7Dmf3eY1QBF9hS1O5QBAw+KkDOsl1GwlWFRZgmCN6A/SGdA/AUzAi6B4Zcb2MObY3qE1G
kd1MOe2xW7fnp9I/j1QIvvDtGxHBCQ2FglN8hP13wrLUCldlrORdrKx8BP4W73zIe3p30918ZzM3
oAL9SwxAbFsaN8yKQrUYcWZeSjB3GoYXh3yqDaYGxhTrvrnnAjVH1bgbJwqsvB6PK6kTArUxh773
Vu279pP6nnH/sv9b0V8kmqcpoeq/hpYYBIg4Mce8TwXmzpBXe9Ewi6978fJ0rLkS/T2BwiqXb9K5
rlAQDyXlb0SP8QZvSsVvj6JutZc7AkMmszWn7QF3hvATQNN7PfimBbNJZyqvgLSoI7y8yZXfbunU
d8dymK3/mldPfj+htoMMUorfdx9kUrKP2Dcin06NUX+YyiYWjpaIz1GiMEAhTe3EGKy9ojzN3DmU
VQn2DYqeSGg5EEKfqiMa1fzcktblEgWOraqY55iaLFct9Nnq1ENnFfGlZU5MmH0nQ5v/CQoOAXPK
7yzkDC1BjQR+3d6829dscJ9Ac4wxJ8jvi4b3eGbWcGH8QN/pGLAMzoLbjx4n4emaaC5LKWMl4VCb
4ehM0HNKomN9CtIodpIxu9ruWvoDuSQpBjdTIZWkes3CN+jObwKKe6KBTe+wv93VfRaDn8g7zIde
vHLo8UgXBSIlidpLjig7cql83tg8M6Xnh6sXL56T1k2CmfRBTK27xvOlVqUvdaLxY2kUrguq4amg
CFn4PuPyOaLQR+Fk17IG0AuVo86LD6mBkjc3PUDfSgK56OecSlo+H+xxuLmeUuQ7o+AHjBgW/FqT
ZLCLaLilqDMrRDRJJQm0uodSwXdupO6UciSOXQxIQ1ruYPfcz1bM7ve/03UhJGWvc6zuUYYcLoqX
UT2D+HFGTNCmiBDijq3L91T19VwUESWCaJSdEc2y/SCHvbDTfUx7AsD6ecAcxNEcCqAUBYHIzTRQ
/2SWoGiOo5xI6SQkZ/pQMDW6xjAGsgGG329pwYkw2cnPFOE/J6J83fhZH9RKoBp5yWvupXBGxaCf
LsoacqSjwE6rKuq9lVtik1O2+BoJ5vJFYTgnwlrSWVKxnaT8Bzh7GwZL02+zShFJ+XWCgAT8Jlqv
W7f2+FybnbSFANVKQaTbCKm2Zd/Vg9XDZIbPLKzFEYKwHbMStUIrvjlJwWJRpvl3rGrrcNzEovQm
rMZygXhdEzRIyEppO/h+kcwk0XvlKZQJzyoTBQz8q6GNAz4D6U2z9SXWSuMLA55xen8LozONTTEf
mMD/VihJBuiZ9KlSG1qd/J8sFdm60Is64fb6lWiF15Ojs0UrBjc1JeW+/gmZDua6gQPeLuFUDNAF
nV7O0iGIul+5C4D2DET+fG/BUP8RkzKaZvrvKIsxblUb6w72EuXKQSPGHXyWd+NaCB/hjSNE2pS8
CG09FG4//26LTxJ6/SwxGRMFzQpeviITgRXwb8h5CKerNDDMUZ80Jv3JKHcXepuwR0xo+ji3uNjr
+hX86chUphDtVWadro9S7vxxri705cSAUboIhK9P7Y2ZnLsQeH1JeSW5qXyK8NcLDtA+f8soL2fT
tJt2ufpO4IPfsKnWCIGCthVmhwIWwJo26Xr/8lSpYhtaLpwvKtmPi8adOPGWp0zV942YT0v8FQVO
0lviITW0oinks2mby7ESPYqgWPZ6cyds1lhA+aQGM7c87ZEthmWe7Ekwqc2lRLlFnF/4fZJjkOTD
BXgKjL2pNt6DArTCR4ZyhVuuaoM54pvEBVe+e9Q9hGS0XQdLOQq0ozgC9//xhz29ll2nPtuJ72Ys
N224mj5vFhfYZkXpujvYN64yzhnwE4Lv3cKAFtloozlIda6jvWvQhQN1Wz1hNsg3Hey+9i5jUyYj
mQNu3t7Iqf8iUMrjU+TVH9CNA1UiP9Us80XTfezR7BEou9eot+AB3bpTroC/fkfWgaklLNR5l6wT
u2/leteXAjwiQbHKHzktch8+e2M2r+TbLTeO+PE8yv1vXTx6Cz27FAM9tjV+/It0nIuHSglSoqSB
88+PHpFnICcP99WTFrP4zHaQYjGMfeM9VzmAi4rIknrN28N4ms3AZqlRQtYBrOWer4qzgP9xF5KP
4ptAvTFLFuhl1CjKrmVsgDIwAZh0rVtF+gsH3NKbv+nWZaw4q9Ruz+C6q4b3cKco/TDcFBT2biTf
+W5aR1L+Exo/o9HROa4d2IB8lUVLPsgXQP+KlAufmQY8y5s/WWeAERrSy7vKuA6KZBY/sMJQTx6w
2guWdmdU8UKt3BBpGPDsvkzX6AbseTPSLMzjvY+RwiDqYDGw7qGFpnTixZ+cGi3Lllnt+8jMnfeQ
b7kx4cU5ADmOQAnNOKXfgjr+jKvIR/tLy5MJzKMSaJGrBX4G4+4ewBfnw2E0TgYCNBxaZPpXCd9W
Ggej1lD7zQsIG0C/TtLFhaFRmsle2mKcgnKDjNB2khMrGVw/PNE1Ey0lREHZGuvp3sISOd86MxBd
tPBAxyLp/UKk/lEczQN9G5EJ6vvl6VNCA8UG88dybI2EjqdH+c+RqWVp0Rq/oaVEJ/KQNbcTOfRu
ynJVj5ZgLXFvOIGd6B6qkhu412OVNycItedk8bXeLKeo9KgbHQNRHK+JBpISyxAowJER+loiw0tD
elzc2K6gk+ur6NFAp72VqhoUceebl3v5BM6iQ1nY/Fnlx0q4BOtFrgeM3KV9RhTUnB8aDJ1Avqpx
A5gVSam4Dmqbs8M3xH7nNKv87dUZYUsWd55UeMOoIfl6kllnmCGwy1+AmAJv4SWBfUtpmpSyyO8f
e/Q4biYA2WYNxvsARu047NPhJoJgMbGbIuYUBT5H5kvRLei8mvjunwXWxkh5+gcV5WMzm2cndMVT
vuMj6Cnc7A4r5A21N9pN6KxQ9F0sBf15YxVnjUO5KmIcXhLOzZuMH2ulpIZZF/47KHpyppKnJkZ2
rhVAdEhCHPflxU6I0g8pfxPj4OTDjy+V3TpEDNk2knEdWzKuyKydlooademVQ5+1XhTyOWF7Udf4
rA2cS1NDJyJJPQ8WY4lYUU2CZpcSDmbwrgBiAEdZrQklwgLTHbTrcdfy+XdHk+ZbRxZQXo78DN1z
lXBvGXZ5abyMZo/Pd13XDSZlusCJyViC9a5M/G1qz0AgSiigpVSPt9l6FSRiDI1U8JJRBwRnSIdH
9x7bHKnXPIcQA2I0vKXajWUKyyVO8EIlEO+U9o+taDKi+n+A8kYsR2lUiqQePbfeHbCbuAX8j+WD
/kElOBpY+rzYYYkttrASRClQ0ITMhbo6DubxP1fGOAzPWGEYGvFeZzXF/prcmCe0wjwXWr1HaRgk
OVWSPlov+w5wAkwH6uLgPKfHL0/sZ/9FB89kgl2ZBDDZhwqi5k+ZDrgfTYh9wLUQCGF+dY46UVjk
nGyDQw08Ol8cT7deZOfxMlRHzTHuxsRa95MxYEocBw+A1gcE/DxSZkL0gj/9fDJ+r682uMO1T6cT
NpLuDsZmoDRp+nLXiDnXWaKKv8rHmwHJ12wZvHWaBSRXtMO/GHvFekbXx1aKr7dn3+WAXNCUSkK7
zq1vmD6yOy+JOqlbY0W16ji8DiBdTTQnWcBnkm8iPkkLu7ax2wfsATOJOoTfyg84CmagYgGUNS4N
M7qN/VRcBe1Sg+ZCvBwJ+cBFHfM6ZT1wky+QD9xKv49uJdjoJ1ymlbvRURl67jbm0Av+nqcJkQ5c
+qt/4jk7szArp/x6hQOv+7Vxk/5+k/8BYNi9hbCQ0viBprWcWq7E1wqFeGJJVFh664oU6ASr+fcK
q+NZxw0b6ehAhas1yAR2awmjrz8oAgmXgKeEMQfl3EM0fWSaVSwoATR2O3QgjvZcC5mRsXuUF6Fd
c+cE4hiX3SBtWazRgk2AIaRG1GyeMmXsFJEFIkDtt5vvdAZROEYicnbgh3Z/x4IVBrJ54LGUrhTu
piXSnEyolN/l5+d2IjrFnjm4gQeWWgKlTl4gPlvziXWoP+ty1Uk2RAMYjsfb8H0+f2xWKqm+hmhj
+RePIE9HZRPRGJTlV1lvd1YQz0PtJ4iTlurQtWQF9zNIUmfjhDTCJj9kTJOXajmzZOcsSh204/OZ
THJFrF4mZK+akjrqMavMAQPMgnA2SjK92Mmy/UbyojDYIQRPgnhA78rY8NtNnB6My31xrLO8lc7N
OioCJw+WdJAqopScRCJN1q0d2SLxEghD6KD0STpFVjBykZrNZ8wguPWYOVejtKX0T4vluj1PC4Fs
nouPHjtQb/S4XSdZ8h0aYylrQuKf3TOdyq9pV1jqNrPX1tZX35SIy6WRsA6D/vZEiNdMWUxMt/is
tn/NqcQ2OtzCtA6CwrGetQpYYx4rBwu8TCdtHAyyPu9Pie0VQDhslW3fn2mOyCqr3+c7OAbNtvxr
TRU183VqoWH8JJBSwI59o/8kSYjjJi0bBygn3jTnvwHdkkUKc6Kavfh0JXAY5MhAgCyGs5e0F2mh
AsrfUzOcCLfj/hjl/1k58BOKEVsqOWDe+SNxjik3SEJaDFlTxJlvCJEeUsTbJQFUK+CYMQn+65Zw
ulknri/ekE6+ZqZXqTbwPekMJteK3IZBQAd47UJx+zybH1p62OrLuG/Kl0NdVZNi+GxBQI68JK9D
b++XmG2OpeJmC06KULFREqlTmB2ThIVaZKhiJoDyqrPM7sihwvHr0lT7DAhGTg7xfxpgQoP4eqe1
jY+fzmeuQr1lKKWEMZHOL3h0MW6swrgFQp+BkRMh6y2UDzDLJ2aI6bcwF86UTsEvJxkh8i+ksp9M
9+AqcUWv+bjjo9XtIAq5jQtSkSgIoz6TAElkSxvO4GlrOHwhZyQ+o69jqwFAYpW5qpVox961t7oE
gbq1tGOp//grbZzGoX7VZna6g9q0mrwgq0B/XrBG34UfGAbZpNfnnPWTkO1covFbsNnyY4tn7Yd7
irmf+V1lJmRytyP8J+auylWRTHMRrYRD3Ca92ZQUAHztHfQYhrYLvAoKw6j1K/HndLobpmRXFUhy
QqmkIl9GF/jndIS6ZXnAR26mgH0esS6dly8r9A1qklRG11oUoDTwFA33XFiQHB54F/kjpYBDWFLr
VtMcIxvV7kuSAbd9w/huVyra71kr0AjwZsMtJN9RJ8s3deyQTs70rHMMVNjFjfPrFy/s/0stAjsf
3OUMyo1jh+Xh6imkD8hXY0vZmBWcFLm8OXmFxtCiMPv7ghpoPA9g4UcR4dlIT9CjaD1r8otdmwwa
/4akn0xiHydR/XinxyEA2WO9yT6m0PkQCdWLjSYsvuR6XauwyCtYFAZKCbkj+DzJQqCHz6NEaqnd
9SsfHREMFEB0nUD2zBH7hG+RDmksRWJ787v/N2kALhjFGL6gU3BRy7EezuU2NtnloP6c31HNuW5d
Z7aHjhG1NZp1/+p3/WX81h3l078lOEUSnKZeoZWFklLu5Z1HI7j4zmFnLTdJIp4ayRLz9FiyiF6E
tainXIy7t0Jw2W4bMf+tqXwRo6fMD9mjyVyQjVt2/PFfTyzvJYkV9SjaW6tyZbPVirfVQwmPJq2z
ShXCX3z5VE3wlYK84VEjCrSk5q9FRYzeMrNu+JmwA1Jn4AVjXWEurWXE0gknU98mlzSpY/XAkdlz
pFp4IDvaGbRArYtjka8LAGHjs1XlmZoO90/UAKlKSU48WtkAyqbpnwDT4BrmWb2yAtx6fYQ6QVJ7
dxTIobsaODA8VRmA9We2dfRiEo2ckCh+U2iY3eXixluNUDAR8xJ6uuFwu3Rh+bE1lhBNyoqy97NK
P5OItyl+UNEWGCVRgpbyladVl8YTwHvhJZXxoz8sfu5EI+7W714Emx5Il51EMgwyrRpg4HTHochx
UOJun3eHpAfyE+Dh7kMfTgsvN8MdOAwAkruqlzzg/jqVrDp0DAe2azUBgCaMzKvVE/8EVBG6EOpV
RcaaV9faE+s/CBiHExwpyI49QHCLKrNPW8trP3H+BHYqsnGCnxWp5qIoXURhnl1iykjLxZcVkzqx
3Wm5IyJRcWYXTXTxFIFmna+K7oSqLkhydND88a1LD6i/PXPw74mZE4BCMIAYuslB8Rm827pKa0ZV
eG4qLfjpmQefGjpN1/Cgd9GMaAa8wVu31crL4grG6kgblqf+BZS95ZSepcjGm8hz+5rTHMc4R+3C
lHlo35TmPg5CDgbEjEFehQ4SPM5GJmlddhiEu+7Yzv/fRd0OslzilsMbPxVdWhAB1j658sdsnMVA
cGQQQZo2r+pVAu4zbro+GSPSoBXN7vON23b2bw9BAW14hIxroK84qhJUv68VMsqVVWZwsgFu79Fv
fvOzuDUTA1/iwNjTAQ7c5exeoiSMMo4zRck6Xc3z5cxGOs31gwnZqV2Qs8RE0DyJanNkanWNbrPz
m+UJAJRUOZeoIDzcIk/ghx6peQYT/yqZ1C+0Z+RFF2HDNfsywnnUMjndnYihTjs3vJVz1oOnlFdB
bsm+68iMEqME2re3unPUDlKlQJjZTMxzlJbS43w6bBj4Zydph8vPF1yGrenSWhfpADbuuksBXfIY
97MopoqdjGzumocm+2yHMIFum+IMIyNwUlv8uCJyrfKr7b/XGB20r1bT9F79AajiqKLSCHs0ThYU
hWk3Rh+Da14/iI729WjA3juyuNKKC/ySThyZtOtj78KQBq7jlMUuuMggg/o2c4ZuQJvDahWsOtiw
B7SSAUpvLCwLV3GzuLeOGQyE/sHmeRQTVD4ANd7dnUgFvei+hAkMN9v8HCd0W/SA4cDogoK2yaR+
u6A2zXbmHYW8TaeigZ1Bc1OIjBEsI5CSypMpo4j6ZpH91hAvjp4E5AJUVUT1CnLKl4Cyln24FM3p
VbfONVuSVSjMw9BMwL0lrrFJhld75qlctQK8gZT9QD8G+4hdY7m3ymaR3P+4VwRjqeDwwfBpj+em
CGexMYKIFIBW+WyMas1cLpXo3x9mQogz0JjcKU14j3Ka+ONasvnhldSIrZWf11s2coFNQpaJQYDW
tHjsnDzjpS6bjl7z7TsOx1BHyzW+xR8TLZciw4NzdaX2/a4WO4OMnVYdB01W8NVigZg8ITSnOKB1
di0NJ9jNIYBFVFIADO5M3EyiC5sJ2bVEEqLcIQ52o+8xpX8F+sp8jkp32RQvRw9NR+8hWQE1qx8P
T93tQRvOow1tpN8FpnIhIlmtk4PK8i1A6F8OvexVdz7cl6RxCmdmtvOIGIZRKNhiWDuvgjEzEO5I
6CgPTdtfSdtLx0UXPGFMoBPZEwLR1Op1dQa8GHCzsK1DmY8pVvu4tN5xlgbBZJnbFNIoNemKTw2J
emG9seUGLxsnlbII6oVURo0X+lExv33TxwZhYFs/2L/M/dy6Va/lQpBd2VoTJ5LN1wkzcs11wD6G
Cg6t96dZt4zC+0bwOxpZftdFgDW+6E5X4xtDGWifUxJ6dmfY8xvFa9IWMPDZLP0xOB+i4e0jkzQW
jAUZDiHJA0MTKZuAVq6VoS/0HpXw2UGiUbw417RpY2Z+fnrhYHE4FrMIf/YH3j/RjFpIxSuUsvWE
YE361CXeS6LqaBqXPjp5SItwuvjdaYZC+CFuMHoAyUJxF7qYW3Mt9Wxe33Tun+pICgSIhUrAu6Gc
XmfoOQ5B3XIeKCUm7sMUo8yqXFKffftjdJTOgblicq8yrBjCiJ67N/Q1+HF3/Vw2qJ9Xv8YrJigM
Vzr9xgbMcK6yajYtCAURxsCF5oRFf0k8DqhWvjvgvFw7gc0W3t/+CQadC4G6zvxUasgU+6t6PXi2
IZNJiWKPjkLmyGb38FAjFOeGm/nD8ByYfC0IFQCS/91/3zyrNQ3998ANQ+IqmJpFqZDrkQFjKpdr
nx2nZV9RBCMKi5MP5zQr9kvFSSqxhcDpm4k7vgtNXL/un274RgvKU8o8AW2PnubXLeX54Q9RC1OS
iaI0tsnEj9XaCiKk44xTMFXNCS0hx8VExobMypaZoDI3HhKDhOBUFdB/p/yfqeiMoxGmreYkb8aq
KQXl35ZuQxcfPx5ocNBCes56LHY/Erb6p/JB4vQ+S7kowzY8yQIQxl1Rpz9ySoUPgVuFtJQkkRSA
aBmkbApjLJRmKPHEQXG1JBSL3FhljYIAXJQJBvfm1oGomuQ8mJ/iwAjHURBCAnDYOFQ/Ea9RaA0j
sLGASg01VYo3cbHr7/XnatRnNBPHjJAoBruEXM9H6U2F/mjKT6L4DJ9Kf8J+Ik9L8n2I6aEovH8K
RbS9ht9VgMATOz+kC3R5gJxiTzWmuP+sJqQnsAP7ZPS1UoC5wDHRWAQUfmmhKLKC2aYT0IwMX+Ah
93QGetNVEzQZhwaVRK/+nf2obPe+2s2+hYJREliS2b7ArVUpz2YTBiYySqt6i3yk2oQK6BCuFfpX
L9ex+DcKFtLbAvQl3F0EEHn3zcpjlkYSKmINqqwews5SIclTJpqwBzYYWf3iINupl/z2eHhpgDaz
Gz+NUA45HS5HsP8HEVVk6c8pYS6kNSB9peHbFvBqnuik6yJAH22nEX0brgL6xighlnMOK2aZBza4
aGiya29P7CqX0+NaRcTxo1Yn7Y6ETiR0z/f+TVSqO0lB7AhUsCfmPXt+Z3Md038GhJ8fp65BZwMz
v9mfZa5qHACQln+foWFltFvkk4iQerj2lEYVnHLEL5WegvskUJas2mhWmuGCp0ns6j3hOMTzx4C4
85ONnr5Fs4WP2xkuHcC7sW4CsICXpg+Nj8TiOY+At12DjWoOh2banFRD8GNvCYIDWd9/SSDrXnyM
DwsrdjCB5kPjSPbmSFiQAgXs4FJsARGulvb4BQypWCPhsNWfSVYsC471MAJnbfV50K1M0W+ftvhu
7ZZelnIYlU5lQYEHabGz6/H6dq4a0h+KRefkycX+VGplMvhd7/opH0F+60SOCR6YKWZIi5caTEqH
0dkVuOyCL/zXPUThnsSacV3zWS0EFpETVGTvmlXpTA1hnDyA4Cwj7WAqR1QWsAyOaU87sXqDJC3r
mFzWvVkbEruE+eZgnRbHqNNyaoTe536qJa0KlwIpjpdqqrnsMJsla+FuK6RLN2p7jqpvrw9tUwwG
ygGfB1xVtxOxuwxPpSThA6N8Mf5DWbjEVRsaG/5z0EvjLFAIj7G6byc2ACJISfusEyW5rRsxR6Ap
SvzAdrM+M/5n8oyt/dbH8+G7IcurGUZV6Pf9dHcr4cJm6etP2YpLv1CO2w+gLeMAZz2IiLDl/Zmu
LN+kNBZlQOfUWEQ+Mpjzxh5ZHuxtbM7WKrTgbaDHqugX5UsXS9gWheVEoSWPW7KbPuYDfWzx5mLX
mGIuOri4sUqlQ0YrqeVpZaS6xrAplIr/D3JqvDevfnUbCIwBU4g25lsVTTNQrFt73f+jCQAMY3PF
e4hmOAz64jcS2af8+3SslPjBaJ7UHqkisaZvkQg0LLggCBV3iQat20DYY+uI6hTxybCTuWa5stF5
trVApajD+bhFH2YBk5NJxiR89+qB+t342z85HQZq9qF76UrQW7IP11rIgUedscS8N5kDCCdo2PGD
S3Y7l7pXhXc0mPPpXVfW/t5nWF/Ww3aZc7q7VJ9BYGFxe1BpubTz0OvX+u1IZqKL53r6183fG33r
FBVV8gzlRpgDmqLU33VjmtmB/Uh1Dh5lqEf4ycD+7LdddcnD3TBZvfApbI//9UDqar/006tClXpv
bRaty6sJY3trhR+gFGjrdvCPi+pkaNMOY4602ApmkFkju58AVUeRRXFB6lmqcwR5eMBiIDP1FbVL
pgrfHGSoZRoRQATH0k2USysfNXzNrjcDGzO3uz3U2+/MRAQrXFEa51aMW41huQSbur0w0wKKLMKr
dna1KZD2dDQZpk3CRDc4GvpCMrU5aaXcvH2nUwCch0nH2zsdXOoC8RvbvYkq0G0MJ+AZnK9pRPUF
l+2eXAqevmRZd5j7srGDPdVw5rr8R/vn48ZG6b5EPDVshWiMuYdqezUTtgiSUD/FlmLYwqVoz138
L/DV1ZkJrejEIrP+ofJ1I8bkXP4QZm3RWd0+m+aDKo37Tq+FPSaFAAN3zUW6mBee26juFwCrM0OQ
UrpqjfdWNqzEAI4ySZd+85ziHuHJnnXIQ3GqTxBgg5k4Z5W1NMFllPc5UNYuS+AgC2peO1X53bFL
qZrmM+XIHmt5PBwOo+U+HYS0uwVJaM2+fTwgJeiolQ6PE+t3GxgXKdVgqFs3/E3cM4ztgPq2Puqd
JOOn+/4+XL4BbXsjVHX2fuxMAExZqdY2hLIfcbiNAavwysxWWxHUOfzNji85HV8HRq1KSEDfAKiF
kzfJSKfyFRSWRKC/yOmbqcEqSiL1OOaufba6CsUWGZkqUz+t171/p0lTQjrIh6nwXbHFaO8VPpFZ
p6gzco9xhA03hVx4AfrFHwT+ZIqKSFOiVUNHD1VegM9dx45SJNZ3lj6GocZkQoJVX+26HGYgL28B
F3vovEZrm4Pohd07TNaQ+jS+jOWxwDGWu6lUDp3oOQrY90VaxyB3cz4vxsL13wsa5XNi2M8sY6kt
6JUrFlcYWn29Kqf8OwOWn4VRAFEkpE3LciekE/hSTAgcZVSLECMyIsXZ++q+hR9EsqGMK1fh1mbg
QKqezcjqq+AMRSG96ugDWffYlBhPb6HxYxVojaWRgkSYLv9g/+a0aLjbsf4+zv3hpwKOYDAtr5YJ
9waB0HJ0eZXDCn0eu1U/4zUM90cYP/peybx6xFsJB+NdVADZNf7oxdFXusi03qA+YE17hLhl38g8
Sq8xEhNSSDtZ9sIJkgx/iqZfRFCtzo7Jxc/JI425EY9ij2SdDdchSQnq2XpwH+qwUnZ9fLoDbeRE
0RoDOJC3kASBpjMhQMT9LzgOwVuWIiba85bZfrZqKqQ9Cs8bjPclPjZ00tWSWLmO3aj4EuMdN4yM
cNgg3VQrBPfW09kZxpO9VbWqWo/LHq2fWT5YX1yzMqCgMfe3ezzUNj5LY6il5TSulLdcEasJXvG9
oMWeMfotVM21+Lm7jO9Y8OWFzgxTjh64DuC/H0cpbyHKCZhrGkHYIrRwy0BldCcyLn7B2yQNhLxS
lwUzmqMKBreZSslcvjR2kIy11r8FqL1LIfHFPgm3yPdIO5Vp5lCVo6PlZWCewqnbmUN/Vyzilm0e
nLqNQQwLz7o/Wgbv1wgiLU55SaM3f2H0m+FOMc4MUdcANhMpsdf1THygAhwfWJYNijl092uJ0hbC
x5SkIYN8OJBRu/CDui9ftM9MjrvNCDzURIPHrSzSmcT7/Cl4LAE256KHrWOjz8I6pwnIvaIrJmw/
HOhK6L85vdivOG4ubPiutR+hId9o7pol8KIk4+y9xwbmG+IkBo9RCp5TZtE05B1sLZ4OmIVUJSRH
NSTvJvsIirBo3nD2borMyR5tjIIkW9R4tPLG9CjqFQNagG3f1WIjf6AAXWIv11VZF+qxGkRlCg1N
5PjHoOixXztLpMZwzDPiANN2l2ka671VZ9luRoCFdPWzck0OW1a9bWwgbMBwNRSxd9hrJ2dTdv7j
LEaptprPpIVJQYnjlnOVBkJPu62StltXU21O/d60Xv5E/6KUocd+9mAhz/OBcqxg005P+fAFafpN
vb224PIKmcDSO2NesaLb+qmt42ZbWH2dDLlR8GQYxhrdbakVu9whC2rWB1mVWY3Yrh0Hwq8foxyo
bV7Mxm8BBAxND6QyNLPMlz5fJtOxoSxhgwotVOwjrhsJ+Ns1IOwDwD0vPBDmFGkMkK3yMhnI0QoW
llNXxVhDLg3L18dKCrmoCsK+dwlGVsNjymhQJwZ1Z5J0ZVUeaW5CNmx5AYuX0Cj05gyf4fOR2KXT
MVNU9lMZRkG+X6/vP5CIGmjhOSaDoaopS2BYurXtSKO1yrE7VCSvOrqTnTAtXxAXq+sRbH3zf3VD
xJDXUTBMcshvElan3/BIQpOENBPkgyX33rXxpPOgrbJtFkJycJnZuTmYSB6cy+lNxz5j4Xs0+o8T
MWQB1oaz3PzOAxDz27wPEGKNIymvKzYKGKmY6y/Z0lQRbMpGkYq1ToqXEfA9YiZBNC0za2G3uYKk
4otRF3V7020p94zVwCMBxl0d/s70MZwmxe/FDY27/iYp5z3kc4THt6rBjqlJyIWXQVcn+1P07j3R
ZejTcT6d7McNnaKiwhNsaINk2qko2zgvsvBD2kz2SJO9oXZXoyvlQAK+DGhB0EYFYfIx7xUNnSpq
H+YqyccPh/N8xLwCFcT1n42Rwdiq6EJ+hVaZrfAZGwRSX8dwZRNv9MyxwOjLJ8S0lWnyFLtQRVs+
LIq3eIhPD00FCguq4h+bOQSDtvG4XVj3uygcecNMk2AEPz4i/BSMI09jmbcgr7f/TPSdywxDJ/E1
lkqBfpue4s9iRJMK/h8S4//SBSB00/KqR4aZKmtXVfsya0lzTX2CbNaNih7O16WVWprgKV+H2ZT4
MEoRzIKxXBWT0+2E18cfhp3iPYrpe/FzSRiFw76Wl2ip28kQ+5bnrKDEOKjsKhvBiwpnVBveUkQG
hkFYN9UxnRZEioVGiL64EXxT16g30KyxBw+8Z3p3WbHo2g1Q2piDm08J+0WYUN7bdf7wmng8GJPQ
NdReENrGsBDp12d5TQYhTh+vOlCUToKTvgEZhrfNMmNJEynNIvqTW8vgIhMy4gS62xVL4hcgdPfS
/zdWuVd/NQQkxBQqdYPdzcvC6OLoryojlQ7C0viS4hazz0siPYh8ZV3HxXr3UQwYfXnQ1J+/N62y
BCWdn1F27yJIfcsOff956wf4OS57p5YvMAdrV1vhJIVVSTmE11ISPvEeyX9jq939chUReVRg7Xlv
5rEu9P9/vxtT1muSYMCU9kkSJ7h7ZP6iqPVuqyzvpYTewB41hsN5UnFZmp3JDUeTD9ZCWolorUAm
yDhdHUUJk8/pQPo91d+M4Bl9x+bdv85rzk2VtUIRHV7Q2RDpmhMKXUjKbNZXCd4UWP2zClsnyVqe
tZ4DS79xqfVa3BEVffk5mTNL2iqESgV5BltuOm+QHdu1MqEZUwzNBZHkrB2kpHzQq/9OWaFAH9yE
8uJ7GdfEnx1OZJCO1dQQKJ3yO6C3D49t/rDksPhKoj7g4wXMT+rNK/FbS0QebYh9qGGBLqjb1FX3
k6k76javBKkJ/C4+Ioe+JHXHaIEKCi02KPD92Jy8jzzCLjSF9V9Z107MnMKXHl5TV3AwBxGFnx8S
LOPlCuadUyX+lEq8oXVlpEzSCCdy31LMn5nzcP854CXDbNQT/rf0694XC0iQBhoSg5xuf8uDF3H1
6za0gFJVwHe1wxMgxRRCdpFpglyY2GIOsdVYIY2gTdczbyui608rCYVBr0/j/3NO7ipvWDRA9/eT
yDvFBNNN3uxKSsyJenLk3dfemXxkheWI6xRxGhYFEX28lSo1uTGJZvn6hPlK49WSvwOBbCZtHNTo
I0Je3Dsw711BICatYL1SVz8e2a6S0rRmHwg71V8HXdrhgod38URGsLa50YV8SvHN6GKgoynO4L9R
GcdXj2W6hVB+EooUOBJWzxXFgeIPbkQRF0A+U6X3i/Q3Y/x3ovZJ0OEZT6MOC55kEyp82IOxIM97
Vqma/eYyaIml2c8y3XdPv/g48gaMpW9bLHwsN8auCI9nClF8LwHfrk7ZiQ3d5PhU8tFmLzCHhRYa
lDB+tCh7fphJCVDxkay7ZAw6QCcmJQjT3GR9/aQQgrjRT1XXuDpyU+eKVkWNkpr2e8kR1GZRMiFB
+oMr51UxztCQiJAS3JF+jKL8VEkOtZFLa6+mT5hthYldGl/Bd4lhNUmHVR+kbIVZErGsU16Hz4r+
03eIzeyuTCvlW2+3MZ9oe+a9voOSdsjizycppgkX3xaz9pwlV5S8HZ1rP6UjN6L8zHM5/tPIMwni
WocoWrzmiTfNUnhud6ZL/lHUo0sv0cD/ISdEp5A2FamPgpQK0LX3vYniZSRHKp53nKxnnkxChSxQ
nrHRYnMSw4qE9p5ck5/gbuF+LtW0TOdQcPjMcIQjcRAOKDykH1P+GaV/dqBonSqZGbIJHxIDuTgr
dgyU5Ak4/yAs320PUI4B2r1bQk0jMLc/fpPR3lg9FO53T5S0X4v7DMtkBl3m7QfOxJ2vwUN8LMcD
vL0H/KaWYnyxeKhFZbcg5WrJ0iTRpq8vvBiMQ/Ct2IzfO8VRf7kNIl1KEJYB3caXH81TehVLTHOO
ZnHUSG0w5YTKhnz/BC3Y4d1fz3P3a+2GIc5PQMnyA0ZzXcEoS/7sPVA1gpCyX9BzeG0nYkm6AJvz
M3qy6WLq4Un98jwGSODqRAYh2YuOEdj11ukfo//hVfr5GcGtU257O7oyAsqftczc3MixGdeZqCYb
qG6RDVFPCMuarRG4mH4VkwE7+5xjK67JqzS4xTcbCk29+Xd3kLPLblOp3Cufcxo+20NAMy095sKe
l/aopGbOAn+IDfgEqBsRR1ClVv8Kgk6Ed6xoP7HcYUM2fgX0p1AV5TIMzOSidtYW6EhWGWCOe0hu
1gB7YOsGypKAAYlit3CdRNnPfhKQ0ok6weq+JiXcuwoX08uwIX5yuDLO35M3KSX16MU7exf0QGQC
YBZsGzjQeizv8Lk97qi/hYU2okAMPFtbG8DqltmslXf0CTD9AYJtjuVGkFVSKHhc4KWQXcTTgyTK
J17JBx2c5YKvfMeLxATo+7InvQNXU9FrgXIfg3V0dPUguNf01f/84UpWhv3sbxz2i0chSDtZOkQX
TueaYHeryy9AxXmqB6+N1O9E6TOgch7plzQmnQuNpkPgEyVKH6Uwg5PlpzTM1EoZmUAYRLRhVHRk
oQfCjKkRsIqHjX1rzmLWfM0KujU++8GSF+T3Ed3CvNcudwR/Xm6H46vdcBmlQ9c0sQFkqBb2p0Zc
9mcbw+K/Yqb5ODYpx1Rpb8l74belvAMzNI4/Dd88JIvpnqQHfKGtR+B3KDI/A5WIRfAvH5UkfTpu
1GuhY+v/5QiiQVcfx6O+NlQivsnMtkZaH15iynqRjfhP1wpdwP5wNGMSrEdI9wsxYn8rZGeyVacv
3CuZp8hZh5p3nwxqfqjS7WIZCXnzgfZT1AhoF0ecNZWPtnqcYiTDV1YIuaiUWniiOanGFY88x4Rr
OVLBbqwPXpomHqNk+i/MmVNEW6VTsu3fkDgnK2DEKhuX5QMPRIs9nfCA4HNCZO1TP8YPxZvYPdYs
wLor57RRwgZ6nmDpFmUYlofywqAt4vGzcfIXoyGMjEJn0OQsWhG8QmbjE/d6EPG8ho9yMSvHBApM
9/078EkIrCRe8YXiZZI9U/VzXjyzgFEE/wYmOvETmSQ/cbPlZUDKEQMDzEtbHiHjIXGvUkr9eMZc
LzBJ4Agu0kqP4+Aj2Xt6eBi+KTh7MfMX0zS/ekFNx4ivv1GgkJz3mFPxcxWTQ9hxbBbd4R/hsuW+
Vz3gPoyyGytDaEeBCFGG7uPYFI4oku6kiMQw08+GS+aYNE4BSeeT51qJvzMO6Hdz0EpFUk1SNO7W
aUZl21kDLamxFrsFTI1jnmh+srbsLpxi5yfbqy6iz+uWzssUF/8roSFHKl7puwlwboLL1+r7MzBj
a9W6JnU5xhEuRB0zeHnnPCoQ7mpehYQFlDkumMSzbPIbr6SlJbcCnyvmhCSHaiTPfiMd8zEANP3Z
VBqfd5S1I4lL8WXWmU4COrxKVbREl/4q9Q8ZAqJwlt35Rsd+yQKtcygTcu6he4Be3Jo4oYZDllFY
fx6aFU9ifVZHENJVVgYr6sGhX2WD2CaRBTgAq9Cc326BI1ScyZYRwl9TE5JA/UuDlnqEkAhX2/Up
Cd2PMuJowhnfTGtD1tF9QqIndTT61i6gTe1rMadnijiwaY49YzUHaSVxSewzCdxxYSM3HVHPXgXx
IOBkBrQ3EGmgNkOpdYcQwG0SHeoR6lpYHAO3nGgHz9RBDoUEF2CjLviwKfe+TtoJRCH+tiX0/ffI
yahHPxekjiCnkd/VImMOdA1w7cHqHm51VkFbV2nLQjsWTTa3tUKDKlStWIKgV50CzH/kzbmCFfpL
wXBt6Ay9gVdOb8FJE3tNZz9nMrKCCDN17bEDTCriSqYiVcGPxkzydzTWCVNm6I3fPOIafGtBEgFO
aZdVGLLSJISaj2OTQdHe1eAoR0k2qL7EUCCXaTzidINOd8FSYRzvAzVy3vbpA+5zR/OWN/7ms4ne
z1THucaxJUUzusLWBoZUteKsLeC++FDc/LhnSrQnQEzrU6PSGOc2afxVnvJ/gBMRjxzaqFQwulh5
g4TkziXqs+KRcmfO+NteGDoT3va8u0tPfLxwQhmjoIBDK3LiMXhOdwnvQRdzL5GEv2XwraEd7619
VKDstCrrXBsj7bNYN1DhNmgpzu9RsAWiZt65DYsp4JUcwnsZe9jC2rxDt6/7lStEia7/DHAqUIpO
eMt5oDBOAA0Ev+aHHmd5ysiFNxoej2KHtdzvCddDNRXwKNnXyA5lTuIxW90T1W9aEuTpv4jIPHXX
q+R8C0Y+z2IUjTjXs/5cDm4P6MZB2Ru2fYFOWjtnrPaI+zVlnOR9wYbNOOp+Kh91+cBW06pKvirn
2fuzOhWa/sGKSJkvECNzhnScgiS8WbTn19grwTW6zpbX8J0IG2HJx/8pNZcenj9KbQx/OJ4iqnCZ
CarmyF9+R4uVJCIVIn1hMLA9wgSng1i+gsu3Y09yKIfsmTRlMGcFFwTa3ai0CH+kbr4Qp8qh6ihx
4Z1ERtFzoiTP4XrC0513I2r8ZGl1yvkimiUZEBx9Q5iN7SaheQKwjw55d/9x7+3QlNteKTTRVDhb
gSs9lK78dIcA7v+M/eXCA1jutZMWmhxp6dIeMgrUuIt03Big2xNNe4Bhhn91Qv0sv5ymmrEthGfm
n1Ce94KWgBPbN8PbBJfybWVxEl/j2b8YhfhnfEtSAPWiO+eofq6bP2T+yh+0q3jWt2y3gXQX3rYK
YU7tuNQ8RjEKV1erbltd8sv1aVc6cLWyHr7H0WGM/a592AKiYXcCHxLJhHmWK+96B1slPeWAmr/3
FPSjV2oCtgrga5KCqNZLibsD9sdqRRkwiJ3hQsriQfUEP06EU9WLTh5sy+yh+PSFQB6G4YFYdta1
S4H033imnqEXZvZgtKoB4zraz4WHHC5jQYPbCAvMnsq1d2DIf3tR2fcYXat/LMYSqsYn9/4KipBQ
Qz8PdiaO0jID/NIGaEnPW0YoYbq3oxbtgj5GbxPeu15lOPlM3y+RyIuF5dW81OVig787EDPjFTPM
ErjjEhQ14SeaFn03tRuhrKankw/XUmwvYYsMxhCPjfH7iRzv7kVeTAS/ckB/smf/43i0zZHjgZpl
bJFQSxkDuvQguOEmocNP2ZqZE87U0TVu6SxG3gVkRQpUpu+xj156O0TLCnWdJZybjntzGo8bLPpP
6j3NbYPl6QdpNIm9egt3vuQ09o1Oq4GL8Oz+JWqQjmBZmad7vMUieTtlIwoQrDPgopHnDSqp++l4
RU8hC6x7XnJ7ssQlbwaLRlU8TzJiNVItNJVZdXBUQho44SFxAa+gK11w8h64kfQMH2FDCMVmLc0O
lrx6VqLaisTurEuAaLaWCXrmkAGYTcjichH+/jPetg1NAsVlIP+Bdt/Mo9Bk9LkcKar89SYJDHJD
19TOBCkym3qdnbqpXq8Tj1LN/rv7pnDp6XAQ5idOA2lwb7uNg0JWYCONvEy5EQb2e6Fzy/GIfbjM
LfNbOseWB8ai/+w5YAzW9vUj8/QVNxs2dn8b2pNtsPwcqQKn8y3lUm7FS6eWMZrBHuOn2622QESz
zMa7HmrazvMfJPylmvCgSvbzT0s9TAVxsbFXGIIuix+LBgsxqMt3UWXzjw/vgYHw6lUIhgp2JvJj
wImmJIkbD5Gn9rR70VAuPOR2oUbw35W/7TRvmfObLQpVm9gVUcWLdeZWUs+fnzoX1Ea20l1yx2dJ
MfoZPazlrbE9JJ9Oafloh06SrX+l4sFLoYNbAlXhYLTmFf1EuBgbw7FQ76Jpu+H4Caf2aBUsXIFI
SDqdwfj8cqMm0+xBjk6pFL6XwPzfrZEf7yfomAKs/tJ9LArzP2LLLDBRcE4icxMfWQhkOmdx7be1
oRhw+SkrYWhL8Lg4E/aVWoqYMi3ZJncyHxYXdWKbXQQXmP7KmjInYV7JBKiObVpw8Cm7v/Euxb+V
Bp9YYymFKuNclbSNE7BSpa9UbsO8pvQxQrsLEy1RlCwgdjxvafT4v42c1LCy4y+VMGBLtxFLygFN
tXn4sg4HgzjtLGJzBoGG7TqADnEnwihDe3yE1xjXv4Ab22VtgRfxOuJwgUeWPPpKTJ1V+ddlCpcR
WXv8fnWgNIXdWfGqyO6K/HDF0KrTAExPr6w/yAwuYqElveH0Cjf/dpvPO3wyKnzNGQLsxMqV9NgW
jKh+miyL7LvoggOFOPI4ZJOVcKH7SH7m96muRgySqLixOruo1g4Lik9QmwPj4s4h6Y3RQTVNUqAv
otoq1WSkuCEan3+gZlplpt5+VjCckWm+Xmf9oH8nYYwUsJflA8gs5qDIvAKjL2nmsfBu0DOYw850
zW6xtMlngYM0g3IZiTj/BWnlOehXECD1MTVZVQ9lPKrDYROSx1eeNKH4vJGdUR5Pzw4SQctw0Zu+
a1uBq4wYPfdWlpPAyiTLWcVkDBzaUGgVq8dxPZACdH1ItMnpxxBNPU0+2qAZ9d7f9ZMvblD8YqqN
vJyve3EzhCDy8MjxO58G+TTdsdaEDU3E17juvmshrMHFv32qx5mm/zvxNzN6CaL1IKMtQL64AgV6
Fjog6TMhefe/QLtdH2Vkyxi472Ge9WSSKQd+esNiBsryiiiBlpYQIxwT0m1m/azAWUdlaMTg2CNi
VkNkFVVMPhU/RNfyhY7IeYvEfsSEpSbw7kQM1btj+RFPTVYRtpB+B16ZO4TPiR9O7ZUl8H/NH4bo
e1HrpTDUUNEl9bZFwq1z9mQ4ppUR1gd82zVpFNIK0CFLih1EsevWimtURBzBo/havNZB8N0/mIi6
aa5NFbDFobG1v292GUJ/yEkxyu4xOSB4QoSGGPvB11sam9eO8L62AzuQSzQX/jQZq3wFYEYwJ3gC
3KTyG3ea+wGl8y7Tn2024VBI+0NsF7KEMN4oXMXz96NeBPJF3uZZgdNHWscS3YjX/EcdAA5s5Cu8
6lTIAuD2NLWrKxw6kstVSxWAGqznYyyPa6+g7Z6QD90h2pC7O/1LvjwoXVGrqif9GN4AlW0mpHKj
UPrnX796GoZSckjrib/WlWPLzAxc8IlhTKvFI47xTHlbw0ve+1CkcBCscuM//AW27QQcP3bxv3uw
uqrSeNiVYYUmUjG5dQ03Gw/YGMoX1LYaLO/UT6ohkiwj8ZP6wKa+cXsbS9rkvFQfBI2XZ7wTHEri
DvgfSalELGVgfKM+hKnrFMnTP8MmEmHZ/Ntz+9RrpgTTvDceFi9c3srHR9jdGnaTyorDfpnkmMv6
d1ALw45IB3AN7LJs9FImO+YYhXQ82bhJCoskI66fhLpB3tYsXrlJJF82GsBs6pjizfb1PHA4bvEW
mN/TirT5en8ui/E05JkzQ8PLuwRLCT2Z1fE5bLimBsqUlI4oQQJozWo9NHPV09fNxWfMSUBRzxSH
zAjpAUoOzAyIkRiJyFpOafapo7pHVE4hhpdpLIeEsOWpwIHPWM23m80r7JlOs5dYT8AdvHuDnM6r
pEw7a3xYehGIutKvh1gt7euxbuwKKDHKwY3/to5rqfeEksepmF3vykk9Wonv0Reh+5WbZpy9RzuS
j6RIq8J2EwjOKPhaFV86IGhkQm3SiE65+oWphQiDuxBaW9qwjXVPHFd+cmFNPeIZg0vaszP4fuTF
e3Bc+6Q3iu4EhuyeMQyHSNYLQY17WsWMS5vUKYvf8gG5d3Wmq304b8skmj1FJAOC80HjugJtI1nk
Eud+Yygr5NzRR83BOfoDsj7+O50aaiO5szh4YeQ8WzEjlL0OQqfw1NL8L3I+AVshRoQwGwgn0Kil
+7m0E8+aHn1+X9tzKp4R1Hk4TiouazOB4xEUiYgMN698zNPpTrWL7OYbr+tftHP0bdXyclcZ6YVw
pL78rB3UPpJoe5QiXFVYmVBhdSERMzZLEHe7Va6pdyLCckMYgxgpxyrl2ipmEwpX//1MWIF8VIpf
yXt0VAIZjqlA6JxE9QsdSARLGiP8lZWgtT/iWlwSanGba6yz4KPtRijddxwHnq71AoNqI4Q7KZs4
8qHFF4uzq4hfM5S8Budf6YprUuia+aCSAa5Yywwq1FWhIzBSViUGWnficfi+6ByUVvUm0+1T27CW
KO81uyjO9nJ3PCQ2cl//hkVYpVWfzfGxDZDf6fc3TjzRkSXMvm4B0F0jCCYaK9GI8z8fPvnlh7h/
WyZs/8zxbxCAoVT0F+SoJRPYm1SpDxVmipHZXgEXZmTaOkIcS2xp2uVuTUEvD9/kuMXCHE4ef03A
DBSoF6cLHWJHhYgASy4cUzO46LELcBxIU23O8ujrEGa5kmuRyuo1Fw95poKeGacm6Rw1wzeEz88W
7NDoXRH3/MgJdJY5KFmD2+q3ClbclLmOOcccODlJvqhe/6GH8O8XDQRfY1utEF2DB1qpqQOPbyn7
KvVq2e9GoOLH9snBycz7DS7ixG0cjCTbeM5B7nMZF3voFHQRP4/uFea9kpln2ouXEsrJvZv+Hxcy
7vvh2brOXuUMq/qXQ3qjz+3djALmk+jXnVhBawkZ5VpiNQxNrv5g+h97gsJ5A9D+QUu1BW8cF2xK
LPzOrrzJ8DYG8Z1fEqiAXZZBQA4itX7i5Mh5QVu2HvL1NYIWpavn8QoP3KiY8DY53KTkM5IbOGkY
JPo1ZZ5Y69Z/+5Y93XkT96TFFniJkOs6hA0kO5Hmy/EEDAlVak6Piv6oI4L4Lh5Dq0hOYPSXwXt6
H23aPJTaSY9rR2bul3A+xC9d2r3EPLg6uPHt9V2lz8FmSELywtO3LqZ0xCRKsC7Vurkx/0OQZ9au
Ca0SDG/ikESmidMbisiddJ/DnYTiNl2Nf62F3VmwbJRZH7Hg587LTjBGSZUZoJ4ucCynkVeotROu
dkwh7lwlVhRD6mSXNftqwPOk7lB1Ki7jzMH2FsWzYJWmb07ENIIp+RBYRy591mFz0hnnyBPP87l4
K8wT77lnIrVX9elwO1l0yfyUw4v8906Bk1QjwZ6yG7up//AJ3MDnmZR/mZehgKCYyXMP3i+q3j+E
4x0suSfMBKtJ8RDW9nK8t9dbQZxyw5A/LLKYhSG+cy70AxdXaO1a7UA8qAnM4LrswJraG7kIpucN
W8qdXmKGqbmv4Mf7Nb6x1NOl7nmaUuSypDKh2ytnHL7g/oguqSQLxlPtxl7P0m9A3on8CgxfTDqB
L2jY/2dnm2zhvdC37FK6QdTn47z0HnDDZxJ8Vf0dkYJYaBCrqobb/8n2CphTxBm//hmhN6m+Kp+R
d2Euh/bhCpETHk023LC9yqhRNAnXCnD8Z9c5iHBxtUUOK4XU64Q9zmR6tqv9CU7lVPzdF2Py/e3n
Rb942rz6MWBUwar4T2mC2P8iWsCmhmbeW+4CR+mzJBAtoj4urclz/pkPL9HCMa9hgIQS2YKKTqjo
jmTL4nha/Coa9d8TPuWcDU1qx9GpY1VR9PQ5ryc8Clb+7Jp9qxx/EbvS84WcU0BXEL723fHvsDqu
9YBv2EgHaw1vKXE9BfjdvQXLUw7LbAWjzjmqpnNN5pyO7yiUpbeot2S+H4l2HBSiCHy2g17lKz/b
QXqTM80Z9EIJMNNNUL/cws3EITLXyUQPFnkIBW9iFEVMHpjQ7SA2RM8z6wuPXBHb3Q+M42T7BSQB
wWA0umLf71BLSZPGjvPH54MNp76XJDl5/BRHA40y4NtB8WCRcFNmZ57P77cv6zIwcM+kjKBn4/ne
WgD+3ljSf/fHgtiEaMFyRUzaUmQpqBODIqM8D3mKYl9GOgq5JkJo5y98bfOzqeTZH+Q3XDgnrt4A
7xQf4BzV6ODSe9Zp7CZ/2PSbaCKG3UbKr1GY7bSx/rShOzbW/8MKM5Y6IIonDz2OLOJSevcSZrvH
9RdpacZcDoNI7sd59wx8QPaF/TJHTQc2IYgKpanDxGLSyAeC3jg6RlyKICUrKvC/bJrGuPLauDH4
MIGTAWM5SZBzpPCR/1islkQXtDhiaa2hxmfwAB2zY/Y4JCDN4iXR+JfOjGPbFBqxMthI2TLMrq7D
ZVGM6RK2jwoAyf89eEHPDxvmtyklYMwbGFytYg1tTDmYwIs0sYNvJVH81tGvLVmESP9+06N4xwiq
iByw/VeutRyaEJTPEIEVKHgxY5nDPoxwb9sxEZEO1dvorcdsI9StPYlZzeQUb4kF4RLM2OmIiPZ0
4fEWuEcDLg8hp6wwcBtdozRt9vRz/tJEamklAui3A/lx2En/1U2umcQ9fOM+JgnkBABLQDMqAWa6
BLAp32ToZr5kU0tbKzc4GYzUHORv0j0hV6XlsrGH679UJE/5+Ky6pUaqbekU/pexExm5mM6cLMSA
wy8rA+fiD9JntC7+LXw5NuK875/m4351++cTq/p5Gx5Jl8jVl9IoW1iDJ1HpECf2TQA8JR2J173X
BHWD61E3zKvh4S4uJE+yf+F4BTQySQXwmzeg4c/nmv95+crqfvVsjlghyHo+UfvamC7Jq1LO/Xcb
UgRrNtLMTakWD5T6mDmxAC8zw+Oks3qBwwo07lNpt0dw2ddzpai2QyhrFf+qyp+xtaGwz8vcG6tR
fNMVINJ1T+nH94tKnX66CPNfQztuP07W4DwT45CtsNqCwXLIQVrpSj7C604qoZfXV+40sDKRAOq7
GA7aB86NEoqBauORTroWEUWnRrIsQLh1zK+vaZ3LQFhLYqHsaxA2oobkAYv1xtNBDjKo9qvp/SzT
ppdJqkZcicuiqcIgY7TXj9A63Zlb7aKnVu3DQXAb3wvYnN+uVrtdxYmkZf4qNRnMdnqcJql7OGvL
+ikYd0I0QhXYdRcYYg1Vjt+RwO4DSLKrrDyDYODYt3WkOXWzO7end0iTge7OzCiYndlcbVTdG5GT
fMtFNvXIsdHxlAfjtw2lCvxZRV2gbzTJuetP02DBzMDs+B+lCiihz0bynF1b1TSbr119BOKD4ADi
lcrBA72+EPiF+1WYy8ZVkvW5SFr66ye+VspRlFUSz+zZIdgKrMUoRRsgvKEnXWlYYFHYJCe/qdOz
PUIcBe3ZUr/XiDutJ37+/aJZStZEuc1aUWiquv03Rvn0d0Y1MbzBXuA3QRNfJ2Rry9JyzO8/Oai5
OqXDH9rbVMYuB8AysArAYwsyyV4SgIGC2TlGxz2qweqblhC5fSq5j9Tyqo+WOjdDEyshjKnHdfYs
bHqa6dK4FYEZqVAdp335JhcADOcZ6i8QOFZAEfQMWl4e5h/NCfFa09gjT6udpJZZdHhZULzJuJUD
sYUts+qCG/NEi+VCnv5j0AEqs8Ec8dkQouUSCrgnkkZoyA3g9GCHRGVDII1CvNUDZwVcLNG2cBh7
FfPjvZtXo0eLzBDfBrtt8j//nvYOOFdl8IidNiQJxpuJetalqtYF9bPqA5VKoSzJ/hj9HqnFx5NY
nBc6eZx28rZLQ7eTSfZ4BbbZAtIMbvsltGrGG7PScNy12zbJZyqRBd2la2+Q1jCthIYfjT6EuzS2
Ixp0k+NDXIXmc95ziIzxV0ZdAlWpVGdR6Bm4UInd2c72ZMb//QORhCx2srfFWRHAqksmdvOolly4
BCz9l8PDEmMYwTEsMijwHehU38r34jUgJv25xkIzVKucdB22iqFpHlJzsKtIwhsvSPSQulkgCe+Q
vw/4giEMk8gAY27wPfo1RkvAWdCwR5bC2V3if3vaDXi/aymM9HjLJcZAY/dSXqJovsvRWvR92hgg
/jAYDmPRGvN3iVxw7Ft6XAL5u6FTyNSB4SvvMNm8yF2XLbFYcCx9SK+CnEzJ89J3bYYezeVTBTvz
9Se5LhQSAyS6gqG2BsiJncLnNhSG2D8EvQAhkiBfmUwXcxr8FbaHFLvArkAkcIL2VAxSQ7wUMWUY
0eHndT8A6/YUlEO0+Dxpva9JimevnVK6jw6EPYS5J396ra6dVwAm4wSu6BC/D9Q+zk0VSK63CwBo
YGFqPwb9OdTV5N7iMXzkUI5wX5frC0gL/CfH74JiRRQJotpi/z+y6U6DOK4Mt6t4uY8RcwpKAYki
iG4HWdq5+UsCEKO92Buq3aym9OGclRIkY1R6aolgBX8Ut6SEt89lgHMsvYfQLB5fGwOsT7ql7REE
/kRRHbu9kImLKs4Pbf4lpA6VjwMbP9iIjqJ8lOPi1J/bN+5iGjzmrfUpZSmFtzTOF4QN4QlTxsJ+
HPEL/qwh0VvvdzzS2uJcGke82PPAXRih7X/wvBz8TmtaMkzELzy5w1tsKZzg/c8sQNZF8gH+SnEk
thID8KqP+iIdejIv/OCdTETjjxSUMacMYYMzqJW0vVfDvCD1CmmtFSbzOsRV+J15cxkDYwXS+gFj
E1qghq4En0xphLPsVfQoveI0nWjFYqkLOHIBGGAVAcu9fNa/zg8w7B8XnvdTaowtuUtUaDUuVwVV
784alLjr2lWTtM8LTiIu/fci4KoXlQsnEPTmFLvZnrfvG0G+o00KQEud2Dqgbk1b4ilkEXOmyCZE
Flil/pXJiXPW4rgAV5aF2zxA3z5E6zqNtoAumUOz/+XK6EzUrzQ0yZSBZ09E0W3NfDPWNAb/LLop
LVz/EXTinJ8NGKTDB5pxYAsRkrI5LVvE3842AocVfeanIRxnSVM6PVyKQjD+fzkJ0KRteAs0dD9O
xAoXgAcCRRmcdwtSoE/q4JW06RfNkVHZIrRAnNFdt/BIJ/NjeS05Y5G0kZps6vpSlzmsb2iXLcxE
0vYoXgsfyJCSJwENk6Kw+pS14eVVrU0g8o21oywTGVd4t+Oq7pWC6RiY0O8J5NiKLW57D4LTjdJ/
XvgbK2g67jlXku1yiGMA1c2YltF/Pp+EVuaXHydZKt2ZqvsnyPlKEtV71OvHEnVZEJ2uFHmDIuZP
h1kZlTaYUg5hb1QfX8+zlcv6xJYSMAVfJQDypKIfu69PNQ2NW7of6ejVYfYVcCfPvE/3qQrQEiL8
uWlFN583arYskVC2WIbKJgxUyF6JdgbELldXR4orfbKUFDBc4Nr9vdpNi+amIwYIXP8/ZymT9hcq
gI6GXlFPYY3x7RJW7ueF11aXXTRnQUn00G4CuLS6umSxus50yI+8cFmV/+DRuQHnNna0BTCGTN0B
/EoKU8uLGs/1bVFQmD5O8oiZWrrHBSBZK+xZ7/zI6vtikKltQqfRjcCJTKy5tMSEo7TJor3uHQsj
CnFgN0u6GmEU7JkxDKQz8Qqmweq6BCgyNarIK1gAES4qJijN1T5dfkonHPTPZlXBEdnhQA85tKQX
0uDQIKwLWMA1ZyrCaoaTHHLEAoEDwH+nF5EynnPLbWPCjIoa5YjEpirdiHY2P6kRSUmYzn34q8lp
WkozCpQ+at1JAY1K8KLNIHYanobhUh9TgqOB56O0vs123tc/p14oAk47HgmFeP9BBPNr920QNhMF
BIhbbl3pabwT91xT/vz9UA7HP498TfWi677/P5vFXBynbz011rSEY6YLiaayrRTC6IkXgw039kPk
5qyJSybRuS84Ho1d801q7dXaf8M1orB3bzksAZDI7tKjez1viQ4I6zX+4znLpokd9JNkmaoQKzMT
ZX1xU1d8cZIlIQHOvuEBciGCDhxZHob30kbdo5uwqMEWpgiUWLzOMcyS2l1P3qzkROm1FqWI687I
Xp7D1knM2l10utuo5qErezjemxZHChFwXz5BoYEboN0IkA/VSdtPmuj3F3eXB+UaeLG7/NSr+n7t
jk/CYEvrQMVJrbKOL6BSkDSm8xC+f7pHZcCsvcqthn3MMSIO3m1ZL9HYsadupb1t2Dbh9Q6+BSKT
ejTD0eFlfF80L8mwdkGHzy35fzIZ2YsDkxDNDxwTMaKtu29SbVzyXj25EN2D3ranqRvYv5CV+gEF
EdoBGUCkeHwCjtr7cUUFsvEvqgmgL7MLIEI0yTcJICPCoRMEETHKkGiGixzirxU2PVI0wvkiphSz
0Qf0np/Rc8ltAYQ+TBaf5mBRumGkWsX1Oo093Ltl28PrMRZ2Z5pzVoZTtLnoMiN+2B4BpndIcpbw
ZBefgnDm0FEsn3mNjpvNXufWhKmTUJjqzzKgKs6DKbojyBTVazYDvO3SONi6gVhKrkvPpIF6htkg
wvXDI2iF5tufw3F6mE1Vg1X0ZzPfHRq9FeCIVA/ohg60f3vi8yf5NLY415oFhD2isOsK+jQjFAGW
jhnke5QP+cyCvt22l4/SdfL4Ob91RLPW1XiljgXvp0y0aFUCiq5PaQXqhUB294MotNYam33PkxOL
GKA1GNSwCa7WMN/lNBDKMjMm7MPKPSIYWsHDF92IS6+9lzq/IPsnsK7hGw9tZ1axAPoCou3WHZLC
9xQv4nicjyWOiLr5bR3AoDa25f4PoHqCAvS1u+zm5q2nbVkZ6F6jRU5brbXWIsJ1J7C8DbVKVfZ8
yAUc+1irxXOrNOIjZmNgMHCqnUiaz0cYMGPXXm2sBSwiAwmbEVd0KFqvYzJO4Iu0+slEhe2SoU+G
qxVLtvTjBQDVZriq2rcJO2Rll8a8CTVFuMF51OiZFelVDL5idSjVlLVAJynI9SQONrgJ+oh3im1s
dDdHqAobSA//cLiFaOFX+TgA/6x5+b1iBAapZWZMqKegtD3hOhCf6OFLI9bDg7GGle4wcn9oi2hh
RALGmvovrimG/MS6vpMo7hUpkTYr+DTZKTdmy4Y5D/OLBpgVZquEy6O9AEL5U7wvqsbCeAJUuRH8
MeZvKJvJObSSItM7xquxRvuvFmhsTl8LaH/7f+mrUy4gnLN1sK2EhrcBbJt31qVJecevzCcqNJTt
Wy6/NChzGNAe0CVn6qR6pN7wCfhqdIKSgSyCkthn2uHxtwWhUhE5yv8y4YqVdFRrdyJkF8odb5xa
BlqlvDY2xw98lv/jZCzJDOMebX3RUMjxiPM8y8LUOFutxXBVGhbQXQYW3xOrbdCeUAVozohzhlxc
p5aBTf/qYRb8VdUnBq8SdbGqx8vIVGWOpfV5asccKoAaDUzWEh1NEExzN2Dsxb5xgjEtQvTuIvJd
Tj3phMxqtDSgjCbClwren92r9Zo6iT7PWkZLaZIV9K4pvTPyD2KmsMHNKCRY2PkmDhyjX+gq2LIz
Cf4djbD8I0fb3UUHV7JBE2CEoqGA82ZZwV1sdKPRtP8a9UL+ZuEzSpX94q4MezlpI55o1q4Eh43B
NVXPK8bPX5Vq1THf1Dpk837CyxEetL3vrflQhvofWb5wTuE5eBkFhptamLWwaGWN105f5g2Bw0fe
DTWBubIDvWvEuuNYojBlzucILW0ITWpiyBFQlC2PU34eG4pmsDj5jx9GdgMu53lVVSddmM6bIUaI
0DrQQH3MeEfMkQgyAcunpa6XTG+8nk+9u8voOPjCTeapYt+pIh02J5j/8ib9npVegmj5MgQFlUW1
+Ax2bzZdgFlQrOouQ4AYFlwENPcVb2yYNo2DG1nj3J89sKNI/24LRLLfDz7FE/fO1m8j6Zak+gsP
sM1OTNZmD6dNTsS96yWHqvHa4p5BYkVgT9XJTJhYfyMwaB8udjfAel8rHqCXh5mGrcmI3Ri2st2B
UE1PdZv3gIp19+uv5vjGSeC83gEUTSI7lsfsNEJ6A+lnp//IRarLQfQrp5WsiB6FTiGkMHHnQrmO
ofMoRwTjeXCTRqQ0oy4CedM6De9K9hrCTZSBxGggX0qzl1rvkTcxBdgvR+PL85MOlBDCuhfNw/FJ
VUfBFqfRGl4j2D3UezkAC3S75AAfiaM4MTKBqVOcE5s+ejORNMATvMIVDsHpEFAusciwdFegs2ak
6Ia4MrrviKNAUh0Yg+1GO1Cs+b9VJvzVeYQpj6SdpKKcIHR8HLXe4iVGzgI6CUjhQJ69Zhncm4wf
eG5e0a2lmLx91m6xwsuCON+ubMzDzgQWkpmVaRv3Bp6AXKuCm9JQoGmEWo6jE2/tHI32/y88usyw
6U0hDo+JCEvpTaALJPmS5Ta1BTV0gbfDZdUpZ7kaPmmdKHwKxPEnXa2btVDarQDWbw95Ta8jkiFN
VPbd65/SiuDzxJ4Cnn09ryY8DFM9wk1SSjWqjmzUo5CTcgvmcDDkGjDfIoqPPFdm4ccqbvKERqXb
htpcpDfa4hOcKoxWK4o4aEYCteebARTQeS0ed0Pq1vo5mOE8hurOfYfwCxzK9vF6LduVbPsVXW7k
WB6iGmwi8iSKDKvNzHOZkw2nsDig5RzWdXz25t6V01SbJR7q+l6ne4tSlUUSR45w6sBTkE6D47Xd
KBUm4EjeZ67X3bXvZoqnadMrkcpKQpnhqnf/UWY3lzxoki0nKJze7gLY6wd8Re5uYRJzRztE7tsJ
CJBcHloyEX+svbVnNJiX/VNIqCXuUphJZl4PStxN97UntSkQE/uuJVaLwiHICwHYQ7Vg60ssFoOw
/eTkvV2RQTRi/G5qZNn6wdRWgE7JV/Csi4DI26PXp08bF7wmV2abjlEvEsBW8axGAGmVsN0StJgP
J+l6Mg8cWKkWRk5IO3a6fjLtqh4nI7+osW2yWaSmaJpu2D4LF9VDXM2TipaaRHl+czdcX5V2/6QS
9F8U+56sQzC7xtIWuL5lKIafraW7xRNLK1UJSxwIGVKTr8/nFoca6MwB8AqfW7rNIvsWi317U8O5
Wf+UGg8N69f+JuLS6pdxu++ie2LxxgX23IcmcN+xcApBx84XIxdvkt2RD4FuavI5YngoSazwDHJx
78JyDNKSa2ojIBOElggXcg0WIgABiSZp50iwULl+eopOl0ZiFFB1mfufOsPs2elkI4WOaEib59vh
ooXAHT7l2uJ6US6q20ua88gacQZILKLvehttJskI5GdcxaI3LCzzIsktmDEdDXOHc3o1TOVy/1TO
sn4RCSXHlxdn9vwhQQqr2X7936PnjzuCQobTSLTSIcStGH7iY4B3yr8Gw2cNXAtRYOcFj4NbpbHh
/p0jwuNoyZClwQOeTTErbONooIBzksnI8X7w0BGBbJ2f8n+AulwrJDFBLY5RBvS5CreWjQJXarEJ
NVtCMGHv8RNyusR7Z6Bt8MPRoTFQm0fIA45RQj488uTFGVLnfZWRMahdKPoH0dmxxVJQZeEwOsla
eDpXlLzpuHx4RUOPY9DMLKs/vcU5oEqjlYGQbjmESlXQVZX1RkuinTPBOFhvD9ZCaBkb7WYctKF0
ddPx/NHAPYxrGFd/v0mkAbQ3WG2d6B8h5XO1XrBJ1fJ1ODQM5dt7/ziuo9QRDe3fc1aGsRT4T2ln
guK1OAZI+AJVaSQDJSPQR13zQFNz/e1Z9cfKyIskiNvY2Np4+PbszkLO36Ar6Bj57fM/SqoUHtZn
CPqihf1DhP/BC13hEgOsRHygFdidcwFov6VGYG3CDOtizg2kSgzUunw/NMhn4YCcuc8OYKrZQCRI
AMqhkaAPmERoDcG69qXbHj7kHl/4SUvP+kOM4lTcbP7skwz5mOLxMpr4jucwe/U2Vb6bz1bNgeF/
iSBgoqJnADSgq0mxhhE3sysbc7Sp4z9VBkbo66n2i87aDxorqrlHDytzLNrqwK4uLCF+JPz8sZRc
cO4OJ7gQF/GXcfWvB6QuRWOS18v3s1r55Fe3iUwOTkNBNqe+2b+H1F6JBC1M4DM1RwUZZ1qRl0qf
bKUV5+OBOVM8PttrjYyS+zFPJw5VlGJqmN/u5X7FZaVV61b5MdUF1594JgoBzIFdGhpEkg1yu7sF
K1IyWZewAGHX3ewMjfBtkcC9s41Ecb7Hjz1IsX5f5A9krO8kO4t6o7+Lnrihc4QhUOoNtGr3nlxy
4syJVYDVakYrQC4v9wqp7YHVDQdj+kqtDGehulzLRF2QlJ3dSCawbWmRIoJt4NaHuxE6VieUEEBT
DOK7ODCL66r9cr3CkxWnHaBsBdlmGdJTGADCU9xNKp26oc5JpgxfE6uST5FkPUz7sfHmzScD3fbA
OICaB2hILfk5d8N8IY5wmvGcOhvf/W3zbSMZFDgz7bFE9f5W8MCpguUuzfoRjmHaPngKmLR8MNfi
8PqJCvLWgOUKxg+5ZYAEJyWzzwP1hDKXy6/C86MxtcAfcw9eZx93CjNMwyBL7kQ5erxfyCd39a9D
38vRLTu63d3RozMQ4VOq67cRTat/yvLMiVhLwMEsVAnw63yUslZZcqj1VFDNC7gN8IcC09W+U46U
1IH6GSC53ar1CZFmsZeelAW9E07QgamDHR+44X9FtvOZd7w3sMlLNdwsfkLrF54hNMQGAU0kjZaE
BXmH+SZjWq9RAKcCWlcWegeYAeG0c8ijPnRex9yh+dQqKGoZioW/jRF94Y8NBW2y9FL7G3Ks6ivB
vbcG6sd2iAQcbsinIfF6umWSNrE1RPdY5t9zvKaRJnOjb3RYKFlTDQ/zIc+2ZrHEsuftzNSjnfxt
+uxZr2/G+5ZdksxcK0ZKl3Zt/f6JxHkeHpYdadwDY6xQQur5S6NC2gmPpFoucie0H8NMVUcMrrz8
+1l6H4wF0ahh/pknT6pWzJis3MrwOfh8/cXGegJwF0Ya7rDh0KAcWna6nHpcgaAY7A6SwRApIWOO
/Y90WP0U7XHaacqoOkrIHmrhKyMMMz+/VM7to0TNi0hEIxBhGv3stNNqyhorqgwACFR7bPphD13X
Taitdb5hB+zO7nD25HCjFpa5P0LnmXFBpcwbcLyVBdhhiLKVIEAZ8ME9lTkDe3jD2h5jv7k9Hmpg
LFXw+yIhBevQjGP1jgRBhtWFxq4GY6UhDSC9+JkBFOzjy2ketHgQ7rOlVIyo3BGbxmuiuM2Tn1n1
+0+euDxS0LZQjTYdVoDaT7uRywg0ysUIk/qwYPrM/hJVTqnjCNLW4WYagDR4KYVJw7fqEMpbKddF
2fbA6Dogy9R8RNRbc0GUo638PgqGKiJXL0RVNMOBUfWNPHh17ut+xL9yNQHwSZF4gh8LaTcxG3gO
XVIwuUr2dJtiN8zy8ApSYTHoxLFw9wAd2+jhwIStIVJVHkgZiN4fYWpwFFFqGbeY6mE2skL6yk6y
CDuyaj7B+3gpZVxbHIq+57wrUWF71J8w2flmZZCBlmusaWMT6gSLV6Nfi5VkCQmFLNB5SyfBLx5g
pPaLat4+Ma9fziLnqxfnm/BaEiKtESGo997XDOqWAA4Ap0KHB3jT3oiyOhIaHHBvZmxf2EMPxpY+
pBL9TymvjkUuecXNkXHK+WyP/P77F25JwEQS/xHNCthWzKeomLhtD+y4xtT2CGam2JnVo1OF/RnB
P5kInPXe0FAevBhqbyqrgmgZLOXc+yrditpNsGEtOrR+V2Y7CAMKnD5mod/UpdxymUEp3szDGBDS
Pij4tVVXn60p0T9HiiMyHq7klYYZoFSlgl6Hasx0mR/8Qy07PDlA2vktBxbM/KQEYxa8JyaHQPFi
/3a4s1DyBfnPHyYGuWY+EwSlkyk8pR55hoq0+Xz+1KWqI/j+m9Yvc6KpAcizYNAb41ZRX//5Xc+B
pEEVJluz4V5BSVFuoXHk6Pnr/uDjq8wna5zeakiWdmihAPon3URmUz3nodVdVRt94ZZuK7OWSL/Y
Nf851Fv5l7qf9OO2sQ5ycyawjEDRMcSa52GMlpQlcSRAdKcusnzumz6kzUN13qJQQt3m4IYLC2ZQ
IRT/ppst631rU3Eb/jidOUBs/+dHlwqzpmeJlOqp6MPbB/bKZqWYRXy7jlfDMcS44AwMJ4rUJ40w
lWgq7uKaJOVklXtcBp5bPPLBNd0DBKdD2z98Amcj9pEoJK9lZBuhdgXG9b94Ae9VhD8Acb6O7aJu
vt4Xt3cz6A+OOU7QEhJvaD0XLMinTcTDKRI2hUEyll6sW1DOqVqG5LtBwd+xO1hz7nopeUmRAEmW
p7C/VzM73x/TnCZQBR7vzdTzmyJhRmnEjSSwgThFU0XeeyaQGt3wzAk3EfpzidUlj4kCdjIWh7Jz
f7FipQiraVjAtCWZN/77lfrUfJEzJWXuK7sx+Zb9BYUGFc6sCdsjrbDDksgBA1tfqkVD3cyZPS+/
S0R5TlHZBYIo2Vq7IKrLM88mZljcRLsC4PKR3FfAZwBwNTKIG1d+7RliIEJ9TKBUP8YSrpopMxIm
lv27pw9mJVpPnlwKuSf3Cik9lkgVCVzPsxeE6cHJX45ms+NzYyUbOBk1Z2ISMWpY1WK6J30z+ym5
8ptDPPvlrfa8FGTh1l7s1O8pbuSir90ZTeV/dW1fC4U4lkEa7p1ymOq/w99uIyyjSe+hZuZbOlhu
YjU/WlDyXLS3T4K/Wl2WEsA1UYLBzRgizsqK9KdwhApEfVtnKucdS1Aj4Vsee2zi0wN1ZzRQOrXc
11DNl8iq2KVrJ+sgCcaw3/iJsLAnMgoWbJfLbdQIQOuT242vo5R7PLgjYfojby5VK9UCJSZ7fW1c
0KTGpUooTQwRFhNpcLP3llCMSPxPIRj31cUFQohXEG+roGSuetqC1TR2roVxHiNE7QMp197EqVLY
HGuN+i769C7pT6X3qwdo6eBFhqypiD3iryfUBZIWuA0uhyc0XDYTHYlymq4sEzu3/efCI/BYgVwA
+xgQuuKYquJAs/aSsjzJMFpeIt/+2ZaprnmgL2RUQwQ9q8+gIqMxaP1zUI9xmMjH0rv8ix/Im4Se
MdqY8YUZCMTHCV+pN0RpAoY98S4/5NdXgf4OnooFK82ncfnFbdRGMOVu9KVg/KIWx4A77COHs8I3
4Z39otJsejprzzknIbL+KKb5VTmPmGGlYnNB6Jn/hX5Jih7+HeW4jkNMdlmn+MeBUzbUR0fW4vUG
PZkIfQqUkU6o/umxRdxlI4iaExgCH8dMec92O1K78WCx/ad5gRQNA9YbmZbuvMzY6KyzY/zzBHh9
1Ec9uxMTwfvhJjdUM16jNUpW654EhVHky9aSq+VLpnrQwPMWOjfD7xqy7Dfcwgd6hz37gMTll4Sa
jSDfnRzmJ1aBNK2t6RuYHrstG1zL09H/kn5yEFu+ypCzkrPHsJD2EFzmhjci4l0tvrwBdIsgSA1P
NmK2qGy/kV7WAoabEX2ghQY6irZQT3Y58llIPe5teDD9l0kFnetSq+DabprJOAMTvs+tV2uL3OKE
wqUbuwXXOiHmLSZ7Y0hB7zFCJU+lBpuJHGrf+0AckGCx0Zwt60kMJVjN8uid9XEkj0Lgpo6Jokq9
UDPxquBMd/wo5CXLMlf2bgdVK91cm8qVZTFyLKsa5V3ww4N2S9v41LLutnCwnv3BkdmDNr4kSnhT
F5D3IFaJRjcyMwsLPacSnYdUi1RMptml8gESYG3R87uO5IhJKC+repobOqCs8bSvq9nwqLcKCqek
wgganYkQ+5zc2CVMa54HAc4urCrrM07KwL4mlUK6Iqd9HZIBCZMGfLoAr+Hn6nP0jnxMG+31N30O
btpy+xYUm/87/ptcdWVtEHjlrW7NawamNycEvLcebsohb0ahXcKKM+HtLu+Z1QcBa461dLt5Ae4z
kO9iVQXFNYBCqs82BZlvacY0R1+i/denANy3hN9FiuT8uZrCXcxfagKa4DYXFbdyuc7t9QO0w4Xy
2qh822sQkhxRtBEuByDNrjvSA2Gw45IjhHgas86ef/hzq/D5ibhHT1QM6HPhn+Wlea5ZZ+R0L3SN
FUucZTl2ZBrjiyEeWLT9R9FayP7jOV1/y06bB5JLyPvT/sNyehMWdHSL46ZSk/j2/RPrVgVKNYoq
Bbnm0KbJ2UEN3cVES/hdDqVezQVcKqvgMzNEgGOE5oXnB1l6+V49RvEwDXobyiE0AufLShky7SPX
CMG0Ao9yEpHs4vY1AunrZR4l532DqmIFg2Zam9UXYCh0PIqAKicZfLBs3tWaJCOvG9iRf/miZTh4
wj1i+hSvnn7dtoZQNS/gACKIlUUKMx9fzWaphlYAXoK/XLk0wfq6Cy/ERWBQKcjbc8c7U2DbEdhY
OIkkngwY+h8mQkWUw6LVuaCDfDVpSKAmKLrIvEWiJjLz5NDgfXP5CBygtAiSoi2LC8RWQKxOeY5D
t5DtBLb9L80w/LUl7MvDZvSaCU/ktAu8OCrJxo5npuX2lBx3NkcRuSGmdfii8S+/IjXf3QuS0IWa
L+ukV1Viz0OKQ7k36438G6xTtAQ77/cdQEvWuSF8iyFEOB+ao21Ev/jdPF/5wyjETqMmo8CP0oIq
rt6Vg4kVZt35tSFqGbHPHcUgAoMu/0pyM7PSz0n5BmrfIWU3J7bgMTjxdNVCGKHb9A0dn5vMIjWc
u5aAkUSlmCKogyi40yax5fqQO3kluHDS4aJPbv5YsH5fqeKLHAOFUQZPPTCVnakrEMmH5LaFb9z5
t+Vd/Nkt2iJHUucE2wPIfIwb20JVf5EqYSUx35AapnuRq0SR07laGY+qdDH7ZZwSbqSNx9JcmolB
T7Nz0jKtyh1c85BwMfkiiAciAShEON/N7Utt8mSyyo1pofatj7UsvP8+cSbveDVgWnqkK9zuKIs8
zpCHTneuKFp4wZlMhyXpzN3bGDe8sGPWIcYXs5fd1HIjMrZLHqDiO+R2Lqtvbb97EpEg44Lepgyy
24aX76Gtz83OyYKoY6RQraL71bv0teTueZ8DH0+T0bz9VZKk0WaJ0o7x5O4UYSKl3+bQujBJHEm7
b0Yilk/usgRvHhAd42PHL8JHs5Lmj8evEGGC6EThFhdxfkrLPXuat67U33lfQRPiRepArbItQKCB
geNMPHm49gx4J5F7S4QnJTEnnonjLmh4vb9d57hWBI4ulkgzuhVnirLAo/kqqn6RIqDLiG4EdBq0
Xn7RtBnV5ckOf3t3jgHTwj8GgWquV3IynnYH1wsluSXDcbd4daf3mT0cH20hga51VumiwkVCTVF5
QjPdAS4ehSMnuR/CYbs1ML35ZI+MVUsRnVh1zMsV5O2hIaVY9YKfdd80Kn6W9buZSBcmXIQGU/YR
IZIwPQo7i5u07OquO5tREHTEFL7ivT9UqJVRa8c1Yj2z65A6kjTyi0ENYe/cLOQxsgpXexi0FonP
OERA7SRqToBOzpBax86kF1vBoIM0cAYucZeYLwlvMQX935gew6Y7PatdBEet2MOUNHQlZ0EAfIoQ
CZpFet5KzKhS2+Zx/CC/sdq/rOFVRoE5uWK+8VMNENahuaMZxkqHabthHT2lkIvgbi1vwkd13qO+
ZD3UO+lphECoD7NfinPe7NjlT8nJfsjt6nSgsvHL26MrQddRplEzvdE5oVJJcuVnfwvQIX6RyX+o
3ZbVmBrMMwrtJiIzAtVWFuXsa3agTiv1c8W+b3hLukSeWNe8YBpOb5T1mbM+ASS594zYjnNSlKb6
9B0W6ZkdoN48qDtLvi+V7a+uSQcJwpuJt36L65jQUiO4yQs0vkQoY2sQk0ZHJXf1HncgUd7msAxI
afBic5ExZ34Nkek6hr5Q+BEJ18GOgdJePepM24NLC/a/nmXdTauHAr8wzJ1oraDJOHpKufnJtzTd
wdM6DupXAlnazDv+SMEezHWr+g2117eLRoRYK29sCf/5wWhKUA4iDHWy9FcJIEdrEtgwwwUu1efH
Bi9WIGC1ALC88rk1fbY3CJYU1dOic4LACPjwHUs6xvRISE8aTguGcFpmNzoCbNCY0tfAE9IwLx5K
R5lP1DUIqAjC3t9b4rr6KXOcAYSXRTE/x5LD4pgeDHsY4Yv6kheQ6MYnZNBNHt03UwMly8/SLV4v
RIZd63gmhbajAu3agI8u94s/V74nia8A8gSbYvb87YgmtPTsDhmcjVr6Cg34Mk4/jptCMMuqMR4B
PlmuvSvNKMIXq6Zngn2x1H8DPleQ0rVrd94nAM2r93rMNkQzlok9uB113npz5MxlZiXLVHYAo/xZ
leL6B8wzCzv1wbtZgOvBkC7R1QfQKa+J79T3P4vS678SShHA7lOO6XtspHCFUiR/7mU2UWvbq7pN
ZLfUYWyvy4ysMW8RfaeHuscT/Ee8D6ze2tY5mArhNLQwV0KH1hLIqVVpYFCk+ecsiUYOxAVXxb8f
c1Xz8p36zcAOtF6zb1IBFYixmiv0v+rRd0tdzf9Z90F0PGw2KFn5G20V22k8WSNjWWkZ4MKJOC2C
vqCkgoKezAc5Ji3YoEnJkW0/Xg7vXWMXzrpynXWpUuNOiFB02xov3ywW1+o8m4IB7Yfo7AZCn4hM
BW1paDGMkcHGCFhvIHB+sEN6xnsAwB99ZMHBGaycS94s1+f5v6I61F+lDS33y9np7bpAwDzG0lTT
S0Vo447XKnoj3tSrn+rg+Nk3Inz9Cz1EKYC+BqXkBXrSir2+hk0YFygYD6JTHCloEKm00t5Lkk1m
J2a5KKBxWY2VQiB/VnyRSqndYNmuTw+QvqPTE7HJ7gLjHOGOQSicF3kRQkZPjXZp4h3z3QGuY/PB
9JdLDoocNA5VDuQMO0fEsRaU05F6d5CwCKx86AofDuW5PthuDtrrOEacwz7p6+Y9Ldp3uIR2yd0Y
xWxquXYga8jgPMSXuEKLWRsb5lLbnw4V0U9twNeTY9mnkCqSn+MP7wgfhVneFXwo7lQGkSWNJED1
xPvvrLGBOpHj0w/YLTgEMMQSxvWuFDyN9afhtGYrQjp3b1NVuNl8pmod76331UN41Iw2yrFXmn4i
R3FRSH4IoKqNewkrBgiVujtvz4MHqJB4awv/jfL36Oi363PxlxOgLA75kityGC7Co4ytqnYmnkTy
N0Cww9KRaV496tEB4/Co76XmuksHEYXgtqhZhTmHICMnEXc8kbdWii2JSTz4RIBMAuOtEMaDNLkb
ENmN9GB03qrU6fN5rDL8Pty4BgQufEP+PbmyxdRar4JF5yoZHjBLGtTswKJPg95UFxf1zfiJohdt
OrmwkteHTjRrawGB/K5l7WEiQjAaaI4o4QqYSZXfhVCsHI0PKZFwUC74DVY8YxuXjsKW9G2KRQwn
C77bFaziJL9hbU2vbQNcdBin7oAGCBaAERkNiLZ8aZIR6BRQiy5UIiL5qGAgIXeeazav4aRfQIFQ
z7/5PDwSIs2/XdVuc2qXCC6XTFiGIacRaxSzmoEJruPAab26/4rrO9BVBZwobia12P8ELOXmmWBY
EMkfNHkrB431ZPX1cp5dlMQ7PRiXwHbujXIhnkfO7g7MNHXjB4VT6+YEA00fgkzpw0VvPjANvP1y
fLforZ4tpimrUpZAJp25QMmHK+hzN+3du0GyXPAB0HU91uQ4ciAbX3P7w6o5et1W2bajZmU852t9
PsNMbVKQuaZL90N21RTPFRpPxCrnyvmrC8WlSYduEdGTeuFW80EGMwuu/yDgkoR79frrtigKPk35
3+1arWUKWbeRCpixwdMX1zkgxf+/2e+SP1YMwawKzmi//39WgU/s86Bu5U5JtUK6u59fTosRXpfb
qH+KBwFH0wmghprrrSPVq/wcDitwN0WQoM3q3cDi3V8/Nu38e9MvEgBbyP6/GS86gwiK8aqJOXqw
SjFOm745IfaBpjbM1O0VsBAq2uGsFvJovZgxf1mKDI6kGzs1XYJSOXy/2HjoetX9Vf+5H++8BLdv
HxAT9bB/pchVTvTBlsHAcVacSB0Jml5RiE2dBuinmxkgtqf+KG1RvS6XoMBDWotuqDhN7BPTvQxo
ZNeVxGoZXRM0+Llo9jm63bQQsQs8wuh61dvvIYbRbWmQRKovCEiPw4TblUk/XQrZsDXVREXn9MF7
tBHSFbZLK/GTMayTpxrMYv0cAMybZFWQkZq5OZkzS/cT2VVPZSdHv1baSGFcKDHJMcn1HRJRsIbT
OlKaAc2pnWzHr0LWK5tWND54+ynkREMx2JZO593Hg0WsU+djwM5KGNiWel/snnRad+ZvElv00UUW
e9LsKQkeIxQH5RHZogzPbshb+J5NvVDO0mSLxcV0swdM5r5clBUaL3QIn8UKYPfAWqPfAiO38e3B
bHFAW9XfDLzIlZJqHvlFIBdVbpXcW4F56YdviYxSeDfMM/Sy0DCcMVXg71AsWXMdoO4E9vjSW07v
j5NBXXzEeD5vCxY2xpgj2cBTOZT0e7L44Hy4xGzyTOsTH3QKH6F7sswE4dqG4vG3gGW5MnJC6MDT
APuSqDRrfrkn5nRC0X2Av2QLV8k21mdNaTbcXQv3RZuhbAyAaGi8Gs2iTAPK00cd6Z0drkoU2ICJ
xoQtnzsgivBBORewICNayZsISMzAdcp9/watKKcV21TJadFudyYmtscI9if+EAMdNnjr+II6YN/u
jLwhP1dhxi4scISTYh8k4xUgywkOftxtmWlb7wq1uoEGfM0pOBrAJbgtx0GQRgUltTdGSo3xPnlY
2xcUjRThL5UMUxQhfSePCMdpiKlAzhqtKkmebTuBTzkOFT/xy18P4xV6gXRHrJms8JxY/VMqpn6d
thPLnhYHmLHfEyIiR2J48w1mrUNaQ8+BLy4UgS4HSQBY2q6ojQzxoykDy6SJRUeizx+3uJf8XWql
jYfBvNhrON0ns010fhtQklvHZb+Zd/gUiqjDrYfHNlSXMTgk0Vq9V/ddT4c2+BiOdbav/ER7YSaX
RDppsci4qaA0pmRc6w+Y0ASyNIBXGzneGMK05yeAKagM7dAxKBHqwTKNrK8oKxmn92yhN7QwtdKu
KQ+arA55OG8r1zCzZ3F56wZep6M/PCVL1piE+JENbSEVa9HSgivo7X1fGUvqUGHJzE2VRUL2G6oQ
Uu+t+pq649V/cCw82baD1OS7pwouG8jxfvWSOLMaT6W1rThRQXQ1jN6+Yc0rIfm5mJ12WOiWF/8N
WaW/ei9i2dCDHVnk3TpH1yxJIcz7InIEY+QMMbKb5r09RXrwFjUyG2lENGaV8k8lNvM0NJBTmNtS
Ld5RR++7r7vmPNZ/m2UkOkWZ09RMDTPwghooSySYGJB5r1b8kR2v7hqC7i/Baqlz5jDBnlqY6gez
oV+/gntebtpivs55+2GF30xcqpSbjISQb7+vFZqT4y1OOLxKvEUgit7gKC9LvCM+d6oI28eYRx4I
R8V1T15Cx734ZCgYTXG3TqZOkeGIo055NuPZCPgMiMzf7qtMfEFWzxfnRIxBaJaUQbOmaUw/JnXj
L4Nl6Wi+E0p1P3CGnUktqRJvnYSnMePhBazrTZe7sCwsDxKh9Pv/T/NcRDyMPdTo91BjrNgoo3bi
W9JfpZ1VTpSRVsRJybte7KLS+dxE5lsGjLhRsVXELzI7loT/lDlCZciMXrvlWd0CewO4plfKxBpy
+9m2PMOSEAulOhwg/sBdc9lyFrxqAUqsNW6WVa9ygk6ILb4kYfcOMbCSmKnPoai4fp+HOC6vdusd
lOpr6SVIEohOf5OjSXi/MATRb2fgiIbHXUPZpCGbJl5tZ/Va5CmvJ+Ky1w6ahhACqosa2IJ4sto4
G85/wq/VwN4yXc0t+RlyGYkNiiZJ9moBK+tdeQgnEQ0hQujLopp2uJ7VCgx4TaZKqCdjjbG738IP
wentWQJL/VI+EBxTnwnKE7Dz2qa6MnKS8lS4hfPQPzImyoYWibx0QbY0XACmAqGHUZUe1z0hhB5h
z0FBqqDjZ5WPlJIOpNFwJ5xUvOGlliBpiKFatJs8Yxc+HiUd/NMLtMX7wZlGK7vzAhj9bDx74baC
r4hvToMa3EVFmZ+I5VwtiDLvFGuZJ8+k/qukw/ReIx1aFLZJxSJkTcfoZurGm7xpVsYu3C2AMjAU
p8E1+nXRoBLv+Napf16e7155KEC9rext9LaU9Rtf0vy1ysTYQrdGKJx/7zDSwPav0MJ6NgwMTjkg
3kEhIWawiwgpzkJ6JY5SQgTPY2qOpq6YOtblK81oIb5LQEEQg9K5zFCR54f7bjXcxlyGiU6ZCymv
iLTnne7ebeRmS0DgyCGaqHnimWVnkoQKLjN8gXPy6DVr0htpfZJRhQDQ2fpc1bi3dyS6P5HezTY5
hidUGoHFxsaXGFiLYxvFkd/TWfVtie7C5KNYL0Xvn2G4n2K1ddphWZ9y3RUK6KYyZ6EDn38/dnQn
dEQncWob2NR6xdfFvc1bf5eNsHXn1WmwoP2KJbSnAU/OGSBdTX1MXME1NrhCj5YllNiiIy58sqhP
QUhQ1DFIm/VBr+uEvQbLFu2yxyQETOovongzdli0MTT21f1GsimVKsQYpJCvFBqjfqJpLQVpANwJ
mLOIm8x0VemSnBBwD/KvbzIkF0KAAxZ1xOrNhb5MDmnCRvKdblemrQOz/YlVXiWwY+tCtTc4/8jN
OZD+9/mCqaElpYWrkWB/X+Ay5HpKYeMEgRwSws9/+vP3ZJbnmeAf+1oNb+yMdFRKBNNGhwj8sc5c
WMmtLkuCllnFYHFXguSNwdD56FbgUCf35jh8+kBePCqvMUotEZnHt9bUvKN4PJ0+uVQncVa11KKg
ANO4J/dfifTG9t8f8jielRrdZeCqgt7y6NQAcImiWROUbrIZywg3UGhGPV8kgymOV4e/X085YpLz
AIR9vQmYx56+S2w5sh531CjhTxFXxMngO1yuU9/HRmdY/iamEwEhNAGgJgKtsKmdutHJXyCd9OAR
TBjHDY9BJG7POw4IJHzuhOLfwligQ8dS8/KtWYObcuHwtZ7lsFwTtvbW77spAj8uU2mNffu0OGhR
MKxBrm3sTNRnh3wJWl+c+PZI4u+COgwYpFgKdeF2uMGeFOWko0llG3GKhcKDpyo7HWaGzHxfXlmM
vivV7Re/REXulixnai00v5rwgYedfUyT8mr9t9VGb+Gw0SRnlbax6wWLwmcXrc/R9s/ifaWMobkR
EVbAxTZpqA81FT+XlagsLWRluoSWy1dFEa1JElm5qEjHFfe0TT9PgwiP/G7LusRQ7YBd4wgs5bJ4
kvylbRML2TxETPvcfXlDp8KzPBws9j6nIi1ntWIvt/2wc9hOvGMKLa0JIW7taz0JlHBClTPs6WJN
BjN/xvK+5Hap3ApaalLBEwMWEPNavMVhqgbZvyYPUA4qpjjn3Eb0eeDOefEoKrh1IHrjD1aK0JOv
tSdA5wPkgIKm43jYfOSEwAaZ3qCbsVozyPWKMKhogLCbyg2/Lv1bMGfgItQo5qu8wgLJXiW6RQes
SmR2FU2fVXYdpLkzCcqVfC4DTQijtdCwS1VEk4ZuaMczeP13inYv5hc2Rn9vuYqac6z1w9vC5Jye
l0DlJv67rkGtT3M2nCQNPdeRWcgXTaDxVwLILANUwkx2AlgzYeP1oD8kWaRExCHwaiW0lz2qDWAR
C9T8Z4KgdCUZ0ygLZBv9aZ6JKCVuDx1ZhlLHK0r1FlEkOF634LGifn+hOl5PfNaebkN/9+pudDWg
G9cBltOLmSYWaEgRcGMwTDtTZhcQPezP22/HXOJWVZsQ9SyIU4YPKRaegQN/NoQWyQG4FQteI1Xt
SFtx6j/SrYr4TS1Lr4tYGtBvDkpo7S9X61EPXayB5iRoNhIta6sfx4fF+ZuZ7GUz/ucaDDBnSCFk
kjlbung+pEpA+rCZaTzMnjcEeojhEIvbCBA1V6k+8DO7m0lvTre7x40voCrN1rHPsOamVskDAAzQ
yN8EwJPHaOucJC5BDxZLgBKvqz9LmZhOrEAcfAa3B9qKQlMj7ZPM7o93SErXRPpyBQwXdGwsT5mv
FYmfMbyxCPAFdWbQuBpP9GLa6TV/BeXUDJWKGIglqgGi9NJGsSlP6KFwqz8HcOqu5xHAWQvCwNGV
KBPdqQOMrMh+hRaDgyM6jwhtmL2SgoeTFsM24DV/7qMKOdMcN5T7pTJsYgAtiU4wJVPVuwJh5tmm
F4q+sr0Xct1uXvsvndKkyg1XcaFEhAfNuNhyKZ/TZ3fCdGQXLva8Aci9gHyw/wjF0Az03MX6c10l
uypU7ce4FRrmc7cV/mKEe+RiWqgd08Q5FQNu3wg8HkaGEVS8sm+BKl+Ro2U1URne7hxf+qdhBzad
bZv8Ynr5wgJN2n6jTqBf+dLKe8wg/efvgXeOParlyYHLIG4tdk9EoA5y2TmZ128PZQo2OXXzLO8k
pG4O67ynr3EVwDRtlqdrCpdN5JnC8boPIfhN6ax6shDIi0oddexb1YUA4AH29+R7hVeahF7LnbzY
DtQOA3dnTo+SEuhuiIL0NraVjpSvRHMStWGPILF68JAA+Xwaa/nPmuabxFwj4Pyj83TqD9l6Kvtl
uhZ/gGroKb0sfwEt+GuGgwBOivbYXuH1Tkb3JV/Q+fA8wFjXcU4TUCeS8MqisYoSVb+7jmoZv02u
UFEHUGmC7DHfW59C8NdTvIJZw4Ci69oBJDibiyYPHJYk2Rc9k7LQsBydgKKIQOhHNn13M+bS8GLX
vWratjV4lReXT2ssoZ8DW9ojcu7qrt+W8aS5+gleC/Tjvh0SEzxqA9wodV5q4930QM4LxiZ1BbSL
ny6UBBz1CRI6vlQm3jIfP7GmlHSpTSIDPmpp1DMW+QBOfhdoQ/gLC+b386JWQCwXSX+FLxGolkPe
Fm25VkGtRRNqCT6qBUNLESKQfB2s3CYtuzqhzN5ABlzd2MWNiFNVlZY7y6jaeYyzkD337rd7DUkZ
J2qGbF0gGs4b7DTCxdw+IMJzyxHwb+1LrNt666Xxwmqo9WPbHmw9sD6jZ+oHE4wLafVakSM0sIzu
bir5NCux1XvJ+r2kteOR2TH+0YLaU08IP3az/0q9SozF6nfDv/po6QZuD7r2RYrDjgt4ES1pR79D
j4oxC9zgYLNw0Gn47XhBWmQYXIJGTsdEXnNIUZktriU/7hqPCI6uO7tth7NrDO0Tnzxv66QIr5Ih
K26GdLWoF+Y6uPkPJZJ0W+Ih8wflKTbH3d96AWsO/jc4GWH8kf7WDcU6Fj5ebEJCHJjirUTxMv+Q
Lv7FdhqzjF/DYwi7oesK98OFxcGa1+/w4k7NurhMORElFDB71jAfSU7gvNEm9gfxgUkvIL4UKIv7
t4dBVJWYGhGiABIOwthQolnBDHNloN4dP1aaBnjY9vFnzQ1imn6GaTQG8OziB7++bFOrk/+u9OHS
88i9sALwytl8fzkZLCsikKeItBflsiMUULtKDsQ6zIrCNqhSqtWW1ewvrEFOkv3K74BCZXR6u3uP
LqCSaL4Chl6k/EksUc+ewYZa5tGBPK4VOSF8CQDbmAurn7wBaLf3Z+vDqOlDyO20Gf37TbmlJASc
+TjKHYocRVFd9SK2V2VbSSYfI4EnViIFlYJQwoBEmiESsdBTQLGvTNvhs+SkzgPUyJ/ISIzwH2IT
Q1zEuLo9Fthbh3WZf0jQf6sN5zf1JfLj2YGknWTSnKNNdm95egT/tXeH9fx3UPFBsnIzpCeyVxgW
kTj9iRtizGC6x71qrcZNHKR0HA3yqbKZCvpVpo4js8zkBmyZsVzInuzpvnP0NZ4kegAXwCaf06G3
uPPQcTyeNFEoUB22Ir0WYyWUnf2R2/LGb1RFk/Z3chsRbmYc6+gHfgiAESP4zWibuG+etYjpHbAJ
oYZqlDMTwwp3qLF8sXcza7S7+BZm8ZZ7ubW7WAL4wFeAf3lpR2d0oQX7HFgzvYcSXqTqZrYbY9Y9
RBmYfy1pyQSO1IM8UMsRpwRnUGw2jRFWW46ZaHJZzKo9C8yRJc4wPpSirOxIu8k9/s+Dw0opy1gG
/jGkxPB+JtTznJmcHXjMEHw5mjaSSkD4YVeccPLqZF2RSL5BMUPXW5gnKXlaFfvPEu9znKSdSWMj
6X8NSYsaLIJQ0JGdUEVnb2nItuz8yAg/+gAW+1vGvXKBEgpQzJTiGlz02LeljUhKAw3pv08uxI7B
vkuEX2rotoVsBOtVQi8dvPgcwj57oawv1Reg0Y5DISr9pEtRT14Vw2KcrwWEXJ/a9uSx63S2bQQC
FPbMSdyGbQcJASvxK4WSgr1IHwWjR4SeZQ2L3cbC/IrLZONKbEXTwFwjNGEMCcXOaYbUPsirkoMY
++BXkEQPsKX9gSz8tN30Fofp/Y0JbUUH+jrOcOe/MZBUjuMVzgkVPybjMUP9v9b3AnTKQfG61G+g
94CC2CEbxAg8Ff9qQERV8Kg2wWtXgTS5uRs6aIrODsxDH401YUfQwLbc59BuN+bNd8xnJVa1sOUN
X/dy5qTt47/zx8qA2PYglO9dOpW8tMPRpOvNPjWpkJ4WTzjM3iPK8ehnCZyOwbwMTZtkYNfHvr9K
OK6YVc0cdgmvxG3Ra7FFh89GytLDqdy8XWOWQN1LU1T/h/1/hyBLHhYYj6QY55DIz0UuunJkujOO
zKL5CMUfo61QGMcjIxq6v8aJYikDIPwB06VsMEjRtT77obr4VpMs6cFKZGNdhKDM4lDxqsDbuATT
HZu5VdebU0h3akZOzDdF/OipqPTV5PEXxzmAk83uVbgfholX4Nz6P/vBIPoWiM5pkgE05VOKx8yy
QfCjWu62PLIxTQHPiFh38h6TQ6ZnDxNIOz/1Sn+B+iDZQ7AirMQf86gHCrlOIz50gVCgak6iupn9
uk4hnaxlJ6zCjsjp3SOTviCEHMiUzSb+5bJwkYAYE+PcEzopudu1Ck0aUFjHLlZLhU6uFC9GMsCf
h8PvnivXtRmXD/w3unz2e/UqSJVOOi6+PWT9+CQT8zvWVyTzT6/DLaCs10U1Dvuvnh/aRow51rBK
57Dk7OQpDWRlgDQz/Uxm+TFl7zqk8iRULZkLo8hJ+r5uB57hEOZc258KtN+PVr43xHZx4F8ESoV1
1JMd3zAdM7xb5dBla/Ex/zm9MrmZHN1Hcdt+dI13HNi5aCxsDOJx5Q/7VZdMO5aG5wScNz2s5M8g
nxXOxe/TvIM3eo9FSsaSsZvR5EOpoBwWi8zCN2b6ETAaEUkmGiprPx5rpA4+hAlIiVNyuV+TtSkk
I6pzSKOSv6cVsv0qCvKU54GcYQI5bC6xSyhHTllZe5Ic+WOyPU5IHShUSbyjuaPDXloH8PteKnCV
A+J9p2zIzk6WBlctIFWCK4W9pL2xI6rrqeWdOInxuSeS4fLBfO+/+DkyADa9BlFNttKL/wOeGnL0
HwdzUXPzbbzu5PbuFbOd9RiK0eS+JKHslr9u1FSC377ZM0DT9ENkwPML7ua/3dECz0119KKkVPKg
PBD/aGRMopawDR0kjTTs1svxzViBxfbwcohhetEJhObuCB6P6ZZScHyJWZeQaUSDvPz3k/aJfJ8T
yvgUd6lcYqQOn/QSMLGmzoVTVKLHyTi2I/os5xv45fRdNrh49FnBNAfkIGcKrpc5Jo+o+7IR177A
TdwCV4xjGNZt3VzNMyk0eg53gpZAaoX5XD/LGT/Di2I6g9DQeAPDBcZwCVzsHKsrjxXrcbQZwwmF
x/V2BUT8ytifFD9QmOtrX26zDRlT750NtGzTO08Udg58MNUg9c3BdZUeDdkgffZdMQETukyigrN4
CeTOAchHjvKYg0tS7XtVjEOn2VqnCWtp2PKoCRYwqUK7PhRxsjXT/q55jJHW/at5Cv/V1wKeathV
D/Guq980emEaZ2Yb8cG9m+CLKAetyvrl216QcxtLBEhyQFj/xAT0+efxnKCIhlKE/o0oE842oGwt
FOPHBpvv2es3EqnAZRbiy5CWbftOgEAGoiM4GyiUKcvGPk5LfyHrTdKcqFO1UkhYnNZd9PeL1sHh
Rcl3uZ/1sutdYCyZ34wTUs301ViGDFrAtE3R3HXum2aUmxFk20KCgta4Xkh38R8Z+QahheTp3Ouh
B3/eTWSs4rqXsN6GC4j3t9GW1bYa/duh2XvFEXuXbubNTtNzGRq6wNQfBzZYVSB7LGIcgzMSmPsm
y5aILFDTWTZPpS278rNjFct24eCiTrccmyvg1j9+f3TmNnPIdBeXYeiNqwrqHy9yLS69VtX4sHse
CcyKYLGqXjEyTfWhOurSmKjyCT5NWL1U1M2wOB1sSi7wmkZgw4q9WPiy8B8bFrUECvh5Av3D2mx0
SLzIHHH0TsLNHJfUQAJ2JuAFZoHnvpYnHnuXgf3G+kSoDPPbQdQDqLfhWuMXQTmjtWFBX7sbjgMB
pVy2z2fuzViP79xD+mVW6Ndh9XdmA3DrL7BHfrZAnnDQSq9LTDbmVIwdUwGspb9R5zdP6UJneGCN
+BE11D8nCmk+2G9EpVZ9g57JrGbQPgYun+pt5VfYxbUfpmgM9Yt0bvu067PW0AL/5L5ca2RHPTr1
c/Wz4ThV98yiDzYJL3GBtFH6zvkJanB5i2zI5+fGSa0p21imKMkJOpxRlYM6O89zc1UTURnFioRv
2tQ4w/rFEuK3RsEdsY6hXgygLJsQjG/l1enfgmRIpOCcZ4B5k5SYsyhfcf56Qbl2gIfz34vnOogz
qRqoWEu1izSdK8xKBIhjd+SClOlaxgar+xHv+TL/svvG8iakqPik5ILGFoeKvKbu30EoKkBUA/q3
kgopiTW34gQBYlCnzeGlvuqzgOSQGa7MPb8aPdgMIEAMP/i7OFn54WBZdH3RQI2ZgH0gzpTFLaXL
LJOrazIqkKhgOWGLPRBY4zVScJlmft1ksAOjLii4U3LZbPLaQLysoPatYV1zviho7LibfpkWcUNs
m8eG9LTffYScB1GEhlJUEKcH25h9j/nvj96ewi/dgRURHsz38cJR6IpiNe7RcQka5ZxxYkQAM++t
0EstIszicwztbuHKpZgWGB06c7A70Fx3KvUsu6V2g2KSswKEdIqY8VrQQwtFrtXh44abV5huaUHN
vatpfTz5dvP++XAmQ+z06jICRd4CpHjLH8/5IoRqtPWRrOWSr/qbT2LR2glE96qoSF1Cj2UuMDGf
S1oL6OFAibo50AQZ8xzS3yxHb9x/W82F5NoR3czRX49jnCwuRgA3HxfPl8vA0FFo/DO5COAUSCT7
l6cd10AE7gu4CWFYb1b0KPRgpSGgGuYADXbrojOBkw1i9Ogpz2i+yu9Swqf0jc9iJrt/01xRXNC3
H0ns1/VK7wdILpvivaZY318r3mcHRbp7uozHL9CAADaSzff/hdOOkWG3Qoc7kTFSq4phQ0o/nyev
BkUK1KZg+cJsitUk8/XyGtLhhyKyf0AEuvquoq4JHq0llDZbTbD1S0odMOT8svyqroVmEY+Q073l
xIgYM9h4j1ydvnpyKDqJ25X8koOsUCwANxvci0d8E+lCANxMYcj8pSpzUehw1q7566jBvl8zM4YH
IVkxYv8Prnrc6LUGHBbPBXHK54posYQNlTp42CZ6rb0zEA3wM3qeAzvTVPAVd+2GgAZFdE3v+cTa
kmcc3dUX/JLOMs52h4y+V/4yTRqeHBkLUq0AW9fT4axSdEJHPqJH/QLkko/vKUMdM+rRWiNCrODQ
h3HveJRJmNtB7+BCG9xfG64EhGJUquP2ok7WhTYu8KxLR1JNonOX73KFjxMzTIdZbvcjKRHWt8VX
bWzoqqY+jUVuq92OQ1udNe/b7mk6jbp2bZGQmLTuMcREZj093JqkoMr3Kwo8w3ofmhHrxxztuZyN
Lazeg1bh9EXd3HXqouk+vwbmKR1bnSTLjV4DBUNapDvXkTYKwbxqIekwsLQcV2WKKA0PP3RM3P1t
dZFrKh9Yaw6lGBjIXhqQbbdAZInXBvED2VmT6RM7PhuZEISECd3jAvJYKWK4mqA1Bm5EHlk9tKyO
gbnuuPp7pdEqE9njdpkl18WZ9qgOUsfq9Zm6i/A373GLpeFjg6SCXDhftipRGeB95FphL87bqJM7
NPmqCGM5blSFG0ZqSE8k6DlNiquCoOo2MaazbPcqGUTbEYb07RYR6UZNhfaJqPTVw9fypWbvaXnZ
aGoWcbyC3SJO8iKopoUo6YaO507A5GTrpq99OTqHkAwhUSFMl8LcVmj8PquLudmuzoiZR924iAzd
SXoKS6QBCfcRvZPef65hcJhqNNQXuYmjI6jJDcXT55i24DvUno3OaJf4lqaFMmf3QM03vKSMVZB2
Th+LovpYdPNHgMoFMfbNVO3VDfKicj3QkN0p0+BDe09OB6Gwpr79mJt5dswyAY6ht8DL0kmoZDRY
f+orOLJq5ezeUqCJ8gpqGK1Ie6p9xhFgZwPEE2utTmfRY8yBXmThyyazGrPgMkQXSBEiMBqD//tu
2RuMuL9iyeu/vaBkfruCRs1Irl1x5wlhE7ib4gSjOMXRVQf0ERovDwq/Md1bYVujZVgG7oXVjUa9
CNHFvVzup6/YNHZIyowoGcDT0Wd3GKB6KDDvrcI2d3qQ2reI/mt7PsUdGBvrkksKa9bAqeZuvL+u
rlpheW9C3LXEOGyfJvnx3PQzkRfrAte97J6YjVSUJlbdKhN1ZIGErcfapvlkXo6JwaDg6FNit3fm
qNmSmI5eJHK9NAcvXveJAvWzqwHIjsi4DMMo1LPJnPxAVUlOpTvA0egW3QiqLY7e7iGPKaStVb6K
h+k917bm9MN7rSubuX5IY9uQP/JH+DvWjxubSOuYOpaod2hW8Fm94D5hJ8kqTkNQw6RBUW4+lOFC
jPBrtU8x64qdDcAbmUGO0EYKmCUSmOW3oOeDSmKXMlcTVLbCBJ6gHaWXRZW/H+6MJQcWi4a2S7p/
UiOjz5VLUY0suPP/v3lgbor9MtbYYKGqIq7cO8/qWz9ODMeYJbs0JLhJOBh14UQ2N0Pz6uO92Kb7
rR+36XlgpOD64JPeNLCtbhk06DSApcJjmdypjt5j6LhAoPpjjNJux8odAIREWLLvxCxF+AD5MCIA
60Rych+pebcNkGAVxumOMKxjHDzXzUYHKuNtd5QZLiqmLwvUSrZiK2hqQ3QYbX5C2/JNK/v+ePXv
pozbahLtis6/uLyJalguAmr5Bea8Q+wmiNhmFq6s+R1/n7Y9bt7Wgz5WVGqeH177pIDKLVDY2TEw
0nc7NSImY1OUddczihm02AJ/nnUpBHhyZ+JvGNdfhGQRUxfDcsii+UMqnH/ZeZqkWj/swNFOFlYA
P9TLrJFt9yEQZWr3TSzV6Vs6GIVAA53fFFWcRd1P2GdrcrK9viwFMz9s3ty+ewhvn1wkuH3m4v2J
CD/SRG/D6f0VzAtbC8lnTNBQ4dpdjok6cyXOoBripVczTKR57nbXy3PhSWligpJiJ8kLSpKK2Jig
p2V5+Cg+CVZ77+MU9TYo925wE6G1Ebf5kk5IEbtnnvozNcRrYNPCaXCtzupSkNw03fQQ2pBrQbSj
Lu+Rhim0NXXKUubrAjD37M2pL6e9XJ6NM9Ff1pRGrA78NgEq4QyyUPdUEQ62EYei7byZ4Te3Od32
qTKiyOaphtkYG3peGfwnkVzYQJj4JP8rXBIw0kOD1mEDDfrnsLBBCLjta9Ia6EJrVwNvXd2CaGe3
hTAXej6ffavwO3z965O37kYVy3QfrQk/mKI+OPjEZB+VdE+uYCAeC4W9NlUV/xzMocYtt4aTt4OL
JCJlOD9UgxtZl4ZuG/KmCn1ZISI9wIU9nbDIdNvcnTdo+f/OHERJ7JJOz7sBwRRrgrUdRzxx70Ej
8ccds3q3gpifM6kVuYlJoc0GsGsQilrlDygRlJOq/GehmqgVlW00zmoh3HGcTeWibUvVGN2cUKWH
ZdnKPp1rl1OUH3tRandegWAKTX+voJXgdZWcCeaxwygXMwrSKG/W2zCX0vkMu16jbqlGf/GgRxM0
fzoofisz5rfyj4CdDytZqjH3MHgf7XU4qF65JgixR5Kcz9FEvXjeY7V7zvbpkiZPIDSz92U8aMUI
zxrLia2E0l6aY5zNRk9dBuZRMNjfzqAuTxmFCDLzsfJ4k1QqtkkDnxGA4UnWI6Q4M/B3ZM8bqqEr
p/48g139db0RK4ZnlR6z5DQASdIFDxRXHVw89K1aDjJpIVzY9zTt6OQvF0li84KJ23Rsp4ijaa9a
jPevBYnRGBTLHSZ8rZXvP8XUz99/rv/W+TOjol5HbLMVQX6xyYDYCG7PV/I9X5P3jwEUkAMjzcwe
unvyRD5mhV2UCj7s2qy9b/mkLWgrPQVFxDRVnfBLALXbWRvcTJwDXH6q3iC3hUx8Sj4/C3io5DmF
6B/STxaSP89ivY95GiQ25byD6Ap3Cyw43FQxMOCIeuMo5yLz+iElsH5LkeDj96HQ2ni8SGLO+GtB
lanPpQtwxYtuNxsCX+NOokPghTtoFcBz7D5fOSCXDLNAohd6szcGYHP8anNyIR+aaiC6+9yhuw0A
h7qCFgTVcdP8hZ08ETKlIfJPA3EBdRND4Os8ZhzO2B1mwOnUArNgiW2xBfcja111Vm+iDb/bpY4s
AzTI/z+0+a+KDa1QUTQavqAML38Atjl4sFBZEZ8wtgjynvLPqEKyfOK+0LQcxKcYBfkJiIlIG07d
zDzS2bwmVL/3KVd2ol1xMMnoVo40L47mcNvpiIWNoRY2082wGRU91c9lmq2nZnppOgi9MMju9SW/
3RWXkxqKdONDsTRV4s/F9ymOY8eEmuStPrOnXfDiuRLTHMLPE6rpk4SnliWwt2z/gtzT9fkzYIuu
ubKH8jsa+cykMaS/p39mG/0JO9mGw8hdPfjf6+4xLl/wHp6NK/ienoixvWxPhJU+Zhy9Fq6QiROM
3fr52Bvib2ICRyla8yKAOOuo7HbUlGuvhp+UpVXDjHURr72ugLbAYMmEnvY54k9A9qUquZAYKz47
lOO4uCZ8AGuSXIcGC4kOI5t08t+gGPUXRdsWL0zAWvoFfLSBNpDCabNz6nPIqnIfH3m1deOBeaIA
IBg7jCxq3G8cOA1DJao51w+dGgM50EiFyptQG/RiaO0trfj2mwg1SZZoC1+q+p2QMyRG1sJnrbe6
ayto8L64o3nP9VcJhk+c3odifbH+3jO9W9XqjYmCOggsEzJ7M+qu8rcFpOKCC9IwPHgUN0y8guon
Q12qe03Yi3OmucwAI7xqNOMPPT1Oe6Y8f6OMHe0697PvSSLipTp6HeIfTv+mtKACrtjGSC+sK+Cf
yQX2dCusMketNNjyXhPp/sGQvOj3lAXOk7j5QUkDCO9Q167Q9wEh2hPeXrCj/WWVqrH11oyyjLxN
Icupj0lOE3QcVwMrUjz9edfzY/BMkE4/R6JPrSP/wpleG4XdmLmSrs6OX4ah2NLT1ZTBiSZEQ8Eu
eHk2blzJwch7B4AHSmy09IfVjc4mH3bgeqeX/Tp1GK0vguVNvHLgedj8bCJoFeB2pfPcHCJOv7gp
AZFHsyGTtsYTS4HDkjrOucp6JlHseyox3tcAuuO1AeSA6igSXuQFG96XYpFwwjTD4nZSGbgV+BOX
NJNo+YzGGnC3f4EABA991eqTQkcfKPdkc9jDOs1xrEIT4HFkaQi17c5BrgbzgyUb63scF3NJobOX
sRf8ru5ODZs2/aY+b/KXyC8pBc/yF6Agc/BPUi7Ddy3hy4+lZSkjHn2wjJ1dR3wPRhcEou8EahCU
vYPWG5A7pi4xKVXzJV4V+y1jfSqcZG77/wv6T1koIv3/eTwAJXcdhK00QdqPY6KYToDhhcrEk/oF
Ql0vItAJe411/SRk5yYHOpwF4eM95IJKL6LYZO2yeaTqYYbw/z3SEQo+mtm1Pch5gue5g2PVYKNH
JaTk0U4GaT5vX4syQs8VjpY7Ps1PAs9Id2geXmynIi+JljiMYjI+o2VRDO/EEvW/3lpaOZTsSLuE
HaHmfAdUMC2MXKEQoBVmRp+aEBOdKOktyjHzYyegrrvjMKpX4WuIXeM3sOs5pGKL+z7x0ejhi0uV
HOZZ/kAu3KVVLIl7M5PaQe5kb8nRoFc5L+N6D/j2fxSAC9s6QGCgkIVYa8e7mwIi9jrUGE+s6zzM
GjoAOo1g1d669nnp+/J9q3sxhmZu/z+XmqArd8QKPNMI5bDWVlzInmjtk1vMxwQ/+Dhc3xkBs50e
WGSoNsEjxXcderIUpmoidcy+z6jZU7jq+RyidudIDzesWSxaGoM+wlHErpRSeT6490eFvCp4xC/q
XX5h+NtW3wP7LifGZ3xDFOHnMeSyab0EHQHoUfvcLt62dSGiWmHHUIPBSJbOs5aVur+fLpeSpJU8
vGMh4lAWnlnzjhRR9LDFPX1V8RPBo4FcJHkUe/wS1hsFXwOD+dy6eVxBgipGf4O6lMs9yoPFoiVt
PGUSP1E+X9TofS5CjkH/CjqDBZCljXnP3JnjY1aWS/EoXHEfxL7n3Fq7N+bfel7wDXgpO3hHtlH1
YGH4v4HyxYSz1ZTyhaz7i3E+zX0lQGvb3wRSxftCjP+VIYK8Fobl4D0UqGRRFAXTA8Y276CqtAfC
eUwXD6zK9qHUaBDwHhuDPuLj4/tCxnX9T1De+YsHgxAuraqhm27ltuEDOnlKVUdYNjPN6LPkjC27
rapvRwMHW3PvcFsX2rAVSpTtFERqXJj+o0c89tjsWgpw9LRf2njli4+WvIYczgxfotMEGA5YkRS2
9kBt1UzKCRM0ubwziPAzKpjfrnmBuds/+fUZWkn+Ii9bmt+Mx43L/doeNcPcHwh1ezwegc+HWAP5
2kyoXuMmcTp3RURcjfuZP/JxyRjhXPuq8VZ/aAWGkKcYYCb71F3ATrhMUNginlSIe7aHj6i+te99
0Yh0vlcIZlRcDL0Ylf7dhmbLJViws6EGqin1tgc4+3+hTAlTB62soWpCMz0nDBUnyXimkHTcGiHf
g/9Vmmr2wscZ9jGsaIUwiC0P7mDKgyj9SBrN7pSZv6qmhhxe4SY10SF8Z1jGIlvnWcyhbLS0KoWq
ZZVPJ7RNeAj3ZqMc62eFS+pdo8zXkVQ7jROXfDqA42zGBokVrJxomCKWrBF1eCWLxrHfw3uJioAA
lqUJMYL1zmMewBa0wqkN58yKxefk1e763MHK2LHkEEiB4siZR0oCmikzu8ioez7Bycr2a+16/4wT
BY/26SKgCAIS8rzw5cQzXCGY5X25z6msRJBCB36zhJcPrzysX57LQGLSRzAOQp/gfAuDn+hHJ28s
aKbcZh+iXCkeLN21O5uodpcWhU0jr7M56PMVJ7HGRqo9RNPUYcdfd6LczFFKJzygaYG0RF8xQsx1
IID4DVnyeALp3pcPbeM8gmgnCHmzatd8d0WGErrhBdjYJ89KgAxZXTOqzu5TSNQJ02KKFs+fwph9
HvUkNP1YyeV/YeROfPPkHLIQDAbO0Fxa+Ny9RsvUb64umgziWVM7iyt2mUTTRJJu8qllQw61nStN
bZ+Mf+4Xm3Q12FAi/Nb6QxLKqEE4mHt3kVM5IdgoqwATcu9Gklrd/sYBlXXcEx+P+9NSGJYO9/xS
It6qrDwJnHRpjdbMW2/6TJ8OIo5qm9nw3tuE3ItYnITMylDQeTWF6P/QgToSq97S8jawOGxMl49Q
/cKr3w7BHSw6ZHpz7h+ug3KlVjL3TWkUSLK8GrrJYaAr0TYwciK6iZUnoCQ5BQ1Jn7vTlvmMcQhz
pPddhST4NZ7cnZvlozcbwafwOeEqJXytrAL4rFnaMSMAL3kIQRPJpk8/H568jpmT5SLUfglyAH3F
x2zhbUZ7/5Z9QINZQT8bc9sf90ITT9J2X331+gBfKcMTpALiSuuhSD17pHmw5WhJ1gbzW3U2jgsZ
88pDNep/lN79moTGKVwy5HWNadJiYxi1J55NL8Bc2JCLedXhe455TtgqkFpJsdSDxV4W4joeN1OE
6o/HZghBfZM/GB8R6A1Al8jaxJFYG8aAVAKB0UI8TMnMU601RDzrHNnm/sTIFhMXHW59S09m5MmN
rR3OBxm9+2jXsKzVSJ9Kf30YVaE9sH1QwrsTb+wSa0+QDVKp5lzJn51KPA5HkPgyXWuXMYYU2PjT
MpIJU2hMfM2eR/zZrL2O8nZk2H5bPfyqP/V+3DEFra5gPZZz6ygO4nh36fmYvjNYRRJlRRxEMpdS
lcQ2x/elY903AkUCusiUmADPP51AAOqiGlql14EhUo3VWXqRVD31EecaAfam9oB8H1QdUdtcHzO8
nXtvO3KYouKkNsf5pU3czkydQb5gE9ZFjn5qheh+PtIy1Iee4syAV8DQWMZqHWyQR0jlYCs4wkKf
Itw7oF2rzWVvjhzxtYYqzrQQYuAWQJK4jmUD3bWqWobfuhYw7YilmZ2Fj5aP9/V1NQZrVzsfkkOu
jfghrx4lcQprCXe2nE+V56WL179xFJShl0qEPRO/3VZSayzM7ZFrDqG+OMKGMYqjUtRz9hZubUO2
pp3pOkQsRXex+Fnpn0BOKhDQVll6taBkbeFjrIL7/KYRAc0MZ+hDUPQPqwsCYGTY0CdK0LZVbVuD
dUhvGFmTARxX82qWbszsB6ckQJvrj+ZlUYJXJO5wByJSUTA3seCGII0wAD2f44tBfPTs0cyFF5hy
s2VMD6bOZ32A+4fjm4sesHb6HFXQD2tqJLzKkNKwxkFKH1TVqeCA5UkgXt9amE+N7nDuGqrXKV68
lwxY2Wi7aSqyPeRQa3160AIUY/iKteIsAwSxfD/fZ0Wu/1A1/NL+9Dsz42Q9lLMkmPxP/iwcdcoy
fPahABEKBYN8a8gt632F6lMFrgP2CCXeVYXc+DfCyaqdkaDzcRjUGOCwFHlNy4ikKK9aY9/kHGZR
svCdUwUIlu8ouI3+fejGed1RR1W/kz5rsIGjerFFWoaxQ8WwvZ8g1A37fpam7aZkt3lNA9dU41CI
75vIlE06M4VpjR/LCCsbUfO+cy3f0jUq7g/4hHsFIAflrWqeg+djS4TXmFvgoTe7WuK7PCgTv8gq
KKE3N4edelSLV2ZsV2OolTx+Nkjevk+KAZyD+T6E2F+v6jURwwBe8TMCG84iG+whn+LvbHFcr2C9
PeSq9nrbvnskFnsM4Mk9VORQzXFaVfaYjTSjeBSWoEmahmWKW3OlCm6m778AQaB9+a8HnU5UEB9k
2Qu+t3wDPtZ3GsoGYgVSwpY6PGfdB2RLMEFwayTaszHUUbT+3F+ucQCHziYY+I71EybXTR43IAxv
C0pz7wVuyaquV1wsmrV1/wJGpMAAXs3nczJcQ4B8N6Fv7nh+r2xEqcmIUbp/bVpnHQQiIAMRyRfl
+R6Mv/HACKlmFAq6ThNQw7IH+gjuL3JTPZS3eEsXizqXQ5uEr+R6iy82XOvKBl1R6ufwViOF5Ait
aTk4ZdDICCBW/qO/vwFOVjrK5CxCWp6FeckxGi8qyr0xRv6jOGFTK3H2nxL0hYiaFOOwxxGRf/af
Jke4a4Pzmxji1iZm5BrzTyVB9mwTOTVfdaSV5ax7T4K32ixS5hSLSLIXH/CF3m22U2uOgIX/dWSx
vUEfR44Q3WF1akWTf2Nx3gSayxFPpuY7FVJcAH3PDn1gCM0d2MmSQOmuHbnXZjOZIHnEmjvyhRgj
TThnvT56GeerO94sMb37YRndkYo/H6hkADjO9cGl3aAJ4hTzpSq+zKd4GfiBi8xekWheUIO/qY3l
rFqdl2rF0OwYu4a+E3fGD4p651WXJfI7m6clN28YhL/rxhgeZzKFkMa8K0OadCEMb5P5W+cWv2y0
lUVcaSfksoiaHzNgtKzi3fRWSaZkXF0MpwBOfMn4cAzE6dtt4z3x1RoSvoTiHbegaELEo74BF1bq
Fq167gWQ6VHtGzHxTrLPpjE7HDkSoCljb6DYgrUj7AcWefTkkPa7zjcYJIf9gcFVQEljc0JDp0n4
uU62sxHhCEa5yklxUTn/8HTDfQVfSbHSQ2RpXDuokCAzSRgSmS0MC86HxW/P/7650MuLq9a1aaci
mAPncewzrqSUUDN2DUXT3DwaDVjQ52+aLSi4YN3MyryjSwgxvAqzCtNB5noT4lz7C6joLOd1QE2H
ECRG+OWC8z+VIQ4IKTmWyWV4UWXbqzU9zkA0iT5O1NCskmMHYYLs7TU4TsCED/vYKictiN+NOKiK
HP5GdRYXYi4b50ZndupCEMX+Su1wZddBeW8mWde4HsBakwWNzJxFs0XqO0cHrMXo8APg2LewG8zE
4aeEzXnV2yhAJ/mrvmVaAeOcVbYzviCVs1pVV7OfiKpteTeWcQnrII+RQNiWKqutfP5gk/wKj15p
ugUtd37fIDfxMnD7pzt/5GyO15WX4t6GSMPtE95KCbXrVpLnAh3viHXOKmy07kP6MGP0bFpAsYkc
ZEb250eV3BWAKO7Dl6XzBIkAgkYDFek9zlVKj6Omd7atjjCUPHb98qlNcwHe80bMq31h9m6kIng8
UMbydMvZe8q4xDYT7JWDbH5Q51N+8Hqz+3ONxcKWaZv+RuERiERY88cRz7BnRzTzWF9SJEB17uzi
v/HWjCipyr5mGt4BFdaZPzDJy4v+SUkGWvJ++hKUUK5Pz5G5djW0AjD/0LZDcHfUlWmEtnoJ4IM/
t5Ci25go3vUWkj6Lcw/oXqd68fVUW88F07z2L7YSX5hzmVBI1XYqrIqCH+yzE67SibUwlX86aNl2
b5EchNqc9/USjkOuFB757/erUwmzowFW67zIbyHEFIft7wN2KO6irBBvaaMZk5rZ1nJf+gKysUiU
qLH1Vx14zp2XFj0Z37tNUtTdWiD0X+UMJ1mkn9hmcFqDeXgdJbyIlpWKTcPl+R7p1rNs2WYn7flR
RStCRYVPAgSyrpCVKGmdclgVwFNDdKEXArp13hAkcKSE/Y2f3rTQGJj7y7cjydGm6+wCxTqPzXUC
PLR8XlvSuTBHAC5qoXME3ecdY3bTDUOnam/uBnMTkufGmC6G0exg33wy4euGPr0ejyzDgDwUCtX/
AZIQ/tBkHxEnjDeeM0y2cbxMtQWqPpDQAu8RQedtSPezbEJOicDymFC4WKDMlkldjHtGh9XdsKrn
/ScVWvo/uxPb2Uo0LTL8pCeOp+Q2jE4+vXoeMifnI8hNmRjApP6hQyxj2rknWnluB5KH0+qE8EWE
u5HaYRVr37ZpOC/zGAQVUIdhuqXbp4qqX+4df3H2rQe0KygsmJrsebBLFA5I+kNK6fOXEtF1DDf6
d6xdLbujGHpJ0rTssGiUM6f59q9MA9qkAZTaFrtJsx7IAZU+wnpP9X6tZZuYTRjY7fAtUUCXH5Vp
9ZszXdzItvQMWiS7b6jkJ2M2MOAiGFhCOqa8H2OZHsXt42AKolM7/mg6Wvi39uNRhLRSv+Dk2rTD
GUmafAb9xCZP6ghDLgTG6uZIe87QZ1ymIQRPM0D3qNSUKMFSUKZVDjYLGAIg1cyvhJC9jRpKsp2n
8v7xMs0DPnkaZkrXNU8Xx1YU7LKv7EPen58QMdT5uJu6C3bNrsQMWjwnQrH+QI5/NVQX4H7h7Rwq
Z5m66xLZXT6g9946zM1yF1KxENDZX0VPurSUEJ7b1fyi0pSpJ6ePhMljsFBn7rna33zUbCmhWl3N
BiLVZRJXi52wPUMNw6G6cX2aTaaXWoAaBa3VirYpKxSM7q4QZCecT4hoqrMy3Ph+4pduUZXtGF1j
jQVkX6sflr5AXpG1m+4K2MVLdKbkYol2fN4+U4QwzUiN9SJqvprDBZMBcDQgk6SlT14tGYlQGDrr
m0bLW8K+1NA0zkbRfLQZcr/ui5/d+6pCDP0yGobKJkinDoH7rL+5rrYXsQSati/X+OprTmpeyTK/
IX6CKY76d0z+OYnWNj3a3CWvW1KhgoPs9YgRh0OrYTgwgKyxAjLS0SgUBXkUj/OSIXSyanlzmfB+
2XEx7PEdSvYzqBNEbLQtt4F3IURMSHe/fFLqQyUE0dtYj4T6+xFLFxzCHFsYDNmWHBZycJZzw0Qt
pH6kYXoA/nJK4See1oAWivoDHq6t9tv/JI4NxorpKFelBd3E3czzr5wdo+5ZhDV1EDiaQDC7A5Ie
+F7fOfTNIE22NeWTWyy3tT1Rb/xWDoB0cnuJGRigdXeN0bIdinfqz59b7JvdukKesF6m2tCtgJrO
nYSI0hijKoRRUNdXGlLBj3X+YBUqlaBhKRhNef3oS3IrBq8BHESKORWvqyxwzFZcMgL9MAbSrfgy
uOcYp8XKf6at6zihVpRFaWb3hGwAJPlqw3Dw2KbnlbDmhQ+6xgcTBKtSX6qq8d08i8YaE4C42HO0
zkFCge0AmiYogsJx18OcPWqOz/UnYdYL+qSTAVMQrhv2Bz7e49e5T0s0GZw6+mOQSW1KOyOjLiJs
+qFSg+DXUwXCM8Zsts4ncuYR99R35mnYK4GxiOt3ZQ7KKqFryFEaL2etJbKhoi5EeUIfkuPtKxrz
cOT/te0Qun0qFLpqa/z3m8VcqIQ5XZOVqQG0bEbM8cDcYqka6TdSN0JmxWBFCBR+DS34bbi8iJ//
DxAi7JoWS6sgFIpHCfLwuk7Dae33nb/6Kr7+KYyWnFU8XrY3af7gwLsaex4vPdDLpiNnSmgKjAlI
IBcMmKrUp4drEc1maLJ2KMMsEt5a+o3EOGU2SnPMU5mFWhxUzfu569urn18tXV2PJbe4K0H457D6
wSNnAaa6PVf3RAfkyymzjInWXZ72EJ3yZzxI7kyrf6XIBujSioQ1nyhPZFLkzl3IddZb8UkH9Aut
xwW+5v5KdxprGb7EviBor6qP/6OVprwwK1H6kvER44uhEI/eFFg36F58TftqJ1rxs2jQ8ls9jpVT
sf23wQ1ZFdwV1TrZVDLv/ImUAZrygJHdn/jRgSDJi3fRJ+FhJqM2Ltfya7xIriNW5gzYU78C2Vu5
jqoE/vpfHhQdM8Q9G5tx3uQbqFiKhEPdxadGUg1f/v2x4a8nRUQRyhi+KyhzqD6mluPxWDsGE787
eQ0hEFpJbYV/aEyobT8iyECPrziG5qRjYjzWDMNrLkviOEIV83jyFxKfnvgTEvXjN5iw3E0cJTQq
dASd8fzXGyD4O2hL3XFvH7fVwe61r7RtEGYjmVp5mDRVkRxW5eJkuWrdj5+5MRWyfcjzynCIsQG7
fXkP9+SBHJD74TOtdqUGdsuHc6/9MxiXcachmkafNArGV/YFNxUsxW1RPrlsF1uov5kvuEOQ84gc
BZCZTdg009qWnayOuijYVrMEgWDJ9XTtNiQ22pFZf2StfA1CuJd9n1QaRHOlEKSHGOcmzQWX01Zb
/3ozc/EWPrtFhqZEttFJMlS20exbaO4J8uD9m+dR8EBaYIcltM8num9F4mRuEXrZThqWimG8jkN+
Q3OQrV0JqaIXODJAZIrRoKwPZ+vc12QIBGW3UWXupya+JlBYATvmkwHkeSUqyJGG17DRMRCkNP8W
6q75do35SWNDTDyoJx1BKz9AMkOR71NAOMHLsMLC2GpRfHJRKHinTlLKQZa110d2dKn1R+zG7SAc
DeshZlKHjdLziJvchfQGCa2hpc9CYcz8MknRsCv5ILLh9ckoilP3LoPkUutE7OdD74Wmyirxz/Eo
mMbR2M5PvezGYZD+JffT/NU9uCKC9BgrlS0iO8+DvlyR92SQheFO2VbbdDUIU5126C2hFQJ4qsUd
BB7iQagJIlNrfpl/DQTpN1nnwDrTOZtNWDDGKYOum9BQSz31tP3b242LXOHXWFlainSoj+a/YkOH
ETlZOHds57lNVIGUM67t9uSWHtFNyyEzxd01uomCOhSRhtOzBWVQtVCvsJCxZ9F1PngNakRfkbdx
r9zCeE603c/HWJWA8V5jIdQYot+m0xD9CPiDq62S7f2+l7uPkq9krfMhbbzZYY0qHunjSn5SvJzX
CUzQBs2USlZsXLYo13E4Fja0Bo6dtwBYke2fiZFSHk449bROKLyp1yjwPAayQacv4EuI5FJZmrRg
GyXOzYgDhpDfo9J3V/HZzUh4cHBrkO+my1LEggv/JF75wZaYArKzZgGjULXGGBc2h8uajO6VAplY
nZa5N4yWSgxAZ9ql+8SHn2cER6zam3XJqZ5iH/nNYiiy6MWMtiaozN/bnd1F0MemJ8if/Z3gzZkq
6Sq0ar3ZzgJbHmBu+njf9Nl07TYi6qaWX6DNrkML0xVMofEndyeLk8DpC4nqFM/z24ZgQp6sjeDT
rsIhSKtrUTcuucNRIT3yPtg/b4YAkjlWTx8oMCiv+3MJySPd3dEgW0TQ0uloOod3cuRcyUIjjhna
pg7NV9XqNnPIDtHKwBav2t1H/Ayk0DMpTH3rI8thKdm5XhWWjDpQCqWz6soaGqqTRr/aUcbXKEad
3ZFipxRne3q/ZPH2LGo966xd0fXwbPw0eEWlJTCDTGLFTeYCFptAUd+ofmOFojF/6dv7h8ohVQLz
I9u+M9Eyo96ZmabrxBtm2+D1fH5HOsfktcrYV6mbBNDGjGdfnRRgm72Xs1m9jiz2eisg29XTID6g
BwGySdfCGQbiAU9nwwl5U5qnGOcMqVHqZAPjPlxJPXKs07OpHhFO/bt1G6uWHOJTMX4VqCI1yIrq
373lh2ZMZ1ksCbeukNLRYq5ezeHR4Sw2hXaSOPeM2r6QxseIlVK7+3eASXT4v7mjR8cEXNt+nCp1
RWZcBAz4dUf1Wd1/DrjUuEK6pkgfu6GrvWtGhx1Nriy4VYdvwUnIt/s1A1N1BtfFWmV1E/DltvV/
GL3KXkfhpHW0diD626hRuGARQaxyDot+gJtnCc8d60ii1FIxs6kICGvrUiH9XzYIazNBErs5nmdg
97EfEwHt/gjz6OcXLRdGFeKY0ZuzXagh+P8DsmAn6xFTcVZRxh1pfdoV+iyXzASskamosVrSKil0
3C1X4Q1neIBt6dkh1s/rDbn5oLt4W/O2c4m+5etngTiCa3R4YMkqxTWLwme9gGbJr7jblzS7zDzE
jN4fFgHgI1oz4yjwMzinU9D9r90rwhi7pyNyAqAFD4n93xMm5nomxdPMJ3Z1w9WV9AfSm/pPcIXS
MBNYqQviqf53uDIp8vUs40W900tP7i10NbGdCBZtL8UoMGwA8qbGtnyGGmYpnaU29c/8u61zkNr2
0QLzDMoBv1EhVnmEOAW0j1t+02Y0u+youb3/G03kVzMGC3B1j3zFBEjLS1osW7FhO/pldnB8Clht
zLlG1ct5B1VJArsjoqUegpnQGcOulasdtMghmapasUhtetrKt4MunZ3MWEpwS0XDHsuVD6auYefm
zbHTuBEjvYOdesOE1SuIl3kr6YyNF76kosp7f/d9vpKEpR+uQLvnwDbWD+V3nhw+2/mQhWYJfXdq
vL7X1e4ytzOnog7JklqqPLsRHlbDnJThOJ/FEx2v9wqPzAQh3FKC/F5NP6O7hRRui6Vxd5fFNhqE
x0trySxxt3PFwf58w52+Z7JLkgWfWLK/bta63mYBpZcWZXwCVlTLo8GdNTuxPsxLNyP8TjaOc5Y7
yPviD6FaUxGJKok4eRjMmDn2AdIbGXAzzjFH791LqxqWk9d07pvgMVoVOfxw0j3V2dnXziCYRzMH
rMUBq5ibYZWD6g64oQ70eGM7dbXBl8v+OFTwVN2ZCMXYRh0AKEGmZdvczJ71YPdUTSwwJ1XBRowP
KfyoGy1iIqs2yjojUmlnw6r/akvitN1oVe/XTZm8eERunnTzONDCGTtUneED937ISjTxu3AtuLSY
mJ1NePjN/lORg254Qjr7DxfECEomldknQNf03/eBcNBo9IKp/kMgZ44E0J2kyAU7FwX9wa0ibM92
2zktkjQJPj5Qw15sFZ8kDG7zqGqqtQpMW/uT5e+TEtvD8YX7Wcu4sKol7U449U4TL05gIbXr7uDq
7DrHzfYqycIJscGBN2cVDh4WPQYythTWXEmkZGsnzBYZKzxZkmsg174Yz6AEMGhe90gJpPaSFjcl
Ikjm+YNei7EonkAEcmXUEZirD0yVhRlfg88MJ1jkD4jShrSn2ISzK3JijZjTkDMx1/yhfy2x4u80
bMf585A0vt07qv7Q5ZpiBRHmmuRY1yrNw+mF0Qes2TAUOvuqQZ9S4LFmfuiUA47wDAGGMQjCLHTS
5wnyUgJlBmiECBzQmcXVUcJQkvm6Aizag/Cki83FJR0lKJoJ34U6nlkMDFXWB25cb2OSiZBF2Wqf
Kb2S3omaWBZAXx9P6tH00QBw5AFxO2WzOx/7dzj9N7E948EV+v2a7aIrmlkYlfg4RY48a1cm1gZD
xcxeVDI0Urb64HjsJGWauE0uMxm3899Ym9iic/vUsN5bSYveDAaB7t0WwgM9hnAZhRhKQfZuEe87
0cSLtaJS8gi6+AKyweSaRJEt8pwbFTvi6GKIc753QETIAbwLhYTSfb+9guxcY+BogHrjZPYYhvNF
CIOsJRs6rNPKQ9IIREh02W1ijDjSK7o4cpFNqrbidH8aHJAU92XxG52yPGCp8bs76Np9yAvsjdOe
5OULKPw2snTHtZBvvszqJsPvW0DJd0r5CqQQ6+0MUQeZOvPqtWB50BQHfJtKhOMxHp2zonR3f6aR
UyPBI+qZ0DENZRflNRScQVsYSnNOCq+aKkQKrrlNXx5fju03Vghqm0DkbelZYJLFSucUV73UhNhC
LKEc/1+XTZ0nXlryDhI+e9Ox2G8P0JeWnBKMppxwPuW/4KXy2LaBH5Bz/Q1aC43aN61MKrfIAIUq
X0O1DaaqzrACG0CNpbXMH7BCTrOQWCnGx3fz9ZKtiaP22H8mGl3jpH49SvQqyb9JmYIld3Rg9x3J
Lb5MSs4uqsHCpPeHR1vW/zvAwZlDTDjDpkwzsDFkO6pA6tFTLy8KAjbJ488uYWE+nZEA5TruLcN8
HM2Xhc6/dktJkIlKJWIKgAc9qNzNtz0C9iSGIeB10XLC63GinBxnr4FzORBRFbv9DgNDAtIb/FST
l4Lz5l9A29CzMLiCLJYwR1VyF39ItFpzrJYHbOopNgXWUie6bkBkIKms/9ORIBSNGGj0OzDiab8a
T4iNP900vWPjGFANx/8Ljgc6pR5h/J143bOn/jwRFs81X/R6560aINzVHirSk2w0RT11+dPTaCj3
9tEIS0HLr2D6s9RkrPUy76R5irDmVyouw+fJ66a9q9c6sw9R1zUu/mvnSkyk8y4nrunkTS0mjNS/
84jjKV6M+Jmqba/HpxWq7dEIz9HfshIJZKPFzg/zF/EosFGtgaFFOhLLe/Cj4EqAoEvRKkrsMmrC
z/XhHBtp9b3wVD2g+F9w8az4NK+vOeW/DTveXekgkHt4jWeOyJ6iFYOnrMrlT3i/2P69+SX89t1P
+cZ6dbgz4/Mqwjno7au6TLk6L/2g5cjT6WXgw8i8DQwomuMoW3IYBTBof3TSCfmj4MNmxYPW+WCi
vDr3K8/gphUAbfsOI4cuzYuqeEk1jQCm184aQTbTGdsttD2jXazZRDm2sI+kEE9njjdcpPrieQE/
z2lEq665MvD5v/mfzF2NIKvSsmtraR3e7sGVxAJqGIAKhM5l67/EzRerprMIjmlSD/JgkQbNPq/J
0ob7mFEVSwYRnj5e+xdTKk6wsH3d8UyjCcg7vCRMPZz4o+ABk8NcWH1Z0wxsdrkQL2I45VwiwfPj
Lbuki2RfHBrkNVxSNN1TO5FbED1feSlbTunnXsXw16G4Tv44qWXkGVTSH0WTT66gcTwzlefISJoy
sMg+HEM7DBYfytu1Y9htYI/XzlDlp2d8TgOSglK8eF0xT8Mm9pq4Zr5UE2s8vBR1G8DQp4aWrlAg
rD6aAacAlsPcZp/OpaxV8Ni5IQPLZu2pr+MhiznIOluk/6u05k97/EvRnBk3zFBTf9kUX4WYURAb
Cy8ZpS8Gy0ObcEPPfkWzQk4+g5IA88Gv37QXHXecBqMnU18b0bDUOFKEMzKRzrYQGHCISnwNl2vG
saOvYuzxzd0b2ErFxJqL9kd2qvyKzVYj/p3P4rLjw869/OZRPfEufodgl7zcsShzO+ZLUKGOUdf2
lLTpjDk2tfQLjwVgPoM5fsNeI3ibK6pCOHPJYfmh4sYjvXEpwSXhRsa1WpM4MZOci91t8KlY2I2N
BN2Qv8q2c//mI7pST2vZbZ8BOe+ZHHLMafzHPL1t/L7dUyhLUEFGbs99GGw2X3RJ9/Qz570QTHtY
kp73ir8TGWWIBJH5h+PbTqFQ6Ahx8Grht7BbUHV1syz7uGdzHJ9EMmaqzcrXMyuzDKW19CMbLCx9
Qg5c93PL/t+ao66sgPLDsfhPy0Sm3ZqWElQ0Hx0aRM75IjkzuDHAVcVvt67+7jraiv5B/X3tiK0I
+AZWDsFpMNb8dnBZ/meg/xq6mTKy1k/gNhYfZRSjqDgAx/WJ5CUTOppLowxgpQcjW/huWjt0/MX6
VOFf04Gn3YeJ4b17hU2bn5P/xzCH1pkzrIOrnPLX1b4oV9eITnECNsniyLoDSffLXSbdbt5NTQR5
RHCX5b6uGwH+oOMFq1RCJ6E2enD2VKZzDd0zYOWZU6oaxlhnu91N5izsUMYm0DiqtAE/XmEQidCE
yIlug1/kYgIcIjDLw3glid6HmaZRWUT0PMn9JfuRwHJ5nk/gQboACI2122mQ/EyX182Fu0D+D4U9
TxFcHAKZ80P6ngh3gWkZy1JmkxrerTwnDIMrYL1XNxWKZBqhLCFMeYsW8/BZ33NJqscDa21sYRxN
xzXuoTqGFxPbjNj3mHh4W/XcapyzOJAWAz/ovE0/esjZhx82p3L7Ww1tK/idQ5k3WqZ9r9MsTBpq
gxey1mjnvwvuWP3VbQE9QtBxeFjHZWPQiOBnF4FVAmZJ2YO6QYsHswAkW8wsRX8cB1Tuahltk1Fj
beSx7Rpjtm05TsbmrfPYWv1x/jMLNqZp5dDnEedkVUbThnPIULq/b9zBjd9hf2r1wxCGcYj5OzrL
u6sI74FHjsqqx5KjKVMgk8ycZiUlP5CW/h57yyOTYuG+zbJNJrD9ZAqlTrMmNGeTPA0KOXlVokyK
fUd05gV6cUuaF+I2e4f3lKiqBtzuMAIDo/sPkx4r2TfbNiHwFWiQP6eYDn97PtQC6juzaGusKA5Z
A3blegSeY3fPOsR5J+l7dboxUw5UN8EvBAaTzHTkrv4lfjvReg9q2CR2ERrYHlve5sJ3r3MjqjYW
XREVqjE9ANDZxGUQv9U/KRrJnoZmpNgVMKEkF/nosQ2AMMWasr4bKC5ypuc7mu/yUJcd7VBs/Rc7
IhCJCeagxO90Jg5TW/29kBwseGZq90gdY7s4AZ60bgykX7mA3l48Fp9FyMJ4+LVfrhsiuNPOR9gk
udSpG4Qonftj00Ee4RkuKAvgwl12gOYEM/vyBhUg/jdWyFzkHiYCHT/lNyfH08VoMBtURB8HetsB
jsksRD44nBxTSeyRAmlXG8PnA4sqNg+9/sfBEqLAnluvcHO7YqGCF4k9eedLCbJ4ZZT5n1Q50UqB
8fBPnXjcc6/Ht7hm1+RTQIJOspm6OE47gJeDqPOjyGhCIQffBXTHmg3aBG3jFxEm+dpzRcaEeDrs
MUuGSfR8YbtGgdqhXV9EscbwUckCgur9OwLfu1UiV0hXMc9aQXVu1YKQRI8yEi+JPe8HWqksRk/9
4cB21U6c1WSsNKCRt71ByKYgcJUWztq8AOYACNO+9jQzabMy4gHBMh6bXUIH6lxDCoMFTnrbrERb
NbEqsVMtNcP8vplaXNfz8W2rtT9WrWUc/CoE7jpxG8qB9sOwIhSDCrYGn4o/T25h+5m3W9FDztqi
PEzg2M9bodzpbLH1mvneuqerjy5wlDxNf2bBi/2QbQlZ6cd45v/3Yeev6YULisCzrvONI2OJNyEe
hT0aGlfCYZB0rvHTLK/opP3AlBKqe1QFL07qf+8WnkEL/QnTDI0PR/JeBZ1lkHt9sRZsOkbhka10
bN64iX4XwfIiqA+QJ2qbUkUL+BkdzDsAz6nx1yV4+AS3Mh92trwm5oN6cTXlALYXtxenzErnaPpD
lhduI3n2j36onC3Esw+nZwXRWWMgP8tBhv0gPcg8oyscOoDC28FZJEgqg4m1MHYKOO969OZBaI8r
7ZEYDBRyf1Z+p0sYiUQGirB+gCMMS+eWJR86YAIMnZCKWClNa0duq2ES0Ai5gObRDo4uZx2j0alm
0/dSS1rBTPXMgaI6o+pGhDoaUFQWxPf7Ib8c0zEIdnttpi+m31JaDbFSkI6W4hsCQcljwSGFioat
NxwWsmaA6mNuv+zoY5yfMwocawOy+b25uL+L9K4yD3LvUjLWuQ5Nw2vU9o/b9Z06dX6yJSnPMxQh
ZpmXq4XynYMlL4WxB/OPlxgLBndwr4rgfCbso/i7Ut5Ae5FKjKx3UlDyUwcjAvD3kpcPlIl+g1vW
7bMIDNJzz4Dqv0sTcNFo0bE05KDkHQYab8QWfVOaFBGgbJ1sWs25Flpekbc2iXHoYZA9r1r4u44f
dZLtsGwmi9FebsqRrkvAuXuhCNBa0OwkD79aqQpRQD01cUOYFigT9ykYSKp5lczJSt9H8Ki6IUU4
lEXJub/cgvNDYp6j7hAl927jwkd5uT93x1LFGP+4vo1YYRm+OptrdZI4HUigWbRNEzbnocQzo6NC
5nbrpGCVuH0a84Si/DjAeH2uGLmDmr0Q2oKXf+1D/4ABd8+ayTYUBaCAIs1TDPqLjy4f9M1Joj7s
HBG1DLyE9lSQSifY53lbIstZdtV8AD92KV1IsnK27rlY+/ehS3zHLMra1vA40SpeW5dwhRocHZtT
xCjMHa05cp2im4QEzYB+EoMuwd3JODgS0GlSNYs+ErKtMB6DGJS4dCn69Er82cKhhzLQ2tmDRbmH
nDPAZVrIj0skyqzWsGK/YMtTytxLgdjztkkx61s3ilM7mrnWedFnYOPXL553FjsY4OZuDx0B3H49
kS2AQjlcTMN8WMmnxSox7yvkK9SdACYARUdMO5QswHSum5NoNvAhch+8L12eTQGRbZG1mSXP3Our
fkOHhE/3UBfavBs3cVwQKvb0mwkEqGP00DK4XaKi1ZclwmTK2/2mulbhndNOQAPsf6zEAw/g9RgH
j7nohKmyHvejmMQple+6UUlU3+ShUOBGnEJ2M9TlaFHJeF/6Fn7PvYyBTWRo2wEF+eBRxictmaWr
xbZH5Uu5lNxsxDvkeNk51VMYRUsv0eXmJG4LkXg0EPg8LP0e7hpiFXVdERShjKsKwkoVpM0O3jFA
w9FwhEu5HcKDlcXSuanJDq5pjVWNYRDfh887bQ1kmsjdPnwbnCOxLSi/TEY28HR/nqCnhiOIkpNT
n05fkjdU7XwZgqAEv4n7DUYyMxYjstDqmWbQSBV2im/UY4PmTFzRNeTMGuawNLx5B3Lfi3d8qDsu
evquONCMMb2GrugpcBF82v1CzbmqAvmLjNz8ZLQmEky/y1VdRY4w7PlsvU9rjMJGXdIWoK5rC8Cv
mWBor07GhlRQCZC1p+wwxB4Biwllc5dBd6nXnvMLNgToC4I4F4OgRktpeDQ5oTJDKn2LRKs+y5Pe
BzlMho/FtEEj31nZnwq8/tpdlPGf+/Cm3+lNWOiJ6NsMTamyEFxPFLYUjouwl7hlq8UQctM9t/4T
kSdK4ORaELW4HDcI+/MAgN9Mwe2ZjWV7Uhb592udwQ5xqmzFNnmytQVAIXRZlQ0pb0gkrlaiF1m0
fFRM7ItiCJAR4e5bGZk+kpXkQOCa8zaBSpYToiJcBU4hJYrUjS4cDBdqG5CjIospPlJ9d3MKnK63
OpsF86ehTBMyWypOFXa0+40+w0TuR8V0aQkMdRDHsLsMnZTrNGvqvBnV+572V6XKJL/tWLs2SUVv
jThGcQCmanWaHM3riyOzsHhzraVezWxdS4G08rjQqy1O4tUE3JA4h73zz/rgymLqMN67kc+oxzw5
BNU78BAg7vY0rKS/vYuGVnvMICBhSTzpZ0bUqWUuJ8YCWyxe7OYrIKrdE3EqZaQjDAeznmWkBhVn
11g2vsRlnBpG8z7s8y/J18I4AiZDlTGxInsr0w3XNpLn3ghcKOYBYPZsXpcFQV+tr6rkg4AVVUgW
vehwnkH5bM92T0lpXiZRT121YA+9CB+dMslgVE0F+PmjKalnCBPXOsuIRx9O7AIt3xGEzkV4cOVN
YwQ06AKQ5E6BaErLn2zp6SPhJ1c4/bqtvYvjIdoiIJ2i2tuMRTO6HPcz+GFMEqwZ7xx1Z4kPXqBI
1+gdWJ+rDkTZ23/6uIx/cGZkCXiZcYGv3mnbRfi6hXLjb8874KsXFqtytJ4c4YB2uxB+RSkp1Fa8
utDcf9AQAvC1v8HovgwMYnFNsi6wuAIkP0dfYnsGOBgdrC+n7c1UF8AMRDyapGbmsA0b2Zqr8UPE
+A+sQ7bhPJ4yn3aEp1gq2lc6Tedb7rJAzoS5vnVv8MKkMvMPG6o2MnQrJqQCMaUyMQcbk9CntJdr
/ACegHMe29dm277spWWIqVJ0T1PNUzN7lBzHl9VKhIPaCZ6+mhI/UHPvWfrUfjQLw+rt73FIYBZ7
A4pbve75xq6MUxrk/TdXw/Xz7LcAwp26NpDlAalTZ879aM2kKGXVbUp8zAs+CDpzHgnudLEqQQUA
ZlXNCudukdHhfe8BaIk//ajVVd1wQw1PICrMuX8Uk8VzRb7896jBUPyLm+Y4qZdsMjcBHv6gk795
jl5Vh2KBA9vWeqyvTni5TFPLnglFFY0Sn7ia/hujSuciK9jBUuAkJ22ZzyM3FMkhNtoGckB+nDwU
TqrIZ6pVFOjNuE9jL5UtX+d9+ksaT/8ubh83e43XTkuL1hHvSdNX+ooe8ITZcOnFh5Isd7Xybu1c
NzzfWEKxyCK/nQyxWVW0puHVQmmEHPredJMeXheLbNq7ZaM4A8odOGQXDv3NPp/NKId2pharo75q
Y8HrzYDNTYWLRNWruTKxz3IdW0oy+g1z5M7U5GV5YOFhxHwnH1SteCSSWE3gq63eEVMb3Xs2lvgj
P1geFYl2xggcqI+mT8/2/U0MVwjRtN3fr4TfXGt+1EH//KaK7hp3BsciErsHEgptrAlySLkS60gZ
sZcbvkkKLSU38smLtLlds/7JAt7KPjqsPzhZ04B3bqnGrsnu7OLin73cyZjzfd0ld3Nx8IRsql4o
gOHvJCbtZnDfwTUBJE/w0a9Kw/JrxkTlmLriLaR7fEyHZbDG3OLOrvhZWKhoYcbfhyWe+jc1TwhV
AJxHZQWp5aEwrtbmrHeBUfvYsQ4RCh8m2u/xHoA10FnfkszhZipXBvBw8074ukZYC+VCJM8ojeAz
mhrYcN1AD5zl5JKVJhykE/YZQXgdMMFZ9GTyte4uJ7XvLqPrx8gkEu0OJtEcMUpL5RVdMAsNStHN
bCyDb0zIUONQxnaKEE6frk5lSGCS+fXqiXrayRgGY3+qPVt7qw7X1YUicLwHPGJz1P/ZHoLRq36i
vbEtqCBXK+L1Bl3cF6rfffKKjvKywPYSu7wN7kf1VG7GjevD8M9JQ0S3+d/Ay0+FiBzXf3uWBl7V
OdW7++a0EChaUqSyTbBAFkD9/HouV1lc2EU785gHtjZFNn/M6Outjwo35qRHIlmgEiVnHw/TUVFs
KS6eShCJ/UR0F8JbZU3m47pTFB/jwXJPb9BSqI8c/kWPhZoA2nGgi5vQ28adR/yxRREAEG80nbYP
cKf7Pyg+O3OvcRnFFqMU67wPZspww/kfXQj/nYdzUCzxOuVM02v61FmAqKAXR11sxCCWdE8rDHwd
0dZpqnpoRVRyaVrlv8S8/i0GiZpwpbMybDJc7QI1ikQXhrZ790LakoBL0bvawfmClyc2eXv2NtJQ
MTyOgB5Rt2RS6ga+c0qQJHrREct9m8kxEzDEPy0bpVx10LUAPoBoz12d37ZnMVwsecj4x9K2JWK2
6xfD5PprSqbnnF//VDONeZ28WDffg8DIgap/7osu78WX8g4tUysD+SuXcRx/64Hql50FNvoWYsnM
gWOpGttC8MyZKsugsIspsMTgMJvl6xEhC6WD5aKv7Fnzy/VBjGBtE+M1kgHiq6j//pCCv7xp1rio
RWsxxJQ7d8rCLLxml5Sj4qR4PO3AkhnsdTMm3HoU/1cdFlASsVTaRXsVBW+Iif5AODB/CQyUr5Wb
3RXxQgWA6u46iXsUo98cjv+zEl0FN6xjS4oBtBsoC4l9qdC3LcQHSHFtblJd5XqRa4uBhpc8eQ54
VBRnOyzaoqIuCFMs97NFw6N9QM4uOuMLFUU3m2oz6VA21E+LBfh6igWGzKrvDCMzuEvYPSwZ++pG
19xAcfmksm7hGvKCsiV6atr7ZC8W9Vw2pi2YiyPpS3Xt5YoBP1SAWu346bFDHspQRn56hbJgotSB
WmzDrU1KTucL0JTzmXbUzKYHZqYBYLVxR3Q1C0kfU1GIAsCrWCtQsMN1joUhhyUOshv9J5Q6xqn3
pmDKjGy/iCW/xKB4QOIZPnbrXnK7BanZCxBLJkVHl9GMrYPgcCaeH8gvIqgW4WxeydLHN3CM+B2E
CLCPhp8NcJDDvDYs1PZPWquDyLrmszibVJ3Oc3mzRnJ8xbJNtktGaoQlvA1C4sx6/3e+VgEMfM3D
lQczH9VeCJiyuRoC2twhBhnGP2WwP2uYNO9g2T+m5bPoGa6YmtvlX+h+o+NrBVhA1+ZParZBC+i1
pmzRPopT8Bg8qc34LK3ggM0rzUzS85F18Dwb5LsM8KFzs4mSVJX+MUdbOGEy/GFalA/0262M5hzD
gGw66KKDCLl5pUhQL6UGSkkUilPnlTRlhit7CGJYirkN3SL16cNAnR6capL76ehOdAxqPrCiCvgn
IxHboS4loT6x82YtO2xXYTo9DeDp99w69PcnCZilRdGEsGR2SVHbLgsJRISENmW5PRGOa5ScnZ1A
8yHJg2+gNyGde15IUlNbU0plncAlNKvqqebXlMjIEhdIJ+WcByiWsG2sJLSfLTqKT+ZVDUh33EiH
MoFD9Cc3k0HYKISuXbyVJe75zWUvDtELSFWKg//U1jsH49xBuxgwGaL9SBLeLRKVdfdOT/YWzmQ5
Zr6Ep25I7NA+oOdUEDrjJu/bvKwRoLerWgSCmqA40yfq96NF+TSV8Vi7ZhI0a0bo+PPPgi0TR+Xt
BZ7iLhw/PCELRPYxe4pMyq33McgYd7oQrKQp06DvlOX5o7WMJVmLy9mkGJLu91To0NSSdxmY011V
XLZApvCC2/02oSWq8u9SfXQJeGDVo8/Lsd8ux1BLUSasVlrIYGYAszo0cQEWJEMyBZKPWP0ItMPd
a5QKLN1VS0gjcoGOECzA/hkWMGyiVl2Z+MmjavZOLwc3MkVjAZgKME0iClke8nKZQ7Lv/mpmSEkt
daqoAXsK8GWTSq7BDa55oGLMTpkGF25DzE6Ob0ER0Ntg+KUuESmwHZQweaUtqp2DjVhnN7MpZYA1
tb7ZQDqCdtCAEEiR2OfTRrgXypv04VC7abdWQdnUBjL2yVvb1qovS5Pxc7rvI61a9Rb9TjyqSLuK
OFrlIpPgMezBnNGiKkxi+V0thpntb46xHwjfSSSGJtDIQwr+e8V1w9n3aqhkJp86hyCC1mhQI+dU
PxoPOqMdj/W2UoIaiwijaseCCM5pF7b3YKIHUPd0tXwEq1iOpxI1/QxWsFyPRpnZU8zZjCyGsyD3
EqnumX+1/HnuFRsnz6UDZf6GubbD4L3wWjkaTs4pupa9NXea8LgMIkWL4dFXMIt76o7u+LZC/kJN
kFqIUKxrZ2Fn0jHJmqDJTMeF1slm6Rn9xJRJGtsVbf7ELRCs+fHVloDh9kR8QHcVJ2DmJkqjOF7q
0gewvoxRUhVabjNs7bhA8B7V2USMBUEZ8n2SjwnfFmLx9XSk37jZatKVdyuIR3wLkbg0+/11rvQr
Ko0C0j1j64N6qovBAids/oH5bkbLYP37yvw2bWaWqndAn93X6vnUN3fuZG6Hka7u3jgAUaSpW+w0
4a/SI06BS3eCHmk43aHKbrCDcFVsh/bz2V9yFULuo/kIIG20a+P8vkH65V620luh3cmUjHVfrgc/
kSGCjgwz6pRkwPXs6fy1XR7RvQnU8g24O8UZIo6TzSdvst+DYk+LXG4PW96KG7BzW9yGBGvm7dk0
7CYke0avH/1e3y1SE/IhsVuCwVl5f5JpAv9X8SAqK1utx7A+cC5rqnrODvBvOrYdEwVlp2jZjJMn
4B1vo10d/Z1zSACbJvzmtGjtW3gtQjDezF9s+gWFB5MX37Tp6E/aPelqPf3JW76l6s9KYUCxiS+I
nFr3LRi0V+q/ihbrFwZyWBizUhIspVLKVsQXICmDSV0G9FhREEcxqia3hQLKjGGefG1m48SoqI2F
Fl7r0R733pm1zcForXHMd+7blDwJfVKA6ucDwLcYMKRnStsjjDXo28aLbPvXwEXlWDqGYMgYf+AF
1yL/ONPAksCqV9eWp4RgCTadDrWhs5LQQ4mLDVm5pJ+RDgkbFbxx9gBe/O5nXBNZD9TvIBxb0lpO
hOnkHSk2RMD8e+lBLQf1xh6Yn1iII5uk7sj/SoOpe2UgMpXPT8URAf7wNcqW4d9vu3mzzS8zHdbz
ehOPTmQ7W2NK3Q79aBzXZoBdMEiNdFSdLZSROpxlNPKNCS7JraZ+GM1Fz8us+3BV6r4jmSHU6gFz
pfZFxoZ5Y1X3mfNKL8cWXHfk7aXv1b7Zbenjks6NSzPRUpj0CTDoIT8hv5eichft8rTj7XnFZ7do
WwGEavcLNPMHG8rvuGXFyOoYoLIB9nAhXJLEs/5dsUawj3wR839HjHoz8bO/go7JJAyb8yEP3cfG
Px8345eY1ZVXwB3RozDGwafN024Kk5gZ4PvuuKfIkr0E59q4DOoZFHQwFTSfldjE4Fqzez0xOpEC
ZGgEtqE0AuB0mHf0Fj0qo7WjCdUTpha6fqTjVHmDCmQDzp8bRuhqJAABc8YID0Z9bW/wsfEWAWvm
dnsbUdlKQRc4GSjJM21HREL1tFmsES5BiXQhpPEjA7FEYR/IxWXHTKy5s6uzOK8e320GtprmK7H/
aNY2m9VmwjAB0TmL6h6mqfQbdQ7r0kGQ7hWy/J/XRTR1FickgABPwT9rXz9x/3y2tP65v47xuK7f
1cvg/vmS9OWSPEBuGiKPFdNSAqhgGIXnOGFyiG4DSLBinPr+u+JgNbH5m7WnJa8Es07mty9UmXS1
oTHwi0FG8TQilhypeHhBkZCWxKLC5IGkbiECdxIJfG3Z9PDEhie67Bnydz1xGL3xS19cExrONLYG
5DBF18YjL8SUhIx0SnH9/85EG7t7xfPyfQOFBR3JNYdQQfn2dlehW9IpMMvwqtpoLwvlZzafuVGs
CkoA3f5LC1MCdDAR27CrK8lysbI8ZbikCry14ufRx0mmzc6XSvC//NDfKjj75pIjtyMnrjdYWRXt
ezEv/UrBMR9MrShSoIHeIZtG5ApFXc+xWAaxeVsEMBgWFzIDAL0TKm5YZoQCJmtef7rL5xr/lLm5
k+3e3JuYbAOBrNF7FMLuEJgO8MLRtR75E+d4RJZM1/KSSpXCaDb2ews+kMB2rBCve7jMEUH3x1vc
SnJtt4d4yqA04Ld7fM29NSReMJmcO+5lY2LqF4Bf+k1RhIGXNmK3D973kP1O+Z5+AFPTmCZZG7Wo
7JFKGQCwl98AZiTF4UeAWqsrXEPE86OMxEemcgVOWGmBjU1QdKo2Awbr2LiCL9pVSrzAP6tywusu
vDAaueSvcc8QqSEtdgb3hJtz65vQuoK58LK6nzhyd40VDrja4xoAyIIwrsoOpKXCnKt+rw+S6l2M
IlzdLTOZPDLdY96B6xw5FitKEdv9UjaKo4bEkC1St0RxbOKjG8K4crwijSiHSPiKc8wi1WMu2fdA
okVJfJRGccE1WeT7M3wxbviAKfarqQ69CIKiE4acR/afoFPGH4WHokvu89JfOR8ucUO0epU7YtMp
ZPo0twwmeHQ+mfLCkQ+nseLLa/PZ3bFTdbmClJaamqR+XEoj52rV1N5ksKsKc7+HfvIYNfEjHfF2
2BcOH6qaCaFksYQ5nb2DIINeFrfI/+AGQJeEbdqZvjWKTzKO/QE9+vgChlYknH7HBczQ++qWIHwx
OMrxTkPu3mNj1lfDJkoAbOD3p3xYqsDpCnjm5Micgy3Yi4ejrH2C4/RCg8WNvagAAI0lJ4w+/LrC
ZXEPaSZwGIPSxQScRZnNLQYy0o0411QgK0Afoh0eScfE/e1JDZvHhS74Cvi/MhWQOMKLfkJtGJ5t
UBbP7v1np80NA2j8JMEQvBDHd5Q2B8GexRgxnpk1TBODvWK98TKK06s8tNygHOKZ59uWU1ejtP6H
pYI+BVkHBOarhZUo/dp1dKirYRIXkgAFUwNuc78+8PEVZedFfI8iBWHkr8Sl5NhAUIyo/V0wQbyO
pevrjF/4fLbXKDaxtA2vIARqzOFKaoqfIZGzu8nuOHfeiysc0WZUmPSZ+P3eeYAv9mkeUf4T5imM
eNpzP6HN0g2yIJc+pXOV/0cmKUnS/J4lek2R4vgoa3QFC971YEqAGcrDv0yZCxJRtAASnYn6tGYI
UmHMsvuQoHcT+Rj/ry9GSNuAHvC66/RmwSYHdeOOe4UbuEDdIWLg4cRMsJTLgqV2RRv5x3TsqfEd
PwVJJWZsEHB4wdWpu/GWSaWBOZDLREbjxCgOMSA9B9uhdFk4GSm5cmEUaXKie2t2TQJmFRMnKjJD
IZld3PN+VVduvc7wA8a84+/JK72qkL0gqKa/Y7d1tuuUmk/okgaGl7vafTBF5BnXoBiWP7DBmf2/
x7n60ycxgiunHeYEkjNp3AGo6/sdOexNDJ1ma0CUKfmO87GO93S1M8WEmn65dzJpMzblWoR/pdtQ
Wpc56UPl4adKWcYWPcZ3uqFF5eI5b1TaEgf+4H3OLpwe+JtIcTqxkeoXGWLjG05oHzrH9Jd+gNeQ
hxJVUd2VHs7X4AydY9kvoyHi9u4mVyqwwLyo3Y+xhBeu+8bL25SDPfNKPhDbFQ0LWxBbROuNmNqf
eIHIB3uLnkQtEz8H71tZoq8SWJmBdpPYJgCHFsldwTYI8JdxvGZtcA3yWfVmohoxX0ZloExSrQSh
eDbAWclDJQFVht5tCiBPSYc49qzAY4F9Idd86b8TLneZsYTJYMqWYyKHAeEFjmGk+OLu4Lp6EKH3
cm3J/SJJuHUD/LMrtoBFxhsv2+pF6CsM394mXHCrYjjF1x/Xs4rPchAXOjw1HhSoN6lJXvJrF8vW
3E8Sb8ZhH8dNzNsGbDa738acIwj0KLq0iB16FvT/kWMsqTX2mCn8nSDifFh8Q++PhH2LZna7Xkmp
N1DjS4RRVeCuBSUJkwaRanDaz9cZLxskffU0Kc2pVLdmgwQ371+uXjVQGN+JojaJrNQ2DABTBJu1
o/mxj3/SRIQLd2Ea3J3vVNgDOhjkecrY2qF069xV8E9MaRE61PeEUKkJgLeWbvob2KPWXAAzMkqC
5s6W2IotfCEEE7mxSIj/sQYjbLPe+4qib+LZ5Vv8wAJrktgD/MVxqVWRswY2M4+bplxJL+Vbg0Ww
PV/9YVFAlGby+7ACJO3WKoSxLHQ6RoRkwOfjuIu0pt6KgTKaNMFc1RDVDdwPfGrT74EjH4ye09sC
WhzNltHDd+T3nkDc8KNWZzbdFXGNtB9njd9hnRGSwu/cE+OqALTvRCowfjsE2V8IwNiAnTHFl77m
0k4eN4vzY4J2xfwfk3PsK5mgsEDTG8hj858ifX1irXIMj/5cJQDkNBlwbGmgNIvHu1rBdjgYlK5h
CEECNcTkK8eqY9d8gHBO4PsxlczmqAl/wU5hD+UV6eZnueZcjzNN+OAa/0yHTqAChjGHon85E8N/
T89PWzV2si9GfNWl+4sulz3qOvo0qIcqjmMyw5zn3ri5newMEY0UAU9yVS+gfQpMd85Zrcyho8cH
dIQGOLVZZGaxAfXwOE5LifLt8pGU28QkI2CBtdjlviyc2JhUTeFg0XMX3y61wavmkkNYyYW+FWZZ
Ind6VcI5a5cm+HW/pboplftiyzm64ezEtvapCAcSzS6Wvg11OFKouULj8Lmr9Uzm0hS95sUTCBaJ
uQ7xvZcYI2x5Wsr0GV34Aj+UVpqBXvMvhxpGo9GOdr4Vrlm7/q/dr7A4AZVRWATXNmbXahpDbZX3
FeRHRvaJ6+r2WobGMcB2soWn2U/ykwh831ymJfIK0DQuBO9SthiOSRQA4EneDpRdqpNEGuodiEhy
/ksDTS48EbRd/FBNaYCjExX5uJnx+vAZE7e/h9wuL9QBD7TaCK3TeqWcDAjpXa2qpHOsCbHVNsBI
TEN4qNweTB8wDZo+6UNXauOUVRJaAchy9ZQzwV39Fnm2qfHaYMqGYl/MV5WnnCRdBX3XaGMq39nA
GnjRbV8mMw/qD5rrc/Vq4HlSOX7Jlnv+NaX/MKdz15FuLw8nLU0neh2oA3C45kTJo9SXZ5AxvNiv
7tyKDSbeb+4P/X544EBIpFSoFDjXHSciXC0gsXwp9qWq+I8n+qNVR8yVtArkN4XJqBynZodpWhBN
f6vXhsZgpPCi7R+pD2VC1KZXIkRDpLEwoKY1SMrfEUON26nf/Dnus362pmVxPDvTcKVsfS7hyeti
IcmsNWQYIgE9r/lX17D1RQ8LpIlnLS9GY3JXjUNDkaWgsOtdFQZvwVqbPMget18vZsTc2xAReY5W
JCJT6goYdYWoF/j6IGeMz49Qqgu/Nxdu8pJWRjZUajCIdvkscYoaI043OK0vTNDvxaRctppVreUr
gfwKbF97T87/7W5TOPb1WBi5La6excxB9yPHZLCwmJyouizli+6l3IyjPTCekLFEXJokRqDsKYaY
DocKjsgbkxzTRY/IkTmckpF2kYOYFJtp9H/YvIiqtSj4BAi0nICBtebNb46hfV+DFL89M7/NVPW3
0gQ7PcZO+7PgdbzStugt5TofWVZtkOtF/7wh93k0zTU9cXBrz2mXWKl7M149wFdV1yC/DrlIb4Dw
eMDpPF3tmQrd7abj8RRkbBelRhd3dcwHal1nlwDKUJYDfzU9gGScNvvf022u8r6JHbFYC3qIYTCc
df08Qj5hFSDUcHfZ4aGplpJV4fNCvEQAKhGdsXyXon2fnk0CQ1FA75uHF5cxhEYb2WlHm+UwqZW8
5A54rVNo73cISm9YnDJzEjGeY5CzjvzKYQC4rYGVG4fChfG39PrY+lf9+coUUkVH050PaJMPV97e
AB21zKXaa6sfg6d8TkBtj31lwo9OoCzsmECKB6azgxyrZsVIP/s/zHHy5WC20K9gcmMkZfgnt5Kj
ukn91KZkSbc5p/ZPrNcelf8whVGOvd+rNfLfbF4lXsqG/uuVbu8QsyJ0lHucBhNAamjjKy1UDX6z
taVAmFgVrqiZ3f+jXHHEFMEgRzyfQNWXoGK914mQB0VcNSPwBjcYfOmETQTclbTSIXcCThRfuk8u
ZIuXuJroEAlFPOt4CRGzG651xOmXD2RmzFnJYQHKVSKuYHOMzrsIBmzUUNo6odYtG49ppLrCKe2H
rGgMVcc2v9z5DKl6QnxMqquuWWScUaqCfBIxYr93enIbmwcLZD5mpHMLft2PYBxWP272S0LOjhfm
IgTXx1J/Jpiz4k2A9MId675qqR4S9mI5TxSPu+67x5jiudYD2l55kD/qjrgust2mNjeV1417A8/Y
zYFzYQvudCXazgIrZcaW2zWisLL9PuJib+fqPSP5uDjfXLJ92iaVoNPBF395e1k3SPxhPbkKC7dx
TgaapfBOrb3as5YFtXfWCwpvCRTmXMcfZbb/wItuBrRTolI+7PM6LdRfoqA1wX4xoZepdci+51su
NTfG/lrFQeJ0cIJQfunyYMw1fY7PL4pb5TWKdfmuwQyVvH+Ppi7dHWba4HF1z46U1L/sHe18jda/
8u62/B3xTGWKk3PgL4+/SGgzWn58wkeEYvMUqoiWlmnRNgv8h1QRtHkSb5VTphBqedr7JB8n0Tyd
gfpUcDLNdGKUR8HvBXCq3kiVlMQ2jtCjQ4ZT6foxagJx0F/abwjG7lBtxaAoJJgc7nxhJqPq6mxo
e2/A2V94iLPxS1quXo98vCLekMa5pX7t2ch5YhNW+LIqTSh2r7s7ACZrSIXVuLQvzC/pWPkUoGEa
hTRVzbMaa6GqhiKz8KLMApcGZ+AYxvOSbY7IYaGuGV4wU8ruCdcDBg3VyJeI/GZSNqGEUViHOBmD
YB2Ss3a1TEzBs0VI3hehXL0S0/SHBQh0rsUh1icGT/OTGBg9tAYSZJUzWFMQMvHTVkABzMxetdz1
RrBrGuhZTZHXpopZxxPHe9XDmPokLkBViTQv6tKVM5wCW/D+2a0oXtvnJyZUz6zKXaIXMNxVuEei
EtLp6P1oZWkDMYb9DtmlG2PVz4wh8b/5dlelRQA09W8d16ccSePDPKojx0aopHeK8ZPSIQ2obbLR
AiGY3ydBJBh96wlnlE6G8TzqiHaIrWM9i6C0CgWmzlPhhCvJWA83W70IL8eATSwmTvpITlAwYt7y
Y4zgLRsk2/Pl8ecbLv5fPkToSlRE2OTtvF0FigM/M7ARf0Mm9mkLU27nuOwDPOduwVg3WgLiHwGi
7BBKAYiNGGgfC4ji/N10L88tvD9F3Ca/lZ+wo4xGAbVghv3Km7/34GXy6yPej1Bss/boXeib1/Ik
iV7hKhKTKE3mkzPaM3Fi4UXbMx8/Idyru87ft1Nqx5d7OAUacopXUkuIuZ3gpAzP0t8zxZk+9LTX
tXz0EFnkpm99+hpT6yyzjbYpzm9grcMnEso5vLx0Dk4M3VAz/SFRW8R6+q8QdulDkKX7PrpWH2yz
1SSn7XHLWsIfgLionezfqdCkb+Sh2MCcr/+NNe3p9LOBGBFeD4NsTA5lJb0lxogXI9TsQraCFoI/
5AqhbtkvngAwXiJGxN5Mo45ldSpKSqKLivV5jAYYBx2cd1FbVDyvawFBQ8AP+LEhUip95xmS8RPJ
oMQepfn4q0E7v+DDPybkjtPSEelDN80tOyb7aluyloqxqzJiXNfQa42K7gTHKTsqfAFJrQQidva7
RWz28lChCAJL/1RAGPdKEn+BaOalN6Xj1gLVgLRtgdIxRnG/wt9fQV057hGClQYe6xbiZOmQehPs
YIhLoh1x6pNEDRGpd6xXx969GuJjtLr7iGxtvNDncy5md9Lxmo+EdCdaFKWKQnArE2Tc/Ih79H5d
yaMHkN2Ktqzt6BW18MO3Uuxo3hUKdqyJUn3xDStlFTfplBJyGk2jzMPRgKbH/bgodAtyVZxe1Y3K
O7OWYkrO/uRlO9dvwczyd30Mi+OJJzCbXnGDXEqaieN/Iomojpkownzz42gaH3vszeygDhI4XcTr
Dsf70yQHiiOLkCwdMmFyMzzGqljIU/XiNkTrv8CBQduD0Hb0yaLT2E9GU2iYKn4sdqxroAoVI4AF
ONTrQWVVlK1+jLJaAA4ZAxcgydoLcY796+XNCyn+BkSarVx4+6sZRNWQiaRGo5KJQsqNw2VCWc+F
wdarC9bDOrU9JJOWwu1ksJ1YhTuZBAAiYOahFIehZOxhZJiTfJCLzmysnA/KsSeTFf1Pj1n0kBbS
qvhxUQ37BQbDLv85etxnNAAinzI6k1i8kyAKX0nQSY3+v6ML/3n/Ncqg0sBzaPZr0eCZt+lO3hSJ
FNsXyWWmdL7BsVb8tbdvl+QF0arAHr1BBY5nUe8fKgfwbl5Isqm1M4QiT46HUJS0YtT44YyXrU7L
DbJ0hOBCnSvzfqRqpn67zqUXx+vSlHB2Ru+WepB7iKgaJkQ0aBu8ykFcy17zuFOAr9R/yfZvgKUN
oc+8EcPZnhMMVWzzjMbgY++5ETcZt77HApX04mvtHPSLjoRppFqqxms4Q9OOd5Sn60h/ciKDER85
CP3xKdXlpEy5Ogh1GQG+ZVjmSfupsGpM3bw59uq+PiNHuKGI64MQ+pTbsJXfcFPdDCgf0zalY749
hwBTkiCOVw+BSUimScXHGKHQDz7G/o4YrG8N+i0MHa2Pdtjm8wsaajFKs/+qLdiOGnpEW3S6qvwL
R1iYLeHrNw4vhQEdvz5VyQQhy1/YBiNn2FF2zdpwh3yhRxOmIN4Q0MNwA6//WP6IzM2S20GssCz3
c0mFC0DXfLWk7pGnINKIoAca4t99ALPSKlE5KrP345vlgTsLsHux8RzOMf29hI5ujUzbbZeKUHG5
04YhT6ANw4DW/k0Ov+370GVC++Ktf7oqsVj+PKScCqO5tx1pZjxa4RLxGYEB1EekO+TykKlXOYp8
j85GERIGQc595yrawK9c4ApfhTmZvItOyhiH48Lcv0EyKdmCSMIY7hp2H/aN+t5Kj6rZxDxHok5K
4+wHyZr+bwu8YCViOiQ3dd1aYecPxEmzRXeedS8G/L/x3Y7Xbny/Xw9ZCrPnM7ilZrdDFN+7x2RD
MUrdLM+3X/AiSfsvLFBwhYedV9aRe0UCt9kzRbfxgq02S1eTBCzsIo8rFZ8ALYpNZsg6voZBLi8h
y858CAl9WwYLa6J5C5D3s6XE4D4jXZohEaA8UexeECnXfYnExr8lwCWCkl9F8cOfFIg6lN8TCuuR
PiFjLzqJ2mIJiqZ89xqjBwgTxVhOKrVUcegSkwRsCPDgp7J0X4sZxjl/e0RpX38EAk/QQWqpSoRG
Q9vf4ay2PG+5AkEc63VUBkussNTLS08x+HsOJ80myn1gxZX4o8nQVBSyFjiFw1CnzmGDnkxSjm8s
d9iD/TgrEa6HqAZmK0ArnYhgpsKm3vF8LbiW2Obh9gwjOlrpPfKMA2Scrl5/+n/20GbiDickXee4
tB1Q6bHFovNNGKtqEwyuFle9AypHEfQ8L8v4RDujbJU4extwhbLZ2nKovk6PFf8oeyGOaaHRF3fw
M1mhJI7CkWuZ/HTzpEFlQ5XB1Q1Hshv4J0m7pImI3GsPFJV/HPKAo+BDSBmg2buDqdoaqo7JKXBf
IvqgMTI41dlVaArDCjgX+TtoIWOM1KsnwcG2hRpRtxXL8jJQ4hx0uY4ZE+qmwquO9bKP851rsgAC
oeRsY2rW1Xql0Dg5KEgyJoGPprUbGwWZ1RV7T6LXRP8WmmbKWxM+AjFPTNvfVFjyZ3sPqJtv+1V+
srns6269HpdyxmkBbM86G47E4/YOXWdxD0qCx9x6wzuPd2XT7vgfukNsDYt7s19jK4Ql+qNEzgrd
9ZrYPrmYeC4G6ZI5KEUM82tRtVbSQSL8D05CVjzjPatG0B3eBVSOectu90wiFIBrIA1XqR3FRzdZ
30R7lu8xWtvD4rq9im6TEQylZKDEOV4ZbM/t8yDyAoHnTrP+n4yfBoAejdt6qwN/yxZkL0cwXZsL
ZaPFY5VjkKNe/0qPk5+m9FZQuVTlJHRudFuSvoScHy9N8efYsIBrtu958jAHDqHXcJ+AL2Bths6X
nrf1iLIub4lVrvEhHdlNmd2SQ3/Z65PaS85OYoRYOB9da5jbKlHXe2V3LhPlWuK6M9aoR1jwAXpU
8jMwOQNcJ2mWhrJiAJE5rMYlfqmVrXhZooUwxJUYYm3EzhY38DYkPWr5w5uZLIFbyhYfmAE4PcV+
2ha/ytqzIerbsjkpRWrcEQG6sYEqdFMnDbibMT9BSw3ZV9TO9o9be9cZ5arB+VRPp2c5eN8O5Ev7
PCMFuf74ySYG/1lGur5wieA20ikk9YgDol4wYkUPvJzcd7dTzdF6A9jruIakjlhsA6T0CA/oKSkf
3WwQkNqiXIfnxveUki8Uhf0XSGdw2aSp7Adks5Rw0/8ok76xoZy7H0C1HjwvwNhkRoev1xNlJR8f
C8ymJfOEU/UvJtaX9okkVMDlg7r8NLelqm08lzBulR/bTJ8m+U0eAIeWYBwgz5OxHJcI4h5hi310
OktM6FyvbRs9YIqMqaFgiXEJMz0cJMF5K4aP3reWsAcAldc62RYQD+Jdr6LwNY+McG6LBz7aIMw7
fxW4BwhaoEfZCYk1l/6Xg2N2AhDBDgZ65sHnoMRE/VhOYo+XbDfax0SCJ4mpmuh01xWAv5dQPwu0
CO8NFInIc8Hjujm6pBok/fqBtBlSUHBiygAVv804jQ6i58XxjDPCplBSAkEJFRyHXBEGo46Fum5r
X780HezCpFPxsJ4K7XDz0BKHpeIv8uIbUMsqCajcSprUu4Myq3NJsTqp9UkXjChyOHdDpWsbwHMz
hin0DSJhi7KQqL85IEf8cA1DoGx4ze+5XrsAm4a53sfDAYVFFP73tx8p/iPwgbLHRwEVi6+7FStk
TD5OZkmSoCc+ugDZk8GRjNVcEVNoPXmcBZBewnIarsA3H4Dw90/JvtRbGHTpvlVefK+bT+oTT46Y
C/0EWPn99EOyskjlTJsTyAk14lsG0D1l1hMVeOpB1mfu1ol4Un7McJczlrpu9XGKyETySv+DrOsj
fb9tH4p6WHj6q4bDfYgmiDXZnFn61s39Qasg3fGi/sYwrJiCnPl1GPfFYlPTVknx3sJqIYU164mc
Bi9V1YJKCpqzLv9qJlEO7MCTV8NA5iHHluMMKmobobIXA/iHfun0XdhG7eN21ufMeZSdJM4OvceY
RDIeEDJnUKkkoqL3IHH0ywQj/CzkI40/ePezC8BsiYQbsgpzn5fX5kn0KV5ScLDCNxLPeCrAd6p3
e2A1JdIH+GhNZ6AfArCsAp7F4qgM0j6AtSip/etjbrQGn+wUyQr3PjWHGKfIdbO0GVPi29667X5e
l6Z0eE9Bi8JASDF3K4NXYKKNSL3vRt9F/Z42XQ8Brkkjx4Zqc4U3YAkYgunPk2yB9vR7U7s8E4k2
7r3FVFWvwWJfgN35WXE7kLil+dQdEKKmv5C35+dJHewkTNEWM93FlZIsXT3xqxwIdgVjMTIQtQFw
jeMUzWWrNaoxrr1L5Lrsv2RffajdMTs/dG54IhN2lkckl27oviwo1bAKlTo9ZiCrYOylipnj/jCI
TItSy5A7D12xUF1Xpe3c+nbwCoO8xEXU4SotaCeujXpoZ4SXoKBsWFxl/ElRapfX2h9+ievSxaBZ
gs0nklNABjcfQckyQv8UsH/ZrwAdXnlGq90+at2UCIt/xmpPk8ds2mnfy99aITF6/ajWwVvrjTcD
CzJh+jlWdG3n90ZCGC1UQyY9IHiMWpI46LO9EPSCOoSJ+dkRkWzk55W6u7HnJUUGjKVub4Yi70jh
T29vyskTEK6IXmLu4N+o10mp+eVu76BCQwXjwAI/rJKdDjpZKNjjBgUWmGkGUZzq85jKsXXyTH5M
JMlUEh7aXdO7FXBuNYA9gPIopgU64i7EM1z/LCqKTh5+3CBLEjJuzKcjQJCdVOoo2fT4f9+cTKSA
88XLRu6bf9948raoONtdhwXcetM4lh0ZHVOnV2kVndQ769rMygpJ/ucbOAONDXgrz8AgOTw3xt2l
Pd2pjGViDs908KfebsnSyNmYPiXhYTN7gPbYCoGdZ0ypu+dvav/h5GXJY0OCQXYWrIQleN28mVjH
pu12dq5nYw8uMZYtqebaFaNg3pvMCrVR8246QMAbkM/J1ZJLPKUx7fqOGDH4rDJK0ZBN/K5ZM//C
Dw5MQJKW+xo6v/7/a8JIk9BIKuuLbKHK0O9Sj/9ngaVzB/uyUyu3XlkeueQ9xFaD7ycebLo/WjYq
N3pQAUUvxNMqwELqLHhqgOss9sYCndxAXaTD8b8+M7iV6DrIm8btvrn+Bx8dJwmP0Y2e1ePPkClw
48O2A3RlSGGZ4CNLiAaqCDD+aWkKRPEZ8IEWfwHgaIs4F+l3gtaX1bM1qcqVMuQxVQY7k291BHBE
sJGqQzfwHxFYqdL2/oB9WsSspobnlexkGOnjwv3fWEoxUKoFqdQD+RUHEt4mOWtAic68LakYhTFx
t8zFekm1k2CFM89tjrrKxLISr71dfmCpoA+5QxLkY4R0eZz7EtqL9GvRkfvGClOyNW4O22/f3uIo
0lUE5BfQxd2VPIA+R45m40rdQ4OkI+9LQi51hHoIPPmwuDePRORQ7tD5o/515VJVqaxD9kOyXQN9
mXztFNo6qylambhbo9HCwm++jr79a+XCLF6TqmdiTx+PoINbkTQ9zam1rImt72PbyMqXohAy6myM
Ytxzid5WcpbyUcDAoCjpYpwUm2ODmD3PSY+7Brfg0m8Vl2PKa46IYc1meX+JUt1soXDx9N1CHcn5
optcmIpUo3VOwXikh+TwwhpXvJb6FG3cDQGztHmkrrQv+5RcfEgfWWCnWN1VMFsBcS2asdS4ylE+
ZWSmPkL0IFdDkNKzCLt3pol5bclKmW1vMakfydge8xAFQUFj2vThFDML5GhAHAhiT6ZMGEmP03fE
IvmoYW2Br0zm6uFEH5ELc5vWNbwUriAGF6VbPR1xDlmrRgDzpvQQ49Yv6q66tsjryApTTohlrfAF
p9a1UuSAwlaNVWT42Pk5fSCCemmd2T2aIrxtLgAlZguJiWx93OsdX4mtwLWPkenYtInk7szpGqfY
XZUtlnDgkcCTAvFYSLjoEI7nr19lQCOdsUBycR0IpkLApz2XiKRAje6HrdAZFlatM5rxIhpBaB7Z
5cufw+Acfa6asw/PoySK06MbqpzHvcSoSPxDAmC6GvbjXLFmYcElzHip8k0EAzmiiGo6yCuqdlW8
/3RWNyinrbbVDOwdTpv05qIT9XxF+xBakJFq1/YwhjXwu/V/OBtqIXJvTlCC06TWVye3KCBmha1g
u4C0naRlr/OFYXQP6VzBt4O+lVq8/jToQwD31Zv/S5DCdWfTWj4LKFVlsHrGEkr8711lNwLPrKeM
SRuj3a+rNdegzFZvPIT03aXjQ2p/YNW68IapA4ftf0j7lq+SEFINDgEtU/ArRG4Ov36RHy6cTFV8
Gly4fFfTgjD41JzZ5teyTGQkq4yLdNxyG782qYS/ADwtehrBzL0XzRhxGGyjUZT7LUQqbxqRAOCH
fgaGihkX6qyrTN3Gjl4X1KQ87/IiLfaeBX4XtRx9x53FnDKOCd4lMRnoMx7PlpHBxGjZf4dT1ZxE
TkCTTMpyIIDjNUib/ghs3IC6L/wTNhFroUk6mkdC+RjqayuLjeQmbH5jguBXdqnpdP43HUxkWTQL
6bcIbwl9aqjK6/INx3YiVdnPbsryuj+bQ+KJtspt8df8fdsFvltqv2ehRIISw1GDbxTtcO9q3Iyd
kOZvSwQqGvnHHPP6492kSn0W0ZaU6jrukbJpb4zWK4/y59t4UdJYZAIjWXfzRZ7plXtVddMvBNsF
FPcucAkSBv7I6y7NGQgnfCiGll0H54JC0aNM3ftjKW4YWHl/mmZ6TzJ/JEfjcf6NmSqNqOBGGh61
zNI65xIEsE2roAA2Txi2TENlQqQYEBR6JwteBVMGjzgYY44qjfPFTKpASBsxKuy3woA/MOwLxXkc
voIKZAxGrrp6B3QXkuJ4dqXYmWGIE7qBzv3Wp7aXZM0Kbj3KwbjhZWcnz63/q3HHV8V6LIVsy1py
mMvItAifzeloZWvcTaySzbsyPZ2HYYr4mhV+ftOgmjv2HJH0uSXJ0b2RF1H+7lwGGsHYaBh+cCr6
vQBe5clg6gn7cPEOKsjworOZOW8OJpGEA6c3PhRxB02Yq3uHUtSVdfjsVLCqZv6B8PUZaYuCmBhD
TBMgWTL03E///BlwiwEXjxufqNe7Behk3AS2nG3rc439B3i8u6tpRFifeIY8MjRNn4Quq+rvPkxM
KKAe/fhNiaCMhoGI17WMK9Aq0BE9XGUTab3gbotbzLj+nZCqF8z5P+zhpqm0zL0ZhbNQY3nkDk6n
HlKh0a3zzRT6QnMcJyX9SPdbbn1n1NkVtbcgVrt6cZ3RX7+AryjOa57kNxsW5HPL7coCEdGqBq+j
zDadNh8qdQSiG+Vy1p/dH3YniUa5DiSIuFYBvVGezUgUJAmIVcN++Hhcq8ahe029C5V6xJ7xaaty
azoqsJWnpptZW2wy0LwZXqIo3dcRNptio0DVfr0lJ0qlB73fwK3e/KYGlTRf3WL2fzWFyYn4TYqa
ExkV3B5iVEWHL+dul8OBC7PeKP9jxS31SWKJsr38aHZUY0zUr7TVUXSKkrZU7dDNRvmfjoqQwuqJ
b9miE88eWnQirg0Anm76732UMhw2SyQN+qtagNodSntzQEwJbr7oXo2z6k+Vzuq2fX5USfD3Qgcy
vC5empoSl+/U1Ow/6i8dGDg8qgYQmt5TplNLnYewbzApVZZW3uSuNazCQ+5osT7OWKFDZfQvXrUp
C13WUw2HzSYg1/8AairometBu1XzdYM6Mp/8rm1jw8+zJdYFMZldqgJpvInsR2plarH9h6qCC3E4
hA180jvYi5+y0qu2sdZpkFSFX21kp8M2i0OPtyGCVHiX0X5XFIl9mWhKnmqud2HHh/RgT+A9Vk2y
r8YW57oP48UByyK7qX99ZlmQ2xaMOxW3OtJZJ1pqrgDnxQe18pDEUi1I3apJ0gVcXIL2s9rj5awQ
5Ne+KR7zeY1TaHTQF/SB1p8S4TdciIgCyB8M37OozlhJd9ELiILAeGxWoId/pg6uWu+2VXXTRExy
7fyBfTPfWVIjIVLYpYVH2i+Z02dF8GB5Q8EBrCSjEXsNauaH4lhBWnLu6iB/D/ej0FAxJfyDfUZm
bHhnlau+LIXjgBSx+uej1+GLWNnqPqzAEodVrRoQfIBsN1FThsl0j8tdOq8g7ezapKEEa96PGs+i
rI9etfGM3cX5b104W1PVca7Pw9TrFF8yHBjxw98PxHGwDSKeIVqCwyB5j6y+GYxGYOHKujp4mYhM
dYUK4BxwzmkfYE1gfS3wj0bXBsNimKNMuSN8gfqlQyHL6PeDKRMNSLI8hGdxFQxhCENlzZdjgf5L
H1f2BdyOhi/663eswN5Fle0TQAkgMLANbvwOpm9T5j65+yLkiha/X/c9BFxZNCRe8EMOYu/AXw8Y
p7w4uQ3kWDuIMj9mNnViLwme5eMFjiGn64lhpoWo4hAyZ3LFFN01nyAICe+vwJ1IsPTln7K6y6CM
ehKHS4gmn/Ym0n4nKKw1hU46EpVaGD+7qGd/PeXlnQ5yp/zHPObM+ey+TMRzPVLlChwuOM6hcujm
1VR94TChpOIskRw84rzdm42mcVExTZ4WJB0YsmGA9cnHwd8l8OSFDfLxhyEH+P6QX2ntjZVzeZRT
A7VV5rIj2ubtFjZOoeC6V03QvJsk7ZFCGfZvHPwjwhKnSV9d4ymI1VXQuX2AHSV9Lm4GYZVjdlmS
DF8IjHb01ZumUzRXtbTPwZBoBu/oSaxCXLUqf/PMpinh6dCF1EOiPfLxz3DHliojN++Lv7YgO5uZ
fnPC/4PMKxc+C6LwTC6LctoMOBDTY3C1Uvz1Vn4u4OQy4cWmfgWm/lg1P/R9lfVU6V6v6bn+GnjF
/kvBf4nquOvi1X8FFWrrmcnwrf7FPn4yKArphruWLeQG4NGMqOv1G4igMv3Lz/c2zqcXheBcCU86
Y99mK/8PjOutCyliIrTeUzEnQHp7doCCI309jIDmhYFSNfxnxB7tCGacl73XUpINaAkBBo3rWOP5
6L/QKyEDv5OXHLeT5yFTMEGARRZf67ay5lNN3+02a5HZ+QGeUZnhNmqwxN9orA++YSsIot1fe6NT
zilPTGnNeUN/F4US/+oJxO5bhfexltZv37qrbXfbfluFXHhmT6mDbD7wxwXCYVtxdUTHd/DTtH0O
soaaO3iUrqXh2JuQrNpbmjfY/IWyfQ4cpzWWHRok0F6cVIYPeHIceg7feA0NPvGWSz66Z/F21vf8
72nmi7FKJvZReiBUXQUDdU/ezEXaDQgKqs5RgzVa/r42/qBiOae+S9S8uMZxD2WANgZGJQPDjtxE
RvHDkFgYGPK9Dn8c8GU7QaWdKIxYLRqY2CX+Gf2Qn1fH76wk3vPTw3JX7103rIolfHHQq6lvc+yf
a7v9+sMzZlPZWcLmwR9SUcHVsG81w1fjgiaRr+i0qFMhcCV/JEwOZ7Fk+LPvGGeV1BhPLs/tV3Qo
Nh/0M8d4HYX+Np91mMZwS0MO1g/JD7dJqKuAMYX29lpwiCGzhG626BZrNwNAR6gxyUjqHCPIYE7r
v7adgvlGmfS4O9KRL0oritdZMqThPl3fXBgUOVT03tfDRA2foQzRfVpzdKc/0LxqRNntpYzx0OcM
Ypgs9Is0B57qqwMbQyu/bWqCf0A2VBVujK8V9O0evuSt3/kwSxvYP7l75nTm+epzyMYeqGFMiC+F
DP+rI1Bw2M7WRNz1TPRa5ckuUPrR0uZSqlcjO+LYABdmczV+b98g1i5pk2Kvcy+zyC0tNuGooRnF
gdELD0nKZDFOBCbFFBMeqBLPWIWznsSKNpATKkeX7TXz5czt7MyilJNbbGmmWvfve8wR0MyJHW3P
6rSvsWtc2GtuEoAZsSa1NIWcJkFCqHW2pXQn2RWCprWRyvXprY70UUGz+/pXZjKiQDJaQ52bUXs4
SycG+MTkC8grHx5Ydoy0NFqFTgYV/mV0x+cFswiHmX2VVd/ivcgUd/zEUBPACmeZrAzo/CC8ylvb
Xf7yBMF2C9pR8WcycA3PsJuIPpRWATsXiTTf4WfUdeCxUBSVdcj+bmAZAukTOd1++QDi/i6kU5Nn
vHtPMQodbKMSoLM4NQOX+p2ALhq49hJxjKPuObljCNWECxD3i57YHrMPQjKeW9Jyb8bVWFBnCMLt
GHjBa9CWG/Wcu7xQPKtVoF+YFz42jfE8tBKlBPhWjtglqRKlRSX+QnJ+2I++p8ajAWCxhILg4Id2
ANn8q2Rt/l507IuZEPqJS/78WUyct9Q+R69UAJSx1gyhmU+fvzHeoptgz6BrIsqhMF9qpeVT2Buo
+p54AXJ4Z6XUI16GDQZlPyI9xvrJzQPUEljRnHk/MCkYT8Xp5jGtiXZAjK9dEyTx2Ve8sSO4Kbv4
FmWTVFKZkxEmBJISa3svMbcqBa7/BxFhxK/n+/RjYZTVqIad7oS6aiXPSyaNL5ZruKtHMK+OpHb1
1D7V66IjFDVXvMmLeazvnLb+97t3YdHGPSh+dWQCezODGxecGtWRfljX3OVgR+mc0PDiHFcO/6vC
y/cidMUcAYLIgDAX/qNqzf/bHJueGzMtsGUmaoDd/uInLjFKBwfWlXJioWEO5VLKtEnbNMAxaXEt
JPx8UeJiTOKWrqx1XqtvESBrLQaXpJR1+FUyZ/WCtmSkfKbmNj1DyOdM7J0LD/Pf5WZx3eDPCiK8
oCwD1wxjrZLg3NwvnMjBYolgFji/0pl38U6ppx6d4CzXJnyzvYwFd5JtOaHu8oXtOuTip1klcIdJ
3vm78ZUMAhn4SbFNAWls1/JYpL7CvoGiJqYZYclqnXBuDqYHrFaOLD8zO9wTrkx1B5Ne0cb0MOQR
HVpMab/Qx0t8AleCn/XInmMDnm842gZVsbci0fV7YH20yqKrDezEmt4HZemtb2dmHXaTIpgBCn+h
czZF3vhn8xL17LaegFeWycZo0IvHC8hlhGzH7JZRHYOWpkRhAo4xCNzZChkaKVr+kDCI3hM5lhbj
ShsRXhFILxFLIqzfaXMLaY9er9D/2XJELmU+YIEem4IDaFp8+1o+ATlZDU8p4MvqJ6Ywc3NVsUxt
ngKqL0WLktv3/vSS0A1G8K5LOHmyEencmcPwUH+/MGx202tSeUhZdxTMWlaAlFC3r/rFQeT4ZGVb
KJrWyv+RHcBcxiz4IpYCbtxlqM084yQBQzK97BEYbPlRBY9hCkVABlXeoWK+qfK+obq3Qi8IgC9z
u7jJW0YuDB+ozMG7H4jsCCltIxwYIgBjujXNbQK6iGe/qFpZK4y5XgrPtNLjnxpgngvxK+a5a01+
5Oddf/MVkbJ5S5x2WCT6X11E7099/++sCTUhWFlGamHbHlmhmYrtu/to5l2Ez7Dosru81Eqob9qt
zQGcF/iGSw4Vm8Jde9yeb1IuksWXIdMstSt9NaXGhRGvqlQKEXt0LNqzY3qN4a8bw9Rmb3inYmXW
YhX68QMjH0E/jQYP5CiR9hTu2sHpWjUlGXgVefRIX9RuKmGSARY9oanBJRCnNgVPM3uaXU7Ahsd+
3qb3U9CxMmqXWiDlYMl+hXv6oSr4R68BvY4W3CDjCRcQE/lqhb8Wt6My/qj9qqCzohENLsHEkBfu
8CBOb8jUJ+bc2co+021OZX7THZylU4dVbB/vEN6SzAfE6xH2rNpIbO0b8Gtgegb1+0PucFTNkSrp
nYVlQEa08ic8gCiQ+Yodl+hnj41GIS4Yn7ccOH2dfdetY0Am315bnbc+9JcId3cF6NvCxEIJ4dJb
RqbDkriwrSzMGkr+6XERCgGbWvB6QvxKj0ljTN6IliMXefQ7u66ioTe3cj7GWSoOkB/NgfvS/MTT
RttZN1f5fVFvIBUchKIppREM6qLbpa+bRWOE1Vgb0YsvM5N9hKfZ2rn/0tj/e2fr1cSYOZiOerwB
kXuh1aWWI4taMhEPuvrKJkVABvO0EjLUPyLk/sOHFhTUCbK/MB0lZbYzYyglvtPBJujxIpvucyIH
UuhL6Qo/tkgeBIFcqAcr79yRbGHc0ejCmgSZhT6HH33qK0uExpGA/BHTYEzpZIBuNIT/NmGkHHHi
ldCwzwMyrf40a9N91us3cBNaNVnU7X2BK9JqoLhNEFmCI2mG+XpB8lxN0RZPc0JUG0ZvFn9ho6pz
efCEpPXOKOAO3BICqkdgIZXQba2w+UeBik9t3u/mwCpxB8pj0K2Hgn/XzLStLXcBGVzREq9L7AYI
Ks69aqsA7tM+T+/owluTfzKUDwYw5753uD8o1ozZFzX6swO4uz58ErKQMXECKBM6088MqVJSrELD
SiGNtNOZjy0on0UjLmhTPVxbH3wuIsMXvP+F6+nX+v9+m96twIgMVTMv4TNPiYg4gD0g9IdRU5WI
5rPgo/8QiswmwOw4WJRNJBPM8L8uiUwG63V3ZQolEUxjXOsX7tg6NhK1rM9atyM20Dj+MrNG7OIo
dfH+QCsMuNjnFxhbfIo9OxuSpZBu6cFqR/q4Zv1RY0ccXB9Bom1OA1Z2QfmMECzoSNyNz9KSpkq0
qtW+VmVD7/uHscaKfzxLADIHpSX3QiBjZim2kRXGrpeseDlK1ulqm0kMrPSbrhwvgNOwyteDpmW3
Bxg6Vtq4Kiz+dEUYEimpMTxwUCcuKp0fyZ7yqdCHODI+H7al+u0G9G6Elil51V+5JUAiJN4hCm2D
0/IzPFc9Rkf7TtlIDHedaF/WD761ORs6SSuVpTqFbbDDjBNdiEe9KZdohXXLje54nQKzxedRhc2E
s1WW1iPdOt5UkSn5nB4A8hFYfdpDeBWeq+NR+fCQDof9pjMJA89IJbQ9QGHpnNxEJ4vjio7DSDNR
lD/Gsqi+TIxLXEWCEzoReYbAGrYyZYxEaGqZN9JsuKFgswEvZ/811qmE1MDNfATEsvSKborED9V/
C7zuc/iaW4z4i7Hdht5YB3ZsTg4uSiFybnFYbWaAEizQh8hdyPH4UsXUbobmHkV36PBoG9AGpuo0
eZglmCeJ/h0EcXNMweqqEf5iCIe436JaBxhSvctxLdsgCK1X3DDweZwMTQPTfFQ0idjcLtZbGk0B
C2vCTLcrhHchU+zdt6tR9ir/aHkpdWUTO9zYN9kd2JcX83nvrlPH4hsnO0NgenF/E+TY35kMr5Rb
GpkueNZxmLX3lCqyfgMR4KllT/qQatqdNiYMAckPJI3ztXn/SHVvBshZpYZld00Dbb3cHcgoY8Qz
v/pzQYZiho81/Pt9w/a2orSsrE/QUmXdOlWaoyFhi58nRs9K7KUnmJo6/klFvuonjRvAbPKd5DpZ
WIzmyEc2B8KqUS+KVgZ/O5NQaMnPFfTlIgpFEzu7uJTQ4uSpX0Xv7wYbqDUZ0eMZ5cwdCKEjnr70
GmHzsspvtCsWbGSjCl3Ny7U15b2DlpSYRE0OnZfhP9tqlRmnVBE+Nawgs4JEzgdf4Pa1oYVuR8x2
O3uPWMduJAip3nJvyJOqSQvIyhAANVtl84PnBhPc3RBp5clcGw0VPqGdLozwWKQi5A8WoysYzr/J
Jzp56kj57eLla3e9rHbR6kq9NsGnF/h+BsukRFrOp9wDS41OoFY/oxHFCw7BNqtHDQGGsccNJ9OR
1n8L/H5/8J2dCKTfnGczDPzrqn35S6jFnjfBWzia+AMXn4a0Y0G5Oawk41cbw6IEpqJKRldXKhSB
iFWc6ovqX8fQYvhco87klm7osHux4afRLtuAt06nE+LWqYQ9TWgCouQtrmDOm0WlWYs8C8p2RtKa
+4IsEjy+Hs9jpRKliUnYjpJW53srrg5Hxrsx+LPI8k4/CkGO46qY/hUfucdWVdEznvrfLh9aRYjV
K0N9VObVlG1U+cdLsyNtKoLGvQSZ2sEMExFmxTxO++tR544cw1VcSCNJOg5drNMAYsomomm0oEB7
HCVBg3X7JPsuwMzEUBBngsbNn4HCC2X1B6wnkuSfJPK6DZQRocz+3gqV6y+hjT7qLpaMS9/EHb7n
z9w4wVPZX+Vup6D4/6wMMTCubJ7FnGJcSEQ98psZ2A1qjG0dV+sKGgc7qjVukfap2QNfVWmT1uLo
KA3nfS+BFczs0vC4U3LqM8QkOrOl0eVwFrQa3QPhmk5bvPr8s0jFIoxNi0pRrPKPvDmfBYdC6jF6
gldj8h6LGcCdFUyyVqSoMMPInOuL5Y+R4tlmIrkX0e1eEuKWSAYy6Vqtk9LL1pMTVWR09/2Wz0kg
FIv5AG2S6CDKGjsRYnY8yy3DisauvuFTvQvG7Tad35pMrPnpSDMlSWg1aaro8UI991ev+IuKQYxr
SP9yYNOXflogUotnGtLL3+waLGuqzsL4L4GjNrsgu5sP1pf/6hfBem8w1wDOhlUFUWxzr93iRPf1
rY4jmrX3705yPS7U3qNcletxgQQvV2RMitgO5M0OtSIsCOVJm7RTJvTy7gu5K4rugRAcicgprYb/
4rO7d3LbBK8iN8c6ySvSQ7WcmmBxYX95kSZSAwLECzfZqcy4tqCNxtsEjzEqOL5eXOSfbAUGn55l
lY5cHUQBHtBWz1wd0NG3JoL8b0OxEaFXHxtXsUko5WITkPIbEUo4ZSjiLB+MWiHTq7knh+U4ekOS
msmIhZsaJBfHzBRPYJQwvVLhe5mnnAbQxfQo81aCKIK0KJj4qEvMknTAETS1/K8mhxY6Trhg8hwx
GjTf9gPyHKzsTznI36FcCmBmdBDg5UKeaAlvaXlBpvhJZ8lK7kZ6eKi2pnEjbUNMlMAS+iP2QzqW
wXMcSQ9UAE3NVVkyW+e+xMr91O1VdHsJFClErruBPl4JNmJ+wPJsii/yV2kXcW6QBNzqNzHSQK2M
Q+mpwxnEwXrFKlx6Thmb36Y4AG/BodjXg6SJqZqsE0s34U13DwFBFjPPJg0RAa8OvgwZ1opEohdb
lsPnLkTH9Nb5ahtm5M5f8CbaXxgeXKGAih8CyUbp6HVnJgVT2tZBNs8b3GoPxLBJ6gvxHSIisX28
mCcv2uOwTtY7GnAoDXK+sVJqGqUHAgHoPKLigBkWhkbeQHls6FkQh+ObJUoHhoSgKFWk8aVAhfh+
ec4GnR0eTfcmXyu4qDI9RmzM04YPHQc+lu9WCterUcntGevd5oYPy4rwoLwarcvbNjhYZp4c4A1a
k7aQ7HLiJ8A3YQO1BITtNQ04AzTq32LfpdT3+bVFdFD+S5jI6rbGST7ykXBSK4S6X62pvPnMuXJ5
BWXfxfpqz7+vp6VYzS09NtjDE8mwvxhHutYUL+gDZfHl7YQoubgx4xwQxfN3bpnCkuqd5DWbZRqh
cZBkSOiw+/X70z/2l1lMLY7D9BEvP0vNUvP47TsKrC5vXEnH5urYlRZyiQQ+e0gZQ0Z4j33yRsdR
XrAMTBcayEoSzMNbAbMvilRDtQl++TxubZQaBzIu9wU6DFIkPVLUV9OocaCODrW6ER/gRWMoL+3l
uNzsda3RcUUO/KiuE3VHnqfWr/fWD4nAWY8UG4Q0hRQOP9ADcK+hwU7/ZgEkffDv+IX2vmS5InnV
Xdfxv5T48qxztyf21xQGcmqriXtsPEAdT+87Wmjc1GZ8CpkuzuP+iupSWd8me3eyaeMUwxdxc8N+
sk5744I7fUDsoGyaXOjPZGxowizwBHGriDuemPvxi1/Q33b4nt+hI36XEDolyirs50YRTWFyIEtb
9ARqWMtvQ7kKhU/B0cpZrcGxnC/8kLJ85y+WMAD98Z26pPNgyII834bFlAJG3u2r5Ha6FOcGxe2W
WJje+b8d0So0E0YtXyZbIk5AYmYPnFoLu6TTVNg2P+1koGT3g+KUhtdunD2U2Q1/QUVcJJn9aCR9
7WwQ3ffp6fWBV8NAnWBg+WBSO1GkVrSHD/88Y1mv0YL3KWy2jd60QtyLgouLUXg+o4Z0obUxqRqN
uRGinOOXrAFwjV5nKpYJ+9GIb6/ZcfswQJ3NOBhZ0w/sJTHMc2NSoov1ic80carQXGwU8dF0YrIK
97ZnwdTawKGWq1jyFgPRdENj3ntP+ruvDVNtrWRmCgU67iz/1WGLaq4yh6hgQA/CKcRmNgtULfpd
bC8cFL1s5VAe6WsTKs1HIxxUFIcFImmXNOu+rru/qcGK4JTlNWjpt01XHgjnA1YYIIy7qCTjSlcW
U5FOSZzNpCJz2QA03Z6vB4QI2ep4w9zfaqUfa/4AeAlluFWBLEf0Ajyma6HUEuHHJabBdd7LFw+f
YShjl0eqilOQCtJcqGcFNpwioB1wFeXUcKmLlz04GSBnY6tM6k7NpC9OsCgD1is3wg0g6l+blV19
fEliUzpA1thX2DADyuqqAa/4ueSjhD8ZPGe5jsAWic1gT9vYFsS+628MaIZKRJr9XlahYrKe8gDZ
Ov2rFGeb0djgqO1Zz1rqgvjiQPKAcNgpKxuKoTsVEmMZSA1HCSqeVGoMP5kR5+0uq6Axech1SWI3
U8anAA1UZzoF0gVlwS8Zg5n3V6tja7WgfHSemmKH7/4Ue8PUhXMrTF8MMjz/tnFBa245daS1P9BA
bAWsANNq47P9JinBLbiqj0Ce8+g2rwZu8ijet+UTWZWwiT7LxBhUhOjVQoWFRUK3UpZO/tzyb/Aw
pEnWOTmko7056LkE6o9i8gCyF70usnIwOMWYUH3OcmiVnxZu9vDPeMbqplyfpeREvvAxMm68ho57
XMSbYsufdHqlUT2uL5kxzoyXHyxuT0gqSXDRXDfwgvtIaP6PcqAKV52p5JbW9lla9aeUDawo/cnx
6vqsufgOycmLPBnKeedsAmazI5+s8EEK5lj2jLP7TPzn6C27cmSmNkiMl+iorH7MyViQ7Fm8gQup
7XgPE2d2XJ3lLUQyrzM26uRGvGBwonjYkDlNopW0TVpFLjUitXvuaGaVy0WLRUolSUcwpkNvH6XG
yt8KaDlFGYH/6xkgHJKkbHd/FmtRpVD7ZtwslcWPF5INpaiiVLmbjMZvuLdN7PiXfTNA/vz19IPb
/MoYHyi/ckvc3YASZI0zRJqsaBS+UplS03jVURWApb6nn1bDKvMxh+aF5oRd7hqjxQEnTIFa6vSN
ib13BUaYHWdgScm9pFkRcFQa0trDdll3JLLnbJ+yRKM5h+ExaV+j+fltgQyKMcnnXgfZqgT3/Jz6
6O9NkjjLx71DBJeXFCjRqyHKGmMJZqClmPyUxPFpMvFDPLB2PPwWXlkS4VSsuTI0zrAxKKDYhNIk
yOsfcJPzULou+Xf28Iaz6fpJbB11pZws2ZFmY5x/gsdDqkY9A9/K1x1vKhH3sinM40bvQ/It2D/3
+DSaam90shshnkqMVlBxzG5P7a4Z4agZ3HjjOusXN1q7EqQHjUtwZeawj49ObQEp6R2908GYouzq
c1sg3TbFIZ5Qc1Xp/QY817c1tX1HAJy+QhGRjQP86afjbOMOXpJF28WF2AWHe0Qiv8lCSAx3KOtE
cT61tbeG9RNYAgQjrswM5CBC3Dc1d+4sgek+oDHuaBE8lxqpqrVPgmQWrDD2jEfM6W42C0xRGqlQ
MQ56yGaG/X7I6C1O7gnRMo3r7nA15Hqlbul290B3+y0Nkyro6LLokkeIozaI8axHzQdmkfJhnZK5
rEETx9BCdHWdBFRlyxccioAaSbmcOupBuLPc5Eqc6XVHVnteSBeH7KQn4aF6BSsTCpM/sPNoANOX
ov47jnxHHQZAjM9cpQzmb/KlDsyRQAZNlxuj3ftnhwQkgWJCDxUaziju8rUN0G3EuhDjTAa5w/NQ
7r2smayDpMYrXpj+7uWTDpmLK8YF0XtnhaVin3FIuxEvhRRcUkOyy16f2ul4TWx27MXljzGIHviz
6/Zu3FdDnplI/8I/4Z/XkChJDG0QKBSoGwUGMadvdMq/alCdLdJXYLB4kpq61VGHZq2LSaJcdPfN
WZ/3ThUjLJ0RXD7oEoW4KnJERIe0t15mdNse3349/cRPDk58lJFxT/ucuzCHSM2fkLFRpzcxcWgb
XvXac/FFah3A3K4lFt/IdlyCBZW/pkjRxvdX6CSFqLXrEW0bciZVoKS/xmpNWAKgyLvAQy/V80k/
PxrnE2cT451532S5JIgyT39pWWV5OxSjDWrwlMbZw7vZjvlHakR0AQIAS7f8QXqZohkP8obUD+s8
tvECd6qqXOq1lKVnUnxCfbzJWi844DWwkg+MGKBz8kjVqFOGL3zRRKV4g5UcnByEkP4EgFQBTgfP
ffS1f9bMoj/n8ZtDx+jKNztiElYgOb5o3noAYZc8wjiE9VxuuqLY+mAfLRpWgOFpX3qBVPQFoTza
Afd8/uPgrRTY/jYUn7bu7Wy38WMva/JPAxLGGMhfYs5qLMfXQwA1lP6gb9+enQWPKSPREWwjOUIp
yAaEA4vg/DYexGf9xO9F0B+IrsJAOKPmPnoW8c7feQGSkSrxWHItQPE2dj9C0T4ZfJCovqQqaQ50
83rCuxr2qNDrNN50rWCqgvAEGKSH9Ytn2GT98jjHIzgKyT7O94csuv8gEKuBjAmzrYUY/4Hxowjr
RJ+00kthTc0pV8vTzW1YngxdD5q3bywc/fcntG+vQO4eu4yW93X2VaIqnbav47ceQ2yxM6nZFzX7
D4HBFzRvgLu3nzbajDX4GG9mtVvmS2cGhx9kB6hDWPFsBTiP7QZikfKJyYXYW6jF2mDLgeoTxqre
KqwC5vIEGbW71XkxFbRPigvSwQtuvEXHtP6PTIOWI4Jgei/fpBWX2DQ4lMRctnrZqAMWszxrSLkE
VZzhWpWfOpbF8kZoRTZN5hQ0o1ABr4PYkU5wM1K/y8z9sVBthHEHZgKl+D723R03+fBISlEgWhT1
zN+eO6jJezbKkJcqvLks43PUmn89s95aob7CQZLLvkjAgHS893ouYaZgzKoGICXHhI5bvADIU8rZ
cZp6qfspFRh7rqokrTugSAUy14c0p7N2bgrMJTjnyUGG+JFsTRC0KVP7xvuNVE10JjYzrifC0Dxu
03s8Yi5OnO5LqU+v7q7Anb/1GrKVGGAfSqeNGCn38dwEgFmICh4vMc3KSWGnU2T4BITR9tUe2oJS
Ul5lsWTfG2uDBzEnsGdhC68rje+ArIGAt757/ZHFfQiVfWwkKOjui+6yA8QNjFtBRNxAULRkDtKh
1KsqLD7RdKy4KzpyK0ECPU3jr2HbNDkQNjowfAaTAmYSXkyoOJbG+uKrUkdL4+hxSiihID/WeZJQ
4inyee8nJDSRzZqyFCyT03R65KBkmhx4U7AHpJmSkMNTM9X9M16YfgpsU947eJkxSHbQgAXc6EiF
Zeg8lfamVXdYtnfhuPbPFZD5v/oC8Njw0zjVWXRUzcKCF+dNswp0OSiEWe93ugGrs7mpmSFq3PUQ
00JQPY/yKhPmNstojmdq8mEqxlsnQgaNdjW2BRpB/BnDf4mdF63SL2DN8x3/5LLyvteYFZ626xGC
gdtmEYXR23qQl0932Itc9qz1S6X/amH5R97+8bX9VfWk2d3lEpaAxQWk6Hcjw86lo7i8PrHylNdh
QP9XH7//QCbqY0KZQFq5ZqCYloKQwW6xW9YKznYrVfHAlDpeCLsntQPzEMU5m6AeZK6S86KZEqZr
+ZnSB5o0xO+9lRTT/eJXoS2abFaE/wX0ExjWcMUPiJ2QCLSMgEsA/ioKmy/AoSIE0J7mH7xF8WUu
wwAntylESvI5dmle5UZuprEZpv335dy/3QGWRaORf8UhDikqcLbnRwQ/XjKglNKyqBK6ZgYqyD7x
JJooRlc0wmD6bXHpO9zfzxpQlL3y7zBKOuhhO1E4krwVASO6hgL5xhTCiSoZsPmrWS6Eu5QeOkTG
pvEUZDKUH7OHWeh5KU6bI8W+GWPoR4J7HjOhHAwlsPWo0+2IkGauwo5NPEF4KTnEAJcDW4SMQNKR
ijbANJYOP2s3+eaWXmxIziR3pb+UgSSJ/G6paoW+fpcmdmgeU4AvpUSdCBEXGoeOLYefBxsf386z
H5hJ4u472pZTvJtYuFpm+M1ZGTsfTtDv7czxbxN6EewvC5/SJUeEJhY9KgazSCLjCAaDht18c95c
Zxf58ppiR4lyuUezcfEeHNDEuxDFPnbtscQ/Di7kItrPlJFe1VP3c7HGJsZz2LqfM8GStdgHG6JT
O0WOlKM3THnSGorjc2Q5IRvu29Xkx6Muln0jFdGEHG4FrgYe0ckGWnlBNj51UI9dfcxI3Uj7+our
szTct9PF1wlzmyNpCkPNSj9LOLG8jT69jHkZ63MKRccC+Xe+jWcapCoVvuRpZW8IGg/vraXArITc
Ue0YEhMEk6zsQO2QcVC56UGQPGZDtrZIQBicd6zoW8NxKXdyu99OmcotYM7oVJxXRtB5NNhDAjW9
HwvRiEk6G0Qq1A+MuA3j08bXOT2gHKMnQjaX+lNlrCFkq4McykRBUHeoFJxrNdqmzvHe7VC8PzV+
94nyevwm2haE7l4z7fzJQYwXai55b+yjkuu48cpOEqd81IvJKlm3GTafBYmo5SkdVnIozhw558hf
nf8n7dJraMyHYmHA+/oe1YhWMSZOCamwqh0zv7E+7UfHHRP92hh392yL+iTZjQ6xmMdsCF9/qfr3
ULu1xp34ZRJsi7QpBe9mwEOQBPg6iLj7pPAt5K3/dVu0EM23hWQSTluMNPqHSiI8LLWsL5rwsQdZ
v4Kxz2jMLHI8cRONDFZVyOAkTbGXceJj1I3RDhTX5WTIFnnkKixjy+vi6lYdTRdntAQuW+pgH20t
aPNlvv1xd0fqa18OHoHS7a0JGCtS5PHYfr9KuLGBRiqC/DK6kqEoK4sofhlJDq4A5wPZwdpioqjR
GlpjVl01xR1SOg5UoIbKKr09b7bmAZhGvcWSvSdnNNfw0rXXYnxie5KtVImd0Cup5X0nF71PucdA
CCZYVkQpMBZ8EHVdxmqGrcH0fn2qRTWF00sZW4YN4a48CAJO3IPRVDV7Mgh0hJVaeqt4a+oUgoLX
iff9Dv6jh3IZA2rvrditqjUZg9FFdY4S9NjDBu8KxsOfjg8ps4xWN0ksgMVbDFCiEpCP1Z6y6XkH
bO1+kZH/1Le7R4g+lD1I5VAgg15iInqyJbNZUxhQP4vMxl10c9h+4E04QjhFy11+NGOskLI+xBU5
G9sdULDAJuvvWM2OvjEhYWINW7vSsdyNr5Ers7BWXTwjJo+zSfZROpc6vaX09nAfWxkt2EQhb6zy
swJXQKPbzACoOgo0c6myRPUhssuM5HtTaZ8E2f3VYvOd4BjeZJ84NX9nBv17PHpnfwkSC+tVQH2V
Oy0vtH85iST9bgF5RbfF/Qlw2MMidevqGkukrdr0JN49cvFivIDR1uqcPIRTAtY7kC8BrVQbc7G1
vCLbRL23pcVKCXzQ0fdb2voqlzgcZ5D6PbbcBIvRctn/yZtrP8OxlA+duGFInZRjeIVF4UgnFxMW
IU9xlNJLALDPRPzPnuMghSauArOxNfLmVv0KxFsjz2USwyN2ZRkyQWng414N5xqLGoSohbTFItUZ
1TlgQ52mJZPkL6aH+fIyNylEWmtwb+ss81F2oAI1q7/yyiqjl3mbv/J4WdHniQthyD+MzqgL6mrr
/F8Oy2tdOQB2sTkJjZEZRPHVTfU6FbwmwDaHQ4HeWUlbispIVuYxkVOi8m20nFwNw7d7ThsX7bIL
+QiWNqCzIPxo2OEWcWLtDtz1fK+egGc+RVousDx/x7iltK5iTSOZtEd5IhggsvfKY84qlut8KMeG
0wEUJOX7YQet9wT29UR5u4pazsEzSMSgZmpnTg5sbJgtOUr71US/XGRpfqXHxFx4dgGLLOwseGhE
VAuVKQiYEkxq2/eEHXiWqgfBorA9d+shf/GHs07Uf9/71v96QG+nVSycW3l/3jwj70j88xUViXez
suxBjAmHVSn39Eu/Nn2lYPcURvKxN64afuJBzQLBsFXR/LrsBqnEYqkA0IazjfVrEhtYDSbe9vuX
dvfqVS/J/TS0LUNepZMHolNVw+pd4aHc3zTC0Qf8dMfgqZblKYMGAxIO0VA3bP15zLmuZKnPCx/W
x8IoTo1BZswTOD/xwGdT3pxxJM+UliS1T3MQtS43tOaQwTAeW1bYPzdD3nVtkQEUYZaLk/f6vsS0
Y5JputyErCK9EjWHeNbF1fyn7t0nZ4v0FTzYPegqeDPn9LwXzXK0RUOfVTGGbayNOOl9fHYG4ZO6
0f99PKeoJWDUGq1kIJZD512YPC5ezBW9fxL9x6DQxzx8/VgLJKWFKRDY2CEO6zBRgfrI/uMmuaET
e5w+1Z4er9w9o7PhOKClh+LyZIVyaAq8xG4gPNZEQ9LGAT4WrmZjUeHAHZEwyb+ae+LDtvuKGPiK
q5ZlSYlhEVwM+vTGOw2ZOtkA/MGzwBj4RW3DWPwfq65UdGzP610vF8umA389T44Qivi/dygo5/ho
dXifE5LWOlMrUDmiWYod1WduzjUYVGk1fkelNq5xL6hFATHFz9FohaDkPF3aKc+lqMxBG1/qnkff
OL0K8OHzkDGIB80pR948/Jv4wcJbUp29OfPC4H3I+BrEQTkOCv0Ko8hpA0lncfgzMTRdCdg8jIro
juL7Oybh9Wc31BXZl+PBxcTMsYRM4iNBUkW+0J9OuWycxgpX/u6Hot4kabPersGXCoT/MCEg1BN/
Ez5yor0T07RSbw7lsrpU59Z189trGxgKNszlU107UvGvXx1Vpz/PYtsjNwdl8Dz6OV5DuJeF/HC+
5Uqe86ckTyl+cSgsWro9qWqwy1nFcKI6Xar2ym835jKcEPvrgQw9eTZuQk1/7HxU4dWgzhJkFCQ0
aHxZNh311nnRQAZBnU+LiAU++PwqnFuXKToa2O2lrL/1yfO8xI6lyglK/o6kOdoIplan7ierCGYD
EcgvdD5GMDtkiJc1B6hPrTY2+T05/GB0G7zli+qpnLXSsbI8VdEpkoW0bqbS1C/45rwmnbZTvGMQ
i8PaJ7jFIASfv2bLLunYy+2DcXSlmpNeyD27TPEzrQvAetKIjVrJh1WlsPPS09Y+g8SFZ7XG75nM
+12h/fg8XaPyzqr3Mkjb1iSjSf4vyUoD+Dxbt0Qf4ZIl7g+spFL9taUqaP0nNeYCnIoeFbaOlUfw
Veg6MSQ/aHG3Llgn5qe9vuWjPk4xJeuymtmgi0zldBaVOd2i0zBuf2CUnws2txHsrnHVRxvyEO89
1bBrniGvEiaIoawQbUx5T9+thtgYd/AF/LQ49eHTBMvAvMaqKSMCfdiFlgBsu6zz5vT8IhOFhss4
+Q7OD1e7Hs7p1bSIK9AHGUYvvpTe90Sjz0y/62wiVYF61mBkFiWP8DreFwI/KMl0sSAiveACzA1j
GR6F1eGmb9k3UA6qo50XQYDkeRdSJqJ16DiAf82PlfVCoKyK59ZRLAqIC2BGAMKoizvfhWjm53IQ
2KzUKZxvE65n628iNKkDTKI0pxdTV5hAN6cVgrfxr+F67Ix9qSq2xGjcjSQmdZwUtrdAGIpRv1FP
n7J5DdXORSkc6LCzMIi6lUVBMICTSi7T0RUkLjrq33mV8KAj98Kgy2P7+yJpPdBZ0k73jTb3jxs9
XCY0A6h2HME80sQu6bznm5U2LBow451msukW3wF+jfE60j00ODyBH1gtAxKczILe+IOC2axS3OMB
zA09AD+iFG36hy5ZQtgqYGHS5iEY2F1eTB0KDkHcYWEG++JGb2c8n87E0jBU+A5m5F2WKNdluQ7A
FmVIYBsPxIeH6B2maRsBC6ZDALLCUs8/2/pQaSxWbu0/PpXWBu0kdy+Ieo6yNJd+a+MyN2DaUt4T
2P/QCKCA71935sgwgkk+Kk1KM4Ld6W9hy6Ntc3zN0o9RH65p3dLDuHchgIKGBe0PFK+TcZzeIERF
ID0iakENXQ2lF/UOR87DOEsLz62bc7PQEukurpoIAV+N5bneTsffDSQENY1JU1j0sbCIenvN4Sp4
zyLYrPcHQPjkAVARy7ElQy46Q4QROHHeZ3l/yx1SVOU3wjjBbpegxXZd3ntcDcU+Q4JqDfrHRscx
hwOB7k30TS2a7V/ed/vxHq07gsuQX1MgDBOdjjR7+l6710odgkWTwJFGP1egCYNd9we2FvFsjy9U
lwDJoum31fQseZoA2IQtI758Tr3cgL2wbcZy1BNgkez49aTMl5PNKEhXtJnNwce6Tq+vAN667HOW
c3gr8sJMmpuv9XD9ve6/5R80kXOjt0x7SxJYcgLkCrOW0qXXsNzfw2LanSpvqQPuXMP+UuNhZ597
ZqlLGvUBYoxt/M7ZYmPaA/dhW6vAozeiraDZfHNMgsruEbcEDtC5rd9BumR1y/F+Rle7foQzg2QQ
ex/9G7JZAN+dbPsJa4MduJMZnePCHUpyd2OrsFBmjrJFP/1ujQWxu0FG6vJW+T7LdSNcU3TZM/Hk
nc/+XVb+TOCLFels5fChTDVoyiAreAFQB+z05b7+boWVHLHQa7Z/c5ayr456XMONOFh4K4DPcx/k
Jm/bfXCd/sX4ni9NegZg9qS6pjDz6AF4gH1T+tPDJLZYIZuzuESs6bzEIAoBDo+3KwFbkaZz0/GE
duXBGc9l2Uf0UGWsZ+pIO93PenbNUto0mDcby3CzcvfMQdiTtQaQJExI5m/zPBjKYboL4KxIX4pf
jm9ShnKnUHFkEuBHnNAA35+TvKV4TrcoPbqN+9FcasekOJvyIIhJFM/DsMmzq5BV2tBOrwpxi+bX
6HVMVTb/cQQbpJG2AKP52krD3YDOQ9+opEgSMZ4dRiEGAsA5M10tR/oobrwXy079ubQSuD0gWLsN
fFXMPZH+XcItT7oZ8dbnulyt3+oAkyi3eFloiDWX/9rWXMvlRxYpzxsTpSEfNCdmESRXnUuBt5zy
ObZMOSW9O1TzjcMjelv9/bx96q8/X8sogxpoUhA5JKzpdOOkRqLki6VTjNg9TOOB/FQ3iC0LP0lS
B0bfklb+rXwzgMwTuHV9LdAL9O0wYP87wDVWLBNOdPWuTa+GnBNLh/i0utW9z/f+j39EM6W1au19
9FQ+zld+1/R1I03y9J/hOeOL+RFGJoMUK/uyX6F07suaJaJKfe9QEIh2/0VwwnP+SFFiNb7A60xe
gg6Wo3kzRhRW4FY74xRZUYH8VgYlZZNeZi3SXPn9xV9Wio2znpS2qLrGmG12h67QOBMpWLzWuVeD
1AC4C5GuN7rl3Dk5iqt+iRQ6jjgaOKqGo1xaqMzocV5K0oOeNiugjZHnTf6J+JZIZYCYSDZ+mg9z
dS9bdLtUunldh4N7R3GmJNB5UnyvPKJ8ZXxGo8DwZMEbNioEONh/UtnSXKk+NNqx2YL6BRE2ZPv/
96Oi48m/7WVK3oVmFYZh4EeGutEq+kE0rRo8F24sn3rSMHkU/UZMvhLprkxibfA78vC9B+nZtXut
nC5dAulYgJC4EWhxUeUsMtFasv1zWys29Y//a4WQmSf/80PSGlBTfBM5gMGKiUBxK3z80k3h7M1c
/2tDTO5Yd3nG560Pxk1kFMZ37A1bEqpcvPMEaF40Fmi0bzfdXdt1ATD3bl1sFa5YF0JWwMY2h8tS
cngrfRDOEmo+moiA/bxsNUqZ6VXk2Vd9rqYW6qkrcW791f3gJ5JXIFT2yo+MfMe37FAW9hX7ImhF
sCFE2gE2ikxDJfOQxmPwAHmCvvTdCJNjYReJBQzWzg2vPvo16xmFi1sOQr51tsTxZpcR8OzmQT1y
zJYP2TE+xsYCSYSO7Qs7rKE8sRkWL4YOAKUr74w/2BsNuPKyMpFgMWUQVljgRXMDQoOWzg6vPudD
ze7MgRPocZH4vae4mdQifr39V1OZB45imhRhuczclXptYrmRbgznBsDbEA1/ATocf2/6oasTmdjH
WTDnxVmwpodG1nxnHnpQL7rW5MqBAcW+THWJwqhsw5WNo41bAXea6v3zOaqOlwaDfCGL9+2EawF6
n5jp1NE8nBYHOiHXhN4uzrLiKok9UlIelivmdgcsMpSlVsu8AG1YJE3N6i0RAqoAGTnxoFQ6DjLq
ainqCDWwEz2t9GxokNDjwyI19ckxVLUOABoWE9ZNJTanNzFcddnU/ZKkyc3k80V4NSO2aLRSV1FD
T0L8V+/r6votNoXtCDXT1n3iq355Sal6tv5N8M4EIccpP+U9GyHM4g1jBzixaFDHhlt9lWTABcVA
vW8iMal1K+avpnt6u6P+/r6UJeDfbgtyQlaR47Bq3ilVnHNGNqzJQEDp/Qld9f2fuMfP9Zu1+Uhk
ESCFyOeE6FkJLRJN3Fp9C36usEC1AWZ1kwd4LpscJ7HuLv0xko1KGgaPXBMkpi0hMWuF3E2zNUCh
hqGyRrf212ArUwtpBa+dcmhubP5oWBm4b5pcBHVC5jvmS/6cy/60UXm70nxGlersqQE+U5INF1g6
SoAyfes0I3FD15qxJbaXkPivRc36rgMzOmb3dwNY0pZlRgFRfyEurJYuqYXyfaAvXJcfGmoe2TXt
u595Ujm9DNmTd5bdNTyjmv1bPWLT/5Gkq7ZKquLM8eZBZES+rS/gjnUeHjU4GApAea7pvNyJ488A
uIV962V6FbBZYxu4XyVObwzIRzoTKyZM0W2fi4f1q6e3AEjZaJBYvtWaQ+gO5Rz3FC9zriw7fLam
IiQAIVYwhZ0CGMhYgbzsoPEcPjLCmbR5ObuBz+LUqw+ExViBabtRg68vnS6DotC9lJDhaaWFIRbU
g/x5p5+2dxcLxwel46xummO47nbzbLLfgsgZOFg3UROcXGYvLAcMupVtcseQ53Xa5fZx43wpZUR/
MTLNhlrNnHYvKvHV7U+K3eatHdYq/xNbzH8/XxsTr6Lt8g7iplcMdaRdn8R04BxQ2ce0mhmp8klC
G6Y0TgsQ7xHIWwqHoVI1+qcnBcyC8EcKB+g6C8Q4ObB9F9XRdor4fEc/2RmtmeTqOmBVfRZOqDka
EF6CeoQ6QEI/7X6vXlOEjIpbQ8O1OrKaB8/HS4cui/Gf8Du/6fOBetjiLWOhW5b6F1pXwvdQqRHE
qSe7J1eSTKpEHQr1U1ZHszwey28HkqY4/qoqBJeavwlQwEIVCuzp78sI+B5+o+pdRWyYGjSSNgp1
nUm6Sr3fn6MXkgzV5TE49JlHeEBh4Uou1n0ucILlBiZWcn4ksyV0XTVshrZVvRUGeQ59AY8vZ5lZ
A6JcXp2WfBigxYOfbkZFm7DDtqaH9oixI89ACs+RGcSOOdvmPy0um4X9x2bl80dxwR+KvEw1xzHN
kLg0DLF9Z4yuz31eEPeApwiiJW8LaRNfsyguy+lQI+wdLopkgn+WnoJbwkOUKnCIdUZszhe20aDl
jocQwTW88SWUya6nPj9L7Yfy2EYFEcd2KfzHkQb4ueaJ20UMbsJmtjT59XAFIPMIv2lfFYTAp6S8
yR/0V/S3h4NMD4Buv+fwjgaDEd51VekDMyjp/TKoVlMR85psfKu7snpWXpFXkaxHuRudOBMkDrta
0k80pFKX3iT17ojcOO5LTRztxHAo6KWNUl8OTngRShTM+l8+0nFbPr/0s+L6XWI8aiVW9+WWhoW/
/ywK4LLp+cf53rHJOJT4O1BxAQ0SYRJLzEtTKME6nocl0bx2Iy9CR4buQ6IIcEaqvigYySrPCf6j
BFtZD0yV1460CVCDAGV6CKdJWNJXe1AQhYa2LX/e3LYuUZpAUibqMgDF2pjWYPbNwA95mP6+k5v4
MlUXN3+ZPzKWmbpkE3UB7KwPrNYSeo3XBJMjbiy2emWpIUwGSGWCrzPJdiMtfYaoriGI2b4Wvbyw
K01c9lz5CN/LdCZc75qLRQq+CoiPWMnmBGS6LggL5qkoK15UPQlbpQlWYU1P/yAjhDFi6lo+tkM9
QbINwHDiUagdQFJxlYmsWtNvz96Rz/gpayuTizrRkTmmiPl73i+q6cI3PdmWnA3Ga3Np5aE1GvPc
fPtXi0YDw60rUtUlxpL9nWOcWoEa3fIlX7R0rZP26YZR1RHB+Ngj4K+UEXZdT6ee3QdIDfyViFDV
QPDWj5EPipK7/SYIlOSUoUFasZPPeOFp1UVRXb2ubdDhC029nHElOy9DB4j4XUzsdpz5PoOZdSZf
goZ4pgJPOnT7LiwOL+6r4h9xRiQywu+nticjQQqXim3eNzB2YPpnPhq4LBwADo/DRaTKeeoey6Wo
eokchlf9Ycv2TbDzJxJ3L09KcVxkoqumiqh7KGwZ0/Wc/dofoTIny+pz25R4aq6rubKZXmbICiTE
jnrW50KxNybTKSThQ6BpR9WFqccgfZ7Ik6++KnInmScHcoeAH67IPSgczzw29bUZCJDah4GPxiJc
t+zj4BAE1QP92KlabecmO6Tjbftf/z2T5O8tzkbzitsy4+31oA8FB9uq8LIGa8vKWDzuV0h9w8bS
d+GV9QpdZKyXIyBS593zfBoSKSHMk9bTU/8Djl4mc8caz7I1oLdnBQxRF7vgV70OwEBCFplE/o/B
R7hHE2fLAv7yubcXFjlamb52GkWhKaKtB/Q15Rg8NG9tc4/5yX6/2AjsFVsWaoPO2rPRfyKwktYV
Dl7HfAhoAgZl60dPNojmZtSVZEUZ+EOwhEU5ldykNVdgEmQW4s05Y1GNbQPXaLPsVTde7yBNHaDE
g4QXoRUGrG+Bh8KSgrcasduI3M5ywcTNQgSlT+Nri4iQcHCtVUz44uNlagKlMpV04hbGNCeyYTLw
MPE+CLOam1pvHarFG+xc/JkYeWpMSl0tTGRXGsNCdoWKPJYBFSfp3ewJTzU0CdyH5T0bd4NUiw+w
XB59DdOVqB6hFstYjhC/Abbq+1WxYXxXGclB3QjAzGEOH48sp4mKDBugVvHhK6cMjNZM0cNA4BOQ
I2SDN4mdDdeKjTW9xcq2CmY290GzaRwju7dagAUE4H8HqfxsVPO2er2MqryoRCtHPibrZTN3iZdb
cvZSjRo1dkmDnXRIFIENecxLRSYBLJCdYChs7uceIqnoQqNOMZB5Wo7VhCn7EezS0w6b8XSIcCr0
lWXN7valkVXa56VquoOF5dzkGjCNOCHwNUxK0ZKtxqwtB7gRckMs5YtrOr0BzixdV74cIWQoGU7R
BQ+I9vswpdBc48Y0WaoRI8hbQFbGX1h/qqXF4GjOrpwjIZCNmavL0Mxe9YvikSdybGQBhOPxbkNe
zKKhpbMSz1sB1pnHsR1SPMgs1sfV/LOMymnYFVZ+jCkbCsU0bptbo+6xRbnehDsUsyQLB9HBPOBb
T6SLsjQGRS8guo4zmeNPpRfkiJVrb6JuIY4iarkpeAP5HyJbXhUa5zbZNABcDwZTH/rApdJxSmZQ
ToR07pLZ8cqQxSVurEfqCtkfT4AxGqzOJ/Mbjw78hhe+sYIY5H+HMQo9IUbfNwmMU0CUJC2S7L0I
F6G1vVscdbI2vuneAAyrBSkC+nBDTR2ExTfH7xG+ZSgOaO1Br5vTdnNmGpzXo3kUPpnu1zC+rzjR
Gef+7FZbDPtOxWkXEY4ZiWXfeK5Od4PyYf+kJbbNWvwYxfYdRX17sbnmJrFQQwO90KGJolA44yOk
++5Pq081dTd38x5iQ2qVaLukM8N5CRUYHU1BzO0NjTfwTRA8uxsxu/xPl25lFt7obIjJOXTNueMw
NTHDnXT7XDbOJi3xnvNeRYG4dG2TLllC/Y6O+H91dudlYlqVKNRlbnmkTSrLaLzZW3C+Ja1uEpu1
hWMqX66nfbfib39bYtxId3NEGZCiEGZFg7OZe3PogDk/pVRyAjz/vNYUahlhKrxIbUU32Z1o/H5T
8RGbI9PH7Opgg7ig+C55U29UyBg5vmUMccFX0y7kbfJS6xjD9+x85iuYsQIkFzccq40cjX5P7Hrw
zrHFrrXtPGCHl8QT14VEm/z0v9+Ab4BiUUGHUw8+Ks7f6nZHHDHfw0fy9H0Qa9/OypVlZCfcEyDE
Is49mkbW7bfQv0aRmVOv802DcO/7lV2DiRYsu1HPZQE7V4/Ts1a3W+dKn/4haDrR+h//MMWBJdoB
YrztjaLTR5XHxxT39g3CEDo/ImmYW3nL/Vb6zXevf8BPc6iRJSArvsVklJ8KguU8DTnCyKg+iDxu
7SqOqm71n8L7KUMATajGhzYmHcJEfe5shQjf5CmSC/2WITxKDYPGPNMjLFcnzpdRnbHXAAQD0sMy
KypRgy0V2ydPj1+2I7XIsjHeEG8eQqzfcHvgHZdc2LDlt3zlK95EiSPBZ7iE/ptOo9ZJY0F+Y44v
EC+tPpJZyf6GCVvG6bRhFgK3N2+KlBqiVcRpRviax1ZxTx3L7u3pNqakbOiVoqVGWzABtq5vNbjq
3lzMYRV9lVs+7HtvGLQur/mWk+lrz5ezA5nj5YXtAiGsEE9dXAZ2q/qJvMFoihZt7mfQKbXqfKUh
JePif9VTHbAnRqrN+yfHm2yWF1kGU2513GIy9n8lw9KYTvod/7Fq37VIIbByltaVj06lrPP4B7HC
m4W2JWtNl47+QXByyNHpjxVPs1BxHNoTXeg/zNij0eu1GhjCs4cCJozHuN1DZ7KYA1NHWAHlDJ7M
olMNETyIOxyuGDsgg1/09pcQmWbULfnc9LrVnTHym36n55KyjXZIf+3bF+1w79T9k2RmDxeL/Fqj
ZNmOw3869ppCyEsXLBAZe4YONQ/C5cBvgwEmXoAQesgebk2bzFhojK4Yk+0okmHasD9U9UFoB0hu
w4VrKT/QxkKI0vMVoHkgQXE6Tokr3ZlOne0qrFg4qWPUgEn/FYY5mHKCMV6Ys5AywuDf6iFyaxpV
nWYcLb0HNcNCho0+DgX6CZN93t+j77WX7AHPR21hdYqq3ub/XfL0bqQbsjYNHLlO55NeFwOAhsyD
5C18b3PDZNWdkZSciG6YWweAWQFClo8c3ucVnlfDV+4xuzlqiNfvW7ZWLPQcPqRxaaXZkQwcpoAe
PvXMSGko+wp+w0EsjuJPZ6GHfHz0tcFewa+r854acXVUAWdlWVCQLXl7Wq3nokKq45DcBaQ5SfgN
ujO+4t61SzQXVX8yUWYHEi5pu6iTMVbl7e8yJ4KiTjvnv/1JJap1nNcHPK6wHAYo5sxt3mjJjRcV
fnp5KelymovKo+cV9D73yMy9IncougXq6Vjo7HU9hSA/bYMvPRnC1CT/HCkCoVpYMJ9u4QPwvVJi
vaY+/SiysjujxSnzclDFiBNROgWNQvJCuJ8brv6DeQQUetxbZCe+AHQdStqNcWjkxWszv4mLhxhS
xK/5wLQvw3U+kHZ9azxr7J5rSQAoTWSCShGPEN7JWqm7o1JTH8ixjjJdY2O3u/SOzqgwVddZHO6H
HTxFTI+60v61GJQuN/jgwKY8B7mvBgdMo+ayykjedWjB9wzvbvxfFYWiYCpodt7xDriZOtaEV+b/
tI+H0cSq0wylzDXu5p/S2M0/orwzUVQh44BH6tDlyb8CwclVNgbvwyiMKrSYfgg06vpUAOd4k71Y
Ux7AsqXKkbPL43WVC2G91Z11H3W8GtjRLsoYPxB5Mzw5PaCKTnXwGpikZ4B9Qj4B7tuDAUUgsGcF
ZsX8Xe8Z3E8EIAuLoueVx884OFWUjVXEKDJrKTHpicy+hlEZBFvP01XhHgIJnAp6Fp85TURDa8vL
K6omR95Rn53tol1qd6lQ+geiypLsveA9Xh688o4QVmE/xFL78JUJkUs7OPH++bYdjCk0lq5r71Hn
OiFYyckGwIwyjQUHlL0Qk6qPm2JzMUlaXKsLNvWMmimKbgy80RFspj/1PNMrqq4+DaNktSJ6bqCB
WvTrKQ05kBQtmU3aVY/LHLRDvOHi2IxxzqLO0aqyE3rzpguCXWG8oIJsxBt6nUOg5oLLnLkvO7S+
mSe0YkD6AkRHUybdYPBjeqTcI/mpnPbuf+e02hLp3w3bAw0cCZ5CwY1k+go5yoIWsS48JKSacrcV
HL0R19k0qqHzOYYKhN45riZ/YNZ+SNQnmyJOkS4QTw9v7wKfqChk9GNIkkwCFixvVFl4TALkHxjJ
Cc/wSjVVTYMV2tVhn59et7SnGdDNl1GHKzJtMjvoKUSvtc21IOiHYSgAzhsjdouqc9de9tznVdBe
i5g4BSbb23ubZYU1kRQ/MA2zjddHlBiUHhTtFNDk9Cp6QU5qNQCIHxtuWWn8DiQ/veClUfJxhsKn
Os6phvu2OJ7twR36iezcCnpT9D/aKo2zjHvrjlc2OPCv8RAHg8wZgC6cSGoCcqeufXJ6+EgOiVka
xzMfCQKqgxOizfA1846yXj0xwOHy2w1i932dCDMdAzY9dXuKVGKpwGy8zfUjYkWRVg9m8BiCMmyL
7iGihmho/4gohIZxJ0aZrv8Acpou557UeSAjt9pQNc5CVa/3tqY9clzGfpcO9CTv6/jBgfayv4xy
xO95eOXDSRV1h+8O+Q3qcntnvG/s6aOuKNThJBCi/mGSJ06b/orkhB3O4IWqOWVHbvS4wgA89xCM
QiQetDhR6mleoIJXMo1SlpPWONpxQUkwDE6rzhnlEeuFg2k7q0pNKFgtRgxqyoSEfYK95KdjBaP6
qCW4ftvXrpmzksItj7q0YgpEDQGSn62MmmTvyD7zLGJtH6Qi4fdtZoll98IC7nJXScqoLYPfpv8/
aa4UpN6kM8nXjVV27S+gEbTxO7gFw7cGzRWMKHYug9jPhb1Ol7WYVMAMwYTjApRcuuP1qSJfkn4E
yFo7esJl3YcEW76TJU5bpGvHzE0OMkfoMM/+9ow0t7vzGBamptwKDrS/mKWT0seReecgVOvQeVS3
Tzbv2v+7Otwdlym3oPNuG8kl8MWlHPBA5YiDx4D9aHKYsvmeA9YiONhYB5P2bR7dIMg69KuBgK0a
7xt9cuslQQB/+KEenedFTeteHtJIrzMpSvibAm4OGiZ1faaToYK0r363/fNwT8U9GKYRemCoVzRw
KbDcfLf2cxwQlZJafFFIBS9kIL/gipenxojAx5K0a7LBcI7RBLUlxMJ59WXij274P9ZIi/ewn+zq
R6Nn60MUwl+AtEWjCqa2vKIN3oOvNsu31wQCGhsLs2cSgMZCYYZ6MbKbzCSa9/6Rf+bcUtQQ47xg
H9/zTh/ubthuFo38d65/kCTvr75Mf0YYm0jQr1mPl39kipa9jf5xOu25dpZZ8Hqq+RauHTuk/Z4Y
nZugvCsFN7hWYZj8h97gwAyr1NPiQmkrMTVOC5Q0iHIRbFi7Sz5Yq3gN8Fx3aNsIIeUUCCmTh/up
tU4dH4PFjq6Vx/u44a1ugQ+vExYMDqW6HCgfQxBB17HbssQhXdRmi3c3NaHiSDmAOHgt7HAE9/MN
wEMaFWPrS6Ay5tE+AZ2iSmE7k4g/xpPcYxB+Z/O3LQUNCc1fsS4rl3pLdU9p6uq6sMqXfVelgbEN
0h5W1hbzRbZ/kKEtnh9tKFxtKHuUbhgwpEej3LLSp4aCl0dTXjJAYLmUT3X+gWNftwJ0vjOOthPE
92gQVxYNwigifrqw5fwjHBQwtZ88e4RJuB6W52OmFOXwpjJB9z+lZWup0GWaYRQOobo4aZPONSAF
cxgm9p0aSHgCzYLaQWyS1AGweGca/wY0xQu5EvjVACKtBLT49DI2FStLT9JtlsjfhcwbpmSKDoUC
SE2Zt4IxrVeOLJM+FT193Is/4mg/5ay+Vq/KP7lakR3K9tCOLOYsI3/gFttuuzEvkZUHuJtNTItb
DcVjNpRfIkbJ/QzzXe2928bsLIMbpb+mYLqhXfBhHM48byIZVZmniu7SAhL2A0PL2gKQByNMH/VV
YQmzSOzHSydzHErIz3/9Cdhfa74Tng7NpM7wnZpnI12q8RRChxDpIolEtngPjFBxOYVZtRXlAnb/
hB6WUwExO98tEffWTn4pnhFqtFTIozg/A63stG8rP3RljCxxNUyTRxpoNSiQW8dqPrx5AIscn8yK
3Jn/Oz7ebGQyY/9lQAoQkxWsDAG26bnqHZKsmL8ZGlcpICTv840Rm9S5s89pXkbxNyiFMdQfWCp8
yfIdMfgPB13lWQlhO8khs/OROHHWa7dctvenfm2V65MedDPVwZjKb+E/jAHP/1+leaJZ5pf3iWmU
JDMZSkapW4Jdf4g3EZB4BRICgPwpBfsLD0KuqmrNVWSKe1RoZw29UhrHWAAacYKPGGDTsJ4CA/f4
is6Dt/Sjt+2V2gcMHsJJf+zAQWTkBPgU4PTctXKyPiy9LfJkaC0wHrPIZieRvu9frlJGoZU+L8Qn
zXRZHcGuVoxlz/uXFRIc/oqcrsMcUj+PjNhdM2Wny2JtwZxWevD36FOkCunWPSBwz0TJiJbxzKcz
Mqd6gkR65mWAwyBqFG8fp072fu/RJ1U7drcrtodNgVHcni3Sgtt40Yu5c2TLJtaxTze5Zu6EqZHQ
CaMFHO/OTf1txLAc3GjSvd5dzP1rWYYzX97H002w75kCC7pQJx4DO71H1pHlZpqkRmKZc7snL0RZ
P9zNaOhpyxjhE4flEk2ysg63euN9lXDUhKhn9cRU9S/FQtVzdE22ZyxgmW4/PagWG0vWI/b86eVP
2wUjiBlwQjLJZr7ckHDGNEHztddMTbpwy4XJZL41y4NwQB8ZK2o/edPoAhj4sqH86Nirh8dXwWKS
wg0guKJJKZuxoV1Ua7+i1JN5GPCGoW2nYNZhkrUSnkVcVZtuoxuE6FEsUJsiO8qCOLRPvYVhlhqO
4PpgTBpUGokUcCcHN0gAPAjCIugu+exszuwhm2hcHA6FmVSWMG82aMxncaqs7mFe1dwFtNT45ENI
weBYp13idLKw/ycRwJ4+T34NQxh8ef1prS5b2ipUQ64253d+v/ESnKu9k3QWZc1igd8BSKLrmF66
dPEhNf58Sa+ddltEN+r2IJjX74iZRFjn++Dhtl85L1P5Tvnqb6IvPmsJDOT6jyICuy+h7ce53NI8
IbxSQtqe4IELgz3CUrfkbVCGImh9LIO5jfkWyqngoDtDAdLrDUREUhxME/eJMXnj1vjb6u2KyjqW
Ngv44Qd343h1TcVNFON/LDtSHCIjmRXBlVuSZUp37AEu59f+XZn70pBddxXJtelRbz/nBU9fgJOZ
S+kCMsIUbymjezfIkF0TfYUBq/0E8BR5zvptHYN2+yT6FEX0dgi/Rr8E3luQ4YiSa4B6zPAvT6Ds
z3jD1h8kU/IIwp0jIbExWIUzbYSxds2Nw2/4kBgEkOkKIdbKtuk92V9zDZpEVnxDJNYXmKR8L2Ik
QhDhdhpL1pTIdj1QmLYtDOpbOENXP02rGbOawh5JYV+s8+I+AA+w3x8ga+i76rOP5XhEMtLkYTPT
ycKAOs8mkPlJRimXfzv+Y1LvHILAE0cBsTqB7A8SvZ8aVzzHG7AVPBn0L3IBqKLbDtP2pChsP2J7
B9AEkA3AEjo5arcR2iAJHSvU9ceoDUpQUy8TSkcU//KQUvvPRuCIyxZi5qR0T6GEgQ78c4p5cA/W
6z84xkX4TwdEqiDvMjw6WEJCpH4Z2bAPWLCW9rs0FR2CtIDFa8prjpB44YX0dSUvbjjX31IrKPYz
KLtZdmVk3Ab6+ZaakPOJcp5mBXwYylATGw3PXjhtwVzDDsJBKMdn7e5XcBQmeC8k66FI0qxYvwLC
d06Lpcs1opCOWqEkp5f3IHinbozwzal3Vi0xFCkAjwu5d6rqN4zB7Tl9+L0fXWTIBrHhqB/A+vNx
ef3o3AWlEWvG/0fbETYI1ygqYLXEcfm+777g1BEC8ijl9DXliwkxBMasfhabu/lKEiNJcH3nLy52
S3Bj+awLnonx7QOEver24hdyC1l25j5SQHrrjDA1EgdlQ02FS1g9GjX0elfEoIeIc1hZOXUf84B+
9AaLAVHYWI9pSkT6az1s9FqFYrbUjM4hGYCIceTZBZAYOpcyrwQ377CJKosgfV+EsN2ZatoxBD+F
CEkwqoAyryOnABGVNp5WXJoLRL6nimeJLr6AYUguXTLo/aOMcX1SbqK4EeC5/z0Gr1ZOUM7ojfZS
AKzrMuVmWHqy73HFPjyEInJlvlxb2vp4c1j6hItkNhcZjelMGdUGrT5lvUfZA5dFN3U+4I3i/SK7
9K8oxII6ddsb94Pg2s1gg8f3LlIlii1Yrtu/12J0r1sO6QYcXKTUqxjhWY3BNbwmD8M5SfxonFzw
wlFKViIOvj3h/WFgf6GxXKaebkdYoHCCLWhMGIxY7sQzSam4oPx+4jv/oKkW3PG8VwITlpwO4YdW
xWjikQC9JuT24UlwZtuT7g1wsQBCaeejvy7sbIkM6835LzRlxASLPWL5T0RQxd3DSO41ivDB9IBk
fAdlNrHSOLyop94ulzn21sIZXPDTLRWMCrvz7EOLGCF8EbDySBFvbt9e3kJt24DGF9xF4gF+WOZI
7LfvYtUXHlcCky2SjCQUcU1ChEea02MHY4+jmjU5SaIbohwUZXD0Y1ibtUTH7HO/YRfTfRe0g1Lo
EsnuIezi6QrVPIl4DNbMp7Ekg7oGSnnUado2iPtskJKTTpB0YNTNbSMvjluDIyqx5vqOmpPXYRyk
nsuSSBbGPPzyCU1RRmJ5TeFm1+ymbcS+6YR4SN7MpmNgqDNFIm6VhaYoyu7HRqsZIhS0LDmdVinw
U2rTrULr8Os8iUbZUzO5YJ31hBiS9TbhkVbGktKjy0x8D29wjw75PhZtYBtGWaYXnXYJLnW3378V
pUSbK38msgAW2hbSr78VNgYlCkuoVk/yAzmUJNFNEP4SmbAe273bSvIH1mom7IPs46WLBhxHZkEJ
b4tF89kluaJYErbZqT4cbddVsAaMyhvmzx7gwUJo5mThFwprjv+L3w2MmYJb4ccNiL5/CFM3GP+h
faJqnXZ2eaC5JdvKbOVL5wGg2Gaaa+YUf7RLqWkvZ6n4PY3gSs6BWt4XH9NXhCretvD1tgFD/Lmd
wxNRsuY09xYh7zGyXCUi8/CCOMyoyHzHjyvI/kW3FswfzI8ZfUQHfz8ax3pEGfEHUmDQ/56YiZP2
yVrEk66OQu3i2vfc+HRDR2b7EP/vDoHcnwaW+bJP3jpkHo6DYj66W9KEwUuDNvz0KPe++YDg1WN9
fBB1S9jjQeA7/HAlPQmZHUlXFcUuHKEFcE74Q+Pkesl+RdUNcyoFeBkuYjG8vjCZ4uu/u+o3i/1/
o1/BHeBHyrBzIK5kj9CXVEtIE/KjspLXY9kLHLZdPUnQi5F88Qpv6kAmCnyQ37t8//WuF+hYWm5j
BmAtmlFlYVnIJimkHJF4T4OWijtuy0QTRsfN8rebJ/6H92RjEHihfmZjpPx/gp8KD5WI4ZfF6sFp
WZU9jZ1eBQc4CblIbvHylBot5na+fuNLbL3G3kpfa+c0hY7q2h993vTQirH9X+ZKNWEr+siNc2bJ
9F+wFVjRqWFTs0mMmw5vpSLbFuvPciCzWwCgNgNjyxuMWpzBBaFSG6f/J0/DIye0MbuXU6LzpD6d
lMqKsmTQNV5hq0KO1xf4gJznXiJNhaEN+lEMWpaw7Q7BIh/7McmdzxdM25cOoqnLYAAg9oZErLHd
vR9mDiAgbL3k5XpDz0E9ZeXw0BpOBrEY8/dE4EggOJkCoClXNVvrmWmq0Sw5m4TDL+b29FEeRFMV
zMM/EHckmkvniwiULV8mURblwmo1+9GFGpbgsMIpHN8utRi24CXu7qh9c3/3AnmT1WVD98zVVjip
NB8kHPbAlYOrM6ptzTPvkvagoqikANcYtzFvtrnRJMYoTkSy13dkxNCM+gQXFSs53oWEfEMAqvdr
5PLHWO5UxAH8cc3TjV2sXNo0B4uRpDqqagCEoVisxTGjtaKdXhTca5AExhVgEZ25uvHyQg9RYpWm
fXkyTbbAAyoTaqgAHnNk59Hhf17xIVrSs3r2oVTmWT97umopkz5t5qN3FoPHyBQckmDQgiQB6Bq5
GiM2w3nCin1TDo1ROajdFk5OCbd5QMEhM03g1GHLXHBXygFrWheaFsGSS4BkHwxzWtVbGkaf3rlz
1HQxdlb4KWjhd9LM2/sWlQ9wF3s3cnM+8vBv2ZmCHjNfhfUrarINQCq9i+oPothv9m8GgQ01WN08
I/ZFWTDxMz9JZq6hjGwwZK2fC5og6X9yCoBcQrcEwmG6fCKReZJ3czqxSyPe/Ha3Hk6vi+E77thK
utrpmpPESsNmwk1e1kRcTEQGJjTYMSzeEIbS7d1FH8bkA9NRnsgB6KaICqjgcoRCDt9I7Yl2jKNG
V6OIpLv6iJVKv5xQrsxmCyrt4j2SHBg2PnSVvozeqUd1WmoQBEao91qkTYOwhp0Q1tooe481sEZJ
/YI4vvHT2zufdD/Xe/d9wp6rw/Del79WVLY8TuUctACtHz7MvwvPhjhOm53LVRmhvSrii4fbvb2R
t+rxdSxtXOLvoDyWa915p6+011gqmV1zCK9gYqTldBCv/B0xbIXIgr0qYTDRFh3J3lhWi8US3hpW
iUZcLkBbKPVKWHHntPVvlPwdu/9K11hNzJPLIN7MnBjuYQP9sHia/MWD6DjS2P2UtSOLuVbTVkZH
x5aVGO2hIN7DRtHPY46TMNe2j1oh0OH8DsS30IwUqnu8/gHXqroKjCYMkDpmzUIySFEiNX/7mEgk
bleBCVUlP0LY0D98sEWekz1G1m2gtLbdHwdU36gmkvCG9XagO0Vlqtgk16jqm+igcWMNRGQ0ha8V
ifNSSXIMXJKhwKtamu3kSmBKPWB4iREajZ+Aw/43fc7sKKhKl/4X9PxZjQd+Nofb9xIRQQ7RZj72
vI+4+aW4xC6F36szlTvRLRjrVyEhchxFIKKd1rhgWNooqwVBech/r6tv+2jTSJGj6/snOgC616os
gyXXqAP9UiMgE8UtDtGjr5sQsH3ncv9wqswuzi9Z9DLgheuXOovYz1bhT9H5VHBQ7gsVofciZjgS
KKg9CJ6CXt/Ar0xJwU5R2DBl7wx2bmh16wauJ+7XrKKdLkqJsK1pwT7pNJ/yv1jMuu6i/08p825u
3yQOGC4GxJiAOTZZt5+W+9PQRCahrjonbnDB2QfNEQKLfveOFfL/kadYv4r9Dym/eAjPVJutg+Iz
56lWON9QVb49lKAW9rPJA2EX8+lFV5rDfn4eKvtTIdNwJOlr3vGpyzgAH+WPaAdTRNwYQycSIt7p
HckdL0RwD+YGea6Z+CRrb+IqjTS/c/TMT+m6xJEZ5HkgA3dfYzjt5sx/pB0ZU95Rq3WpHE4q5Alc
76a/hjewsKZqW3QnwgcHcdJcqAPGyL5A+0SFFrdhwzJcSJ86L80seHIrBbefuzYLTMdSQdvcNqFR
SnfEEFGVr2alKDxpnUGkxMG0ajYOMoN7UKBcS/fde5ZKAtKmij4xddW0Rxr+cqmLLJ1OVwyvTKNj
IvbTfU3bwJucdWtg0WHaghVzQDRvECzX2/8MBSzZHB2hexKnePmku8EXyO3kNblXlDXKvtkIFkin
ytJc1dYMzt3poJCGCQBydbRVrXVw0ddzl4vEq+1Za658tYXziK8OTKSPnWf/7449pZC2yaOR2n6c
0NnHE07TnZtiQDxTTODsNIvAgK0J0guI0YNu+loK/018E1jrUSHEab+IBA5uZO6EKUUL1Pvz1q4H
d5LE4CDlK4F2dm07x+SejkfdKQsi3CIVrsJfhpw5sPfdwNCvW0ymmLvcQLDjUQd2Wl8pAQa/Xmd5
jqzWwekzlkYGGICXMwG8cuwKgx5+j7fb8bbDxMbhTdZDn09y3YHgETIeu40lMPRtuy/NU0gO5pUh
M/eYy+RoBDNkzOnSScV6npkbc7bZuslnHM88J+fcjHMVNdKI7bi9RUl7FevKnASN81JZ47nv2qXg
p5qFrbav05mWHmpbyA1s69iopTnoWNCvvBW/ftlGaCuLKutCVOLctkX4WLcbwvq+ElGc7m6pPJB4
iVpvLxDimYP3gJPSSgBSLoTg/HemO59OJdrMIwwfN9HjeFRrtJK3cik70hjnWRHom61hQTo+7pJh
f3um0nn/iM3sbvjYlOfNgm6McY8l32oLlWzknVVf17sL5seW8PJiUZNUvoUD2OUqwVrQ7eLVOlsM
0eVyBjUwRa2lT9flP1O1Xif55RzPPZAuNR7we1Fs0hVCeEEgspmJgYn0djyCOVpAQzw9kc9WR1Y/
cNFU11YIJ9aSTTwVExur4H9ZS+J9Lg/KOXz8lxwHBUJsmDjcYova2iB/T/xCVEJsqjn9UBGDXQyx
yS+3AQ8kpLFd1+7Y3WslRMoi81SUHOxHd5zGXvWBJztgc962J5DF00e45dCO8C1kqMkAz+LvOgrW
8qslX0nxOPP2vN+YFmT3eFE5icDfV+Y97sUycsVoCQ+iNQ8C5j50dIoII8Fj6Q7NbkdgAfNvdc9y
MaIwnnjHWNGv+/jmHgdxJ05lK01v+nVfsuMisqIQjZmPlFqmKYdWoD+wCtrErXNQETdyVg2DNyH2
lZzY6rkAb7t2LrFcI/ACcRQhtuUURTjZEX0Q+BEMmRKJSpEpg04MaRGFF8IfvkLRRwgvB5y6DS5z
3h//a2uopOF546FL7cSNExCV8btiXlrHhubbucty+ALMXK1g5ZGfxHWfXpn9cFPkaBBg0CNQ9BC9
ri3ht8IIzU2ehFVu+hpTBcvCELkrodeuU9gZGn9NIliB+uAVIRXjWE3b4JBDd/uY/CsprwlWw6zF
zFudXerAAG1LttTYCg9EdwzxGVuTd9JvvvPaBTZo/fBC6a4Xj5feiyH529+z5YH0enH9VBp/FxEv
2StvWgprJRV1yO6B+B4yA5VyJxESzoY8HVVRngS5p7wrgCYUd03wzGYnulhl7TinJjo7kK5DnkDC
Szh8c+kpPp8n5Jy2KzrOUwphIfSuzMwRIrDhKR7X0fAdTaM796VRngx49w3vVw6HppNWdANPZMnz
HD7wy5m9J5kIyG2CJthWWrl0hoTD7/7EZxNzxuXjEhOc+l2/h7KVed6N96J4oyjyg7EisQeomYtk
Jn7MjQ37D6QiX3WHy4C1Z0Od3Hl0oPqV1tzrhZneBIMg7AcJ2F6UnJD5sf3kKcbpQj10gZpxDEIH
/HHn1/15ig55NE7PXOCsIt6Sv66Ah+DjGqVkWtR4DktPJLTnzAIdMfljlWyrJ+Kq963D1XXDPdjq
Yh1vqq72fYc/QXxwsYweSorzN/2n7VGYvOX6dn0XAEi9w9RNffpaigkMuEoK8oM9p60c6QI532E7
vcf71B4Yzi2uqTPsfyPBn5ttVPVIab7DOxqOebvhR8IOQFayas8NFsut3PcIKv8lUInb0ZZcrRyj
BoGzvwAPqLo0LG4VOLSu9dh2CrKC+D3l0DXu5xno8lmWrfcpAxSzdE5MD9U4WP3xzDUeRaPr9xe6
ktB875OZKBB+3SYs1kxQxFG8sAVJyLsAiSKqJ24eQ4xV0kySlZK+yrdUBxvQx0GO2lnF7b08H+TT
9o7Lr3A+/FLP2/JcO7OnCl1E4D3PhSV42srhc1MoEkfG61Qfv90JSwg0oxOtO62IYxuR7n/BZxh6
wW6t2IXuW8bAXCgqij2zYpazO+j4jbGN+xTn5ztDvi9IYj0rCjQdAR9G/t+GZK9l20W8RGCxCT83
jpay3lr5bKtynnADZG9nvf073tk30q1TQyfiVczyxH2ItTEdSPZBcaPV8/kgtioeZcXw7PIqTLsK
t9iQw7FBKHYWnw/HD0lWoKW1ROefMilb24CL8ocqmppuRop6oD7Dfse+PDnnp+CfdzWHRD2K1MYJ
uesk0Wm84LgHNVJG5zP1VtkDKlTS6EYvX++Ok9gRz5XgW+ZUP/q6N5Xl5TtDqB/XGrMNcIiaS79q
V4HJMYQQPeBEyj4sWkn9/cL2DMKohB+KEEveGNdJg/V+1K/mvQl4jeP3ohI6C0yo8iu1eiZ7C9I4
PgwvbXE+ycFxmmKJVVJJj1qet5BQcNghDNTQWVLVDUrAOYP8Sw6VQgjjC1ntqaNpgRPzTna1B5md
WVAjspmRUArJa5Z8iQmqiHPcF+SSznx1Ao6MFphg8y6oWh7NHRBk6qhG82mAdUZuhAmR25wcRUat
55Xi7VD6+gjNazzEdg9f2c2aRZ/QMxTNQ9obUqNqM95+qhHmWBAhQR4j8FQvrJQFaKNz4V9n8Raq
7Pbrkxz/2pdOqRbEZ6N+t+I7d7LBeiRv2zOhC9KoP7EpUPdSCloxz4oQe6AJs0CN1oAZmJ98bElc
IBiz61wZOd6vWx0WcDGdsuchH89p10h0hBmAYxhCr6oO9IzcsuO68mBdzsAoG5q3iHnRpOPqOmab
rccJgTIcGi3ukEUrb+dt3uJVcoaxN4Wv/hfjGMK6faprlxOwtPkwX+74PrVNXIplP+hIlHrWM4OT
IKxjG1IWoArz8TC4DJM5tJNDIg2MMYEush3RG35Yde6yjoqHWkF/k1kblZLYyYK7s5tm0Q9QCpSv
NeVK3taxuW80XGyLLyALqIf7MhNw/Gxw6iawMhwjj31JVv7W1SuDjcVpCP4LrZVb57m5rptcAqMp
I6cdIn7hvP8SMI89XMN/tUpZLoX+jEolm+hX6JIYR8K/Wh6iTbYfkYiBi/LzAgyolMBtzlGuv6Yg
LwM+E2Fe80v4afPRNaCaYL1Z3fLOW5CvDaszxlR/4fyDeh+voLGMgviAAjb1vXWi8AR4Lol7QyRa
+E7ZyQSPZGfrOxKPWuU+JLeqCSX4RmfJzvWVaUkj/4e2EhlrrPGQssSO+Pto0gyIN/wM3IUN71VS
4wmwZ4rELuHmWjI5pc/9ZFWCk7A/PCvUd5longkSfRHt8I7bEMrvYhIGC5Zf4KhGzes1UPZ/zK+g
qbQxGY6UNkX5lEU0iG7RlvytQnR7t9d+Lx1PseFWGJv0FWCbEXL3nTNBDxR/c0NP0HkA34j97WKI
58bHZacJoWOe9nz4ZVooXTzd3+qiJgTD5FEHh+m+MQEqy1I7/vejS2/HdcgcRgvn/ftTrBlk8tM3
Eu/nqYOdJLV1r7H4sVlFEtSGj89xJHQ7P6eOAud6WNfR7OHV/lNXLh2F/nqVTC4+KuDaWYrlYRkU
2S6SnfmGjOxyBtzSNz9xAyq/IM+aXZ1V9u/irEFD39LL1w90hOvSOHjd2OcCFnaApgSxGiXsbSnw
9L5tQ16KOx9A4xwiZudq4V/fGuyjiO2wmjVZjqOxT4K1o9L4hB5uR2wBRxr5QtOEt7ufvrH/DhpH
QQfOGzZ+7c2A0IaqTpv9wSJoFGtSj4m1horqF3wQ4M9x/QVgWeDHLVbwQtZx94OEUbsK3/xROVou
OVGqOq9N7+PeyK6mgBRwoB/9CkNFAMDGGw050MQxMKE/WChAjWuuF0L7RoazvYtc6CSvMdBZ8Z7q
7Uu9NgQb5/UsJOBVSvCUeQhOYCqjLT48kce7FsW0p2hpwv4q2KiMrUiYZ/WGDFeFkuMSZTKpcFfI
k3CeCU33n3sINU2joJWGX+KMfDLvIVb8s0Z+weSv0hCdASwRjxxS0BY3GmboZ8z1YL0YaLFN58bs
m4y0BldGoKpqvRMJSHNarg7iLaStCyuUv5ar7/ddNLPcmvRXD9yTfBf9Mtv8O1UlL7sXVXPtAxyy
wELbqokunqFisQM8C8TMS4FrWcw8r31sTq5YMbKr6bQg5xyGGVa0i4ugFj8hsZ9q6doaHovkFlyz
+o5qt121R21U2xpMsG4DiN0pBB1+zcvP77PUkY+9vl6p9nI9bsyndSBy5id0iM9YvDU+AmlW3Ex6
l9ejTg1fd970ulyjXV3G3QwDaEdOGUDkke6fDPZmUuVZdIGRVIUvgDDQ5iZMDTa/yomoV7c+DQ3k
6FXtn35Vl8yA8oN52vHyVePINhafTMqGlV4dxJ9gKoUAtoEILW5vWOezJ5qU8Kl9F9+PzOlNMyW5
Rw4xL2FcmVzzrjkhbV65JMPH+MD4UWPrZB7KocqglEiN3jh788f5gYNX4IepuBP3GNTR0PPpZ7Os
IKqd0uHZwjn83zYLEf2kUK9t4FQQqQtTklBUWDAyi3PfB3QBQqWcsOfkzWRmotSZw5rtQAOq/ZDX
hGKyoUmKD3Ilq1OxD0Q2aN1Tujq6KrT7JVHafbNvi9oAKZfPXnXQXNFeLA0kLpXaYde4OmiF4s6b
4fl4tHGLW+naIiJReAZTQuZf1crjZp5voxXcyoJg0wSMEPLkDO/zsm3jTC8iCw7APQYb9edhY3IJ
bxgytjmlQ98dInCDUQDs8WRxWvhAcxTF4lh0Tqb6ViSM3BmcVBcJDmJqZV5E4CQ3ljlR5BQyZkcC
xOcOf5MQGtcOvF98FBL1A7Xx6j71Lv9eUCZQhEZ0CafVd3osmbI0Nt1O30+Hrs2ZuBuXNCV8w1LZ
94dN0OyGI5vaeciqIrVT3PA3Bl5zRnqYFjwj336PBCqDn3Nkajxee3vuqsUzcvAfK6P4KRVFfjze
G2Fl/KUsQkMd45irwjiJ9iEG/zPppbxuhd+DgHu5LXjxa3HmkfJyFLEgpRuTK38eMQ5ljB3roApY
eAPL/kJs6xBNXZ1Pqlnpi7HK6zQpRYWpPNMnzOS4GkZoMoArSTRLZQt1b1rSoY+ixXIYLvfTqheK
ArEPDeM6XkSMjpfHlNOFzjJ1LJp17h1PZMxN3ZOwTnZXrow7LKFktV0fnuZZ85BYBkbCiB0qLBcD
qCFhJRtoLvUBrb5mYnNu18ams18dmQyLFxzZUXZ0m0X1JvXz0A6WrBaSGEjwgfjA/+SrJGrNFy7h
/a62PDKXoioPq201G2CPRdizjqlN4O0qu0LF/+ic+FX70IBAMxhCllBFd5iemuDNKwr/3z7+226Y
kbVxbCgbN+YGKzgBDFR4W7b0qk7TnjYZkydP9iHyYLAm55I8QmwxMfLkZL2Ov1qnKf3PiUaoOh/t
Q84q5WymUA0B7yfoLJEK2EsqdHDYmwkV2fypjCUB6V2E13+PaN31U7JcY4BCJssGOYfMFISZRqIr
ZbclzQRj66o0mZv0SP8fbrylOApjVLTBWEIrEuwKEU90lX4fxfPHWB2yB/BMz2AgwVpaW2f20yPw
zQycEsnbi6IasEZqHRuptb5VA2dDA0+nCCLTuWQGZ0Ea1NAEBOCjDsGeSNUCcwLe9tAFiquHqDJe
ujljieQT1HwcD6SQiZfXPDR6ieFCnTnNwW8NZ/n6nkU9+kkBd+3u7yunp2SWGCPYgl+ayql2kfBU
SGPOSCUabU+p/AQUnU1DkhGtcMEmvAYqGnfvHAeugVp4B+U7UJ92wAPoLTfnwM/ByENw6LVGsT9Q
By2UPcF+vz4cbNl2IOEpwVN/+ldyWxZeczQWGQlukcNDWXwz9i0oEc9xT/CpjySmRwhTAkz1UBLN
5fAcI2veIWJcnalNj+2x07j9oXcQyC5Wc/iYedPatSa5fvtXuPmhdVAZEIjaoFyWemB/DXjOc0+c
btQxrKLJmnRxNSaZ1E4TjKPQdqL2OMqMPYCezIn0kV2eqHpiX9AZlQYG8+1hxHUr9du3UuXEY17/
UIPXV7uaQsZzHldP+kKo1ANlGO44bHpOpVJGFcRiQZAK1Gx4Vesz32gc6eBPiTXeJMKzRn+dv8bo
9969bViuXn/YyKDgyEal7Lsir9G0TSk7yfZcBR/DFc0mExdyhQDYlf8VAiYhnHI7wAeDGsWXfe/I
Uv77bXFYEMrfHXWP+i6Ax1Ire2zs2/pdg12rB+YFOikWCcr1EmeA0Kvj06xst2NoS6GqZzSQ7CW+
z9SVjgAehqqTnpKh/0HdIQ6tqMFALnU+hNrhi3qhpjCzs9eMT2L5nSS4spT8FAqUGNVJVWzu7O7d
KhwdYG8o2uSv2/2r7AL+seURp22nozQR8aIf7kby8M4EwfKq7RkzSOICsVBxz1goual/NbxBVknG
SVVpuua8RBQbZS7eBTQakI+JxzlmDEFpilz8xrlSDjtPS0B/YUKhOrP4IK66vr4p/WmEBy9sAV21
Wm3bCWCFNRhI2wjauHjb4MTjjTjC3vJMd7ambDZSe4YfHRJ71dPaOKYXysn25aApbJNjlQ7bQrKo
przy6c5TtOYDC33NlnQ4+pKzCbhIcFhWNDU001zR1REcwG3fmkL0UDkIb1Cj+vL3cn4BIQ0ToKib
vVSOwrf6MQH9Osjgr9Db2+9/3tg1YfzbsMv9WAUJG2IfJ8AW3HtnYKM/5vLam0JHXvfCeESb3pSP
5/9Rr5eGMXHyYgs5odIo//E4AovqT2x76j32ajUOSVwlLOI5o5A7BgA+kmEOr/6417XZ6OeXxfXt
5TGnLxdKn6WdZzzE/ANtf7ybVyr73J7zJ/oVeQUgsYA/MoDD0EIDfu5DGB2fqwRNC/u+ZZRyEQ8J
ncDAqZ2/aiUmvBoDeLww9ZkroQ+oaG76kiBtnnunISh3lhomDSoBmce8v+5gAGNCxu/H7VofBcSj
6g1DfyHzPMMI8g9v5hwpqD84T/3pAEQrGNRIYg/suhC4r/+0+7DyXm36pBEFG1zVkRkmByTic4n0
/1TIjJnSo39Rdjk95vslOZxMkGkJSLNAlRaYzK1VasieYNsuUN58ewMOqPalyK0TiN7UVAryZPMv
oRumLNFQkgod+mNR3rdns+MLf+3430wYVwIXvgHRQEboftng/TOQAv/rXbXdzl5jqOVCUzbFv5g+
zmoc5JFTv2ktVw/NYgccAFUTY0WfjJFEsAUd0BY3iJurfjjKm+CiW0n6iS9StvTt37FNRFRKJA9v
DzYs4RFdMH7cCt8aOUXKJKB8CKKUZHCvfiC7qqZqd7S0c3bi9e1Tf/Qm637f2VNeEh+AK4YFD77g
UZ6n8EMpP7av3KGtAY2c2LC5xA2nsUc/cAZz87+FWAFOSQP9jOqa/wBu2aznOv64XDRyRcaHecJX
habokVVSKTweCcra4dhiHwOc8zf/+xrLSkvOGXL5At96Bl937zZgvBtLLXdwbnvEqcMQxXpd/3d5
0TYwq8lXV0yorZdE5Jj/U/LX8WTjArWQIOVx4WIWjYGdzCubP068npeIqrN/g+6TsyoLzUyxFTwK
OaeBSwUfPbZJjFzTKe6/6HQLs2DA+O9HHCsJCIhuzX3tuCMJY5+4PDfH4pXn17kYLPCNzusnsS0s
9A56NkM1tR1YctuPSNemSw+slkQo71x83xXRzIMh8bXfUlPBmpV5KFNWURLaOLBJOu8iaFlI7ZkH
2fxbky/b1+WofbEROiaD1nCiHd6KjLyjoMdsEfkhaXxN4aEWnnv747ZtJaR+gOtmZ9BS2eI9m5Tr
n2fDREGAvO7rlVykB4CpnIft76n/zWp6hL95RApJ2rHdavOMzyNDa+LQ1ORX9RNpDCDs0B6ifai9
3xRKhs29fsl/3x64VSLoeBqqX+tS/Jeu5F8DSikj9l8yDJhE59wa3Y1I1W6VBh7KxY7LHCD8MXgl
/S8r0w3D48ZVxmelCkKfnFwYRsIrudGPm+FQ1q04tv/RMxP0wT7QSUUvqdvHjEeGRyPCuTOwwzBx
daQ9CdvfddHM/fTsvgJiug60wJYP1Nw8rXxUPMdLxaFkyknU0ybcFGHPbmP71hWc+rCMrhctP3g2
1S5mGYcboZbpzooGaqFCzfQYVgKmE2myeN8ouNZVbj7q/3V3Oh8eIQVQ2Q0Jb51k1qriki/L5wjr
LrknijA1tENN0YFs0iBKRVLrP4gpZq8d3ZXNBXQu5egQl6Y+K97HmFxg7HGQoA7zVh5PLMfkCDMD
Opma1gT/Es4zYfgBXcmR9dbuQf2Qf9RnFLCEQLHGnrAsjN9YaIGG6I4UST1//96Z02zsDGkODCbr
//+1O2sy6DCjiUrVLTeHDuQ7l/BnVD3RPrHCdQCzgtJdEPok+ddZiQwKVoaRscBVXBzbWAI6uaQd
X3TGgbUsRZ1A34igZdBhxhvjC6m6UDwQSXM8kq+HHVwyqzh3365Z08Ylg6uNmXxmb/YdFf7LhMRc
n1rtxYwsa7+3Zfl6eTOH3hVb1MZir2fP5pGc23OEHZCynr9gUHtD0GtEAqDOuHn7Q1jg7XG3/doV
fpjPbA/LPlgrSn4jt+rSL+kLlkqfLoR2g4I/sWaTSdCW7T5a28e97OghRm+NrC0DyDprtlt2A604
I46fIzM34O5gb/p/fVFtP0xZnvlrrrzBvg+FA9wP2TtMk97OjgCvS4teTmGroAi4uAuzFt08wHNZ
kMrad4JVYC0LEFi3WMY426W1TW81lhIPYeuEU/Q03V+2AGQmoChjPYKcPT9FASv75r/k+kE/vsrn
XAHwVS56BmoA23bqQ+pg9Lc53p0IY2KV2zo5jaFKkUu2PTBJ+mHg6125ZVgInWY76aVvImmLde92
bv4ZjQkHYnonT+upYVQRtGAaPbsRB+0NbaEtZmQLO0TuIvnhnAl8rkU6nmHhYWS5UFEdkZ+cc2rF
fqzkTx1sATfChh0LKC2k/KIcUtCTwwh3WvCpB1LE1tZjZi7lr8ihYy6Gd5DPLEA3DpWyX5+ASR8C
NdbfRL8/SlAIXk0GHOpg7KmRxledvnGuvfRm/T09upmOYjxqsJq0qfMozWel8ocCo5obA0KsXmkH
fKuSFNaoIaeXmDQdFKIjhQ9cGTHSuIuQhOpMKzFWxwgjm2Rq2Uq+rMlMPbeGBXtT/NyBI6QpwEtK
qluvbJwPLHTgYM1m4Ne964KCaxHqdEx0uHepYCC+JPWqaDHzS6v71pgO8wDb824ai+eFZL0zvPuN
N59apmYF/B/DKNHzS8YGlPHQ1lbhLTBuEstEzKPPKE+28NrCKBEFV5I1YnSS2kFUe6499Obs7deo
z/pTIDXksDvyTO0u8Ra8soXB6f9qF1PGEhxFLwA/6uT0OFW0fI/R5ipjJBNWHiTN1mNpPMkjppro
/g77qUc16Krc9ODB1TS1vmeCvXb7CqABm/ZQMGC+cxPSO5uYvtdgAF1LX+ay2AGhWg2hc11lkPTa
Fs4J019+3CLI7giK2ni9/qAr7bnXb2959x/v92JArCvOYPN3tNn43vtDgw7XJvvc+h0TdXg4uwlh
ScGxCXF/DyVgZiMpIJkFTg4CGw6uM3UVnI3O4MoAIcbHTf8BxKkOVV3PF75nolGH2kN/PnyQFn6b
7Tkifh/VohZ+mc/YVUD61Ld8px4GLEx9MS/8KXDQ1SxXtShuc1XMSVWxO2h3w6/zzSbXU0DMFI9k
+AqLehpe+0+8MndWKhwdhDBz6xerfuuHkx86ZEC33G3G1sqLpsgkrbBSPtRFnDOCAfemJ5pIP2MV
39BddSUpezTVHt5oFzP8/3RytG8h5l6mFwxayN25DvhxqjtTVsGL5V8L1IrmM61es+WsXKt+adHe
Ye30tmFORmk4WQ3gv+vu0wvsWeELQMqblXiYcuTNtKWdfqHih7i9w+ugUidpRI3Pscx/AY+267Xz
16mfOFTNFdNOMm0IFRcsPk2iyfykQjoRRGE1FkkA5CuDnCGpeVwVvTjmNdLpqgG8B6G+amIKA4hC
I25JkSor1khPG1jw7tEAA24zrNMVGTsQbn+VHGc22Lw2kSXGLpZ7X1yVHtT5Uzg4UnU9BXMtY92w
N6dXO0atruq0Owm46lFkN9oNwUdffNs58XkQ/DQhj/UJZS4t5/ln5eAKUY06NiZFL2wlC+OLZZqR
BjgEexmGfcFvzve5sYhROPsx+J4fdIZuW+ZuDUynenUKL4wYg1CaN3AdkHjOFl5xB2mbCFAhA4Ex
FKmBPxRobN64jd+6vbPb/732uBvFvHe46HbLCJGBREYpMmedrjgHmY0JOcZl6VEzCLFtRO7QFpg7
46i6wCSGnWc7OAvvbrzrVuA/kQ9eTlvJtjFfssEbL77HEIHjDdfqi9istDliCbBbszeTiVZYabUn
nOpkz1v7qwXq4HDQXDxMtP9IYsJcAQogbWUCl0qcQidwsnlDG2jm/Z+ym/RHs5QfoZlRByqLJsIC
1iIDyalfNXhu95LQgzp+yP0Hrsi3NEMZbWSniwVpAmDO5tm6E49GvR7i/3ThXeaip7ADtf82rDCe
0031I3aYUAPvRWjGvodHbos8ts7WnV7L8h6RYKfafoVTgHfBpYWEHFMDjfPBviq+cwWbJTaPJMwa
QmMDwoN4PblFj0Vhlo6Cl1kZek6vZFX8lzn5KbFgzwKmLgSbixLNoxPHrZlavRe7i/s9teDWcAgW
IP5JMjABVXhCoHa2srBwszEL3Vzgv7OWn+G3MOF8EjnnQBON8fQ6xrY6eXHNNAATAfccBgh9FORD
OHXvrJC+IolbAlIGB+gtroF/dEikpzaO2/cR17It8h1FEcTQW09AYAuCCiToPAqCh9Y42AthnGkl
xEIBF3/g7CJN6KnIb0b3Apc1C9It7edtskMNXskLS4UqEXeSrYxJGKamUhbHvpSOUKvSan9hYgT9
QONlT8oIIF6SN4U3XwYovfo4lQE9i42/KI+yDXsRXC7bOvNvv4eRjK+pze366Sc/PgWHhRkgqZO5
q8YjwaDK4/re8xUEfOjVeWrSq8MLMGb3LDnB2rRAdPjf3+m+wUBVz+hTSKy66rbKmlZT17Wpm/SB
iRVSsZhFhQYRHOrEGF5LIeQAbURxWTeuL24w9wxWsaYcsg0bSxCvW3YIdsBpXEqT/zPH8gBHuohY
dLKSDwtbSwGfwouPvo59/4WVt7AHmHvZcJfhIp91cHsyjfofriS/u+M696du8Zkeu7NLtcSRKcJa
5yGEzUvPi8R2j9rGNXx/T+TjJT+oGXaEZNMk5fFk9RZCv8LJASd0/lsfEoA+mTO4qilq0E3lV8NG
wzIKasbrbe3BkbO90gHqPHPh8OvX05kJG/2igBNqZUDp4hZQvjhKW0FvkBfdKx39iW0Dm0Z6jF29
/luqGJYH1d7JnuuReqoUQRsp4CDKr37EDSLKeUoooZMpqnOVOInh95r04F9Uwbio46w9fG+HGDE1
dli97I0YhmGXE/Kp/+eUphexvuQchLybyN3J5yuB+7R/GslbnP+nRiHqtY/O4GVAEqAwAo8SsnYY
piRQN6NItkWxDcotZw7pDOKpmhoXcBs7hz6TgN81dz93jSaVNPRpTZLoa5XUOaKm4J+ZhiPhakUu
7MhAi082nFZ2p3ZKh3dN4aT6d3VF5NI45PwWm6UIQcdWlYMZ7Ygj3hoKdnebTHVv3mjSnENVGK7A
e8YbrZUob5+8iazZNlxDGKinKWTaj/9aNiAd56xkVIYkfvlqsAzfjm5W8bgILA7Lnzn4NnmjHKtE
HLQutlyp+FpTUahZFTWN6l4s/jLEpDgrzfIxsJLGDTyhkeMH+UX2bzLg//TqgPy7Ed7kXTTIRFN9
DVZY4OhceJvUYqlHcLONa4ZRUhJuJe/jdqSckVnLtpt7BuMpAZVWZnx759g3a8WabWYZzqdRGiiF
e3BMkksKYwPe+yFiXzQ643YfxLaAmKkRu6mby7IisRVSa9CgGqrvXFiVtM6nDUnq/z9ZNWreeXo1
dplDVsTPm1PCTcCSDlw6k/d3I5oANRqwxY6VhSy7kzIdcfEDQvFzkGYw8OhIrt2PUfXI9rlEoC2E
DrhHI+TfdJQ+a8ghWEKPNHzAKlruYbnLTWE5FM7XxCjuPznWK3OoR9WOHKz0Dkb2J/6p5WkC/Ni6
WutAfV8EANdTXtA0SFMLgt4e2fIeK4rFuADDet91ZINyqkxetJAaMkmD2D9lqhmtW/xDzHQQHOIE
IrS/p0gUYDqavP64ruGv0OgoSZfoO680/ZCMR89tldQp3VbA1FA43LXFpIYcmj4ovH9Y0IT9/1Yw
MV7fiINf8d+iW1gYwBJ+u4dIaZYRAuwWYAn9DgbmiHWF1CwG6FgSkl1wjt9EDMU6j1VliMQIdScG
TNXbUNFo/oHQupdIB6VWoPOPx1uMOcqdDkKEzDjpCcY0axS/YOSDljnOUvNju/HCbhwpTASjD2m5
b3c3FRajddCwiKjrLyiAAqs9ehcEORIo4CIShtS0fPSqvawkIUy6oWA/5GWwQPDee1mkHIpU+7i+
EU6aIHLQaZpzTixNhfzKCH0w+qKy5xshUF9YX/6P/4pr5UjUAIrITEzUZXCGkP++deWym0vJNlz3
oDBNfylZe33s8iiAGCk4W5vUK6qSxh9qCm7Uwc/Vare/KyaiJVuFIRsg5YSHVzcuM5LDlNaRCEId
bPEYDKcIYFiD/jZf7sYLxZuQVd/wPNnVS/luNKZy7YQiYb/Lu0/m7RXteTHcJH+aJ12hYiqSMTcn
TTyUoP6D8RWnp/ndFO23YhlbSVc34Dq0JzIUmzkWt2p4j43zRoeTPwbkrPL2GWX85Oom7f8Ygvl1
VU/uv7kBzwIfVhkgoQ//RQ8Y4xgP2NZA94I/9aRBJ03CFhGqJMvkC13IWhN576Jjm0gJxX/5mcB8
qm8bjMFriIKSfFslIkbiCkOaFYsaEBGNxFUW9byzqxk9NhKQCUwVw4SvXKNVmLgJtIeZPgkNXgvn
P4R60Mt8cc5q18+hJi5WTS0dQW4JVzPBpSsUQIvbliqts6NNn7DzsUcT7G1LZMXEyi2UjJVsvK2E
GkQ9IqiJDGm1XHBHhWjtNn4vvBXqNDfCtbnmTWN+PAqEfjkHZ+TC2/nJq23Q5d6NoTgXBQ1NUq8r
FpnVqGXbVgeEini2OcInQmoli/81R+OdkQVqDca4gsG/hHYqyufHPEA2KcMZBKV+bONImmm5pd1O
jxnZZOqFs0oOBODQaI6ZghiMJ4pPxU1pKnyKNOXjpUL8J3qHKlsuW7HMo9d8n9CvryEUtdx3m3fI
8nNMLRCrhmDLXewwVLVi8ZM5CFQRQov0PcBBKnzJsjPpcAOtKvUHql12QaZ8ykOgHJetd90dFJ7o
Ptj5BdfjevNID0vFp3NnWILvgE7Pg0MUi+TmHXg5IAtLfisRHIdmukPm6fvwpyGOXRlEffiK+HuQ
q2mBAbR9WJR/EdMByGrDJzwyTpxxspfzFd5UsaoIXNleJM0ClWcA9yaTBZEBGOuaogYOJW0Z/eAi
6OekaNu8A3MZ4vXrS6SPLOnYGkqwDJCS2djGvZIVEGJLPmMKWESUxIEh3i4dZvvHPry4G3+dksMr
lCEmZnlScyGm/RMhK3GOj2riv2iCWqwWf/dgMDGgWNnGKezNia+w9I8g/eBfooTqHIfI6IiajauC
jWnAFB0MLlFnjp+eZRlUCGnGryeIPqA0cg/9S7GeDRq1OjIbEqK/Hbd9ubEdNE2HtjE4NwxNulS8
46JBlCogcQ82Agp6i8h5vIMg8OqoHN2WBtdgB2UoIk/BFH/xnfIeUktHlhycwwl2sQPss0u+jWpt
wPfdBORSsocnmsNwiuWmftZTyS+Z/p7Rj2hIRXwaw7dUEGx0Z6tjdV9XZZ33pENctq7OqyVoCU1o
yu7fLDtDEG12+cxACaX1rziaofmiNJeyfzggW3U8Ovvw/NALZqm7eCjSugvqb9x1b5hMxZSlmwGQ
XsKjYw6BWsqtwykTNTLCcHrtX7pYB5jmEnZWLMZ+TuTnrYXw+FVX9+AENOWgmkWIm0kk+C8gNF8u
70SwTEvqJ0u5CJKqLg4psWh+ROlI+4u/MI5867j7zXSwxHrsxLvD3dfxyKy49t9TJsLIukqLDXFY
n+Bav0ayMa183h9TtPIPQavdq8wiSi2N+tgYnH1r3IAdG8nJbjuSvkwyISzD+yI3kGNpzZBdQH1g
DrozjkvqIZ2Z+unhhYuZgOZcJVbAXMlXzoG5T2u2w7S9L09PjjAngSttSJzKuR8+w0PkeI8OKhdO
wBKh0yCubfE/h17xZWh6sO4N6qyxAEntotnWOMfLjPlPLx7pd72QL7v6tdmi6yuNwnTDRsmAvSl3
LyVkuEh8p4hyi9dreR57goDMmRbNIRXnFLkkJA24wSShKNStvpuPB2A9e6nwGzrcwMC2mAm/Ri9K
GJm22V0YMeYO7UmwZuQXBSccH9pntfXtzOus6TkvVdJpYxOP/CfWffTOeUB3hQROr1CqCDgHos1h
fEjHJHEGOkyXdd41sm8M0Uv8sV0VCfdQoPgwZCXpGN9pDUEiLIEufxJu67F8GLI0k82pwtCyS+6j
52klJ8SENysrILiCB9IZmboOZQKrNkVimHsYcmoVZYFCymhi4B8yDr95AKLWngtSiCzBaJN8TBAV
8pK+2y8WvWj9X0S1MRCUmL9o9UBywWQ3VVm3RT+BJqybjnDwOQunpEOhH2TzAAvu0TUCJGVth4GM
VR4AcsqS/vu/O7C4Z7oDv+Dp1o7yEwgXbt5LEN2S4Yu7geranmmEBezk0o2DDMnpmU5Nu+f8TXAD
tvtyZvqp5g8EUTZ72lef6K9xc176045MzINvgTyVQrw1xVpp+hMeiW1wvu9hr5vcYHIlVqWZzCCU
Xp8LoZBqfyWbBaSTykyLR/Mj0MXenGYGF39eLGLv1/9wAdevQ3QkVjPV1ItrV9G51z4nSsabAKgn
nGIzcWlP2u5WwoG0wv4JKFgy61fR7pFY+vDNNSnr6sLbQMxEPjSSrVttE/mMC9hWa0tLep1YQlUt
iwmgZ6p0BfyN+G7KaavFNiDNQ7h/g7GmEBx9K3o+xQa+Si1XBR2mcWow+Z7thWOjGi6CbHCGiUbz
2/XnRKjuIIhDi+0bEZplIdOQRmBnZ2fJnmUakcw8eiuJIlxiDfaIK3S3WbxpnZ+drb0te3wj30Iu
W3k0S0nhYXKb+x69KA0PbN8Up382FGeM7eI7PCZHlGntmEtwRi8jZZNk1y7Fy4xfG6Nf3sSA2SOr
4cfT7NDXl3Y06P0//RAJuAECv7GDph0Ne7quRJghHQZ51PVFKXyRPpB91mKXLbFuHlm50Yho5eF+
T4wy+sOixhFS1jaxL4P5YDBHlINh7qDsX0jSdSNMaS2dESUqn152NZ6n5DdpGI3N8AUduww6rw3n
VX+fJRS/WFRnyCC3FN8Hq5Dfevl+3Q113d7GspU2BjMaqcPgSxqF8MQg1E+taIWR6XypKvYawmI5
6lYShhk8Gy01bn8z3coB+IN5XkTtB3weS7qkl9zkYBzG+4ycUihQznBeo+IFEOkxhBdMBbQ1Z6qI
oFC04BJoeCJz3bo3KIDGPXLFuWr0DMWKAEQPAauB9waLVAD0RJ9hmvQFJBTc1NmUWdljzE+dQXHf
xcpOyKNFmG//yDs6h4ACrgXD9TJzFKN8KA94DGPnI5haRurZz6wPWj312YEJqcC7L97y/ZQw3fkG
uZ7AnmNKW0PTpVNNx8zvqaHhTPeTLpfR+uqdvM6m6PUaBukeqSaM4syrlvzHgnWN32KowwGe3FEl
Phm0u/U4Psxouq/8e4JVD7ZC4gI58Kq0Iz2wOOKJUoOkApTZR7lJsnwtj4669BpAz9ny7o7EJl+s
7hXwtTL9k3xJzjLOuWkzEqBUhZXKvSqTrMCCc9DSEUApqh6Qh3BmRynRPQfOkr2fvjgH1NKOuoHn
pd29J76fSSv6pb2awaZlJVKY3FlOIZ9Gu9g6oxxj2OnTvCU3zOGcKoXYLkaYoDuzLhVrw3BCJ884
wNgFtr2FB1ykj5ep91Brk0lysM3EcUqhW4dt/NIqpVTkAvJbyC/iKLuVyIKQYGb4IY7rjRhnpKZl
yYp3wxZq1Wft/8EIpW+fHCzl+nyUOjELRnat0di87IBj5xc7XpskPCMm4OelQLk9RhnpxwQGq1Tw
WBbOEtBhG8eM+7NNDA0XcPqwgCyT7IA2vIKuJeA0CFA0sbdB3d2HDWV2ZpgPV9Xt3p+N91+u2Bbx
Kc0p2pl/8Iq8vR56+XLcJ6N0YjdBCXqCxPP5Z6fQ15mpBhMY1k4/UCqWcPxa/KpRbYn25tPNoAog
bfWY1uQTCsuJN+MdOPbyjsOHsz3NdrT3Cbm0HmnhZKPivyEi2k/+9QgiVVCZHESiXxkH0kWxCr4/
rHlMciWMAF4pAVT6AD/Vb66DkDAxo84LVYbYo9fWHuFZJiLG2guN62yCtMvTV/+tZRWpGoQ9nMp2
LBqdintBSdkdXp9tGXKuxecUbvEXfj5wSYiU72sa9102pVEtVN8cRD7BoqmNcdKRABtW4eNP4rtO
tleO1R0fpZ5cFUNnWEYGEOgwV3v9B/vxxso3Hv4ygq+e7Zu58EicX7kSny9nvGXYlJUB0CXyrXbd
UxE0IQyl7zcdjBuxMLd7vU+mx+SRdAw0NwbxmGCpHV4I/uin1aPygnPJjT2Oz3pmzjv1tT2D91+z
sL23DzC19zFa4YqTe0KzEEXTaV5wQmgpqY79hTfcFLewamA4FDMW7kxfVkxzfjtwvadm1bGCwHrp
uwqF11l015MwxbJVbJQTnL7W/7J6Up3PPgXSV7w2TuKIecXHk7rxBfTEGHpd/mwL3J4q49KvRMqt
eZbspzMGCUNa0oQQOdvp1nxkig1SLyrRBAr7eN5XuwlC/ictFtN+EPJdgzynH7Yn3YkaVEB9i1DI
N2kb/LYP0zilthBDR2Ulx4cro15fQfc5JakceAjXd42KTq1ZxdvuFUG7Wzk06F0658stFe55m7Fs
3yhvGAopu363Es+okW0PkO3iNrXOD35WSAqES6pwIDQ9EFMy2fR6Aae8bSd6r+OI1ZyoSHaa6og1
uh7vHXe+KxTTkkNGcC5RKUHGmj4fRLPj2khKNFhOoir/vhnzlenjXm2m02WeMX5Cy6zRsF5K7/Cf
lNS2WQN7zzEtVZOA8eCsMv6N3XUgPSlstUaYkJT91Hj1BoeTWbJjDQ9BjYnV5rMBAl4/mHg+focd
PT2QGrRkOdsCiQpNin3mm+zOZs3LxONHund/pzQREQjXq+ipX5OIbK3oOadr/NZ+cDARbZCeApw1
6H59OUIbi5sRVoVO5oLdPnvv1bX4itfTA227SCsfVyIPFhMi7DNmiBV8FdHi3htZJpg5NARY4tNg
zd1+hEuzrwibEr7dJbIoJYgmsoZskSRnX7tg2v8Pv+oerv4MIMRFOihRZCNKQ5Z9OhVSFxO05c8y
DwciI4U736ubD+Vz6kSeiEMMX9HM+kCVNWS16b9Q8+gaPiYYoWtggSZyV+tm6gPfWG4tbb/2Pu7A
ECGqD4NVSUFKd2vmufmnD7GBj+Yl2wofihi/5Gil7L1crJtlkPQR4Y4v69Ivptm9xFYXkDj95SEy
1c0VaD+huKE1BoSegztakDVI3edQe6E0Xjf55fhLCIYAca2clqyDMHSqA6RwVvyR2X+z6385LUPY
9VIff+w0Tvgjypb9Aa3iuqbnTPGh2HrwNfBPvUQepsW6psCS+vwiAbA10EZEiwOMbombTYrgu3gX
ItCzxN3PmdtkMTDLJeq1bR6UpckBh7nhYYic9XpJA6qLBM6yLowEpUzGmDZrOVzPTFdZBXeRclKo
JnkGyRqlzWFe/hA8QTzfSNo0syrx/0uhUEqj+9ahpQi7lYH+6UprqawElvNHShMzJRfbm4DLHk7/
nSj14m9s6gV4bxpH72lwWDBQiCVSJu7vLyq2eUbF69TBNMHn7GoIzVVqd8Yn+drmBVF5Ehq8EGku
qFOI9hpBslXd+kux49ZGWcT5iwPJhy/ampiulH7pu66pBlSzbPCxjGanmmsrNQ0CyJdlQEGuIVsX
s18GFiDXpK8ikRgXC6bWqPX8czdE0JRn+VFBYJTgHIhitCPxE8unmBBs4+HH+mqMYoYYtPvh7vqs
7kFIrOmGeiyUzXIVc9uAoYhoPpMz6OYXa66f+8F+zbe4W6m7ee5ofyQUO/3PZqXz71wD7zUZg8Pu
QyFndQMODiDx8BwitjYkErBXul3OTDRzNp7himVoSXsu+87l51i3wKTlKSDmCRShLJ4EV3Yr+Xav
dKicKymAW98Fs8Hc8A8XJb9TSe+Fq8OKFfNh3bxLFHU7SZb82eMVCDUOvYofnWvBQYP5HB025Dt5
Ve88L5Za2W6Qrxb1zepBPEwnCLXp1ttpEyTiNWfwc6gBh0WLfcnO4kGsLQsniAln419sm73okSSH
pspM43iTuvkRKxSaEUNgsGy8xPrk3RMKBx8QwAYvs/7ZpVjnaN1L1jVncr3tCsqQJNmAb1yUO185
I6MojjwaJABK0cXr6bcSe+hwpN17i2kWGw4o2cYGxz4Sb6GI4eA6KmkdjPTfDLXsNcMJDmVFTOir
fFdKxjdITZsJnvXXtjtXx8RfHAo9PMDRGm/BgDnNjeqBYWVY9MNETH5MtoBJB7uaji6yRwvcmNwM
L/1moX4MZKRnKbENSp86owZoRsCOxYuSO4XJ54GqJjFHl0f+c1v7ylL1qsIlQ3yGqLyMBegZ4DeA
rRqM76hBlgkS49eQY/XaZoHJ9b02EZTEmFZc/itBSocqMwfAyN4UjL2qRoOaAfmjAYbN3dbZqFrw
FcYxjCGBL7+foXLZKNUSiOXOxNU5zkHzYD5LSInZGOasTWv3yIZbrPtBOD3Emx1Jz0eE6WFzcHHM
cEqNBxZXZqGa46bCh8mlitMrlpuTcYWCus4T/tnH6pUraWwI88LS+XPb95mHbRrr5n32rkKUKit5
UGkQB+hjRUhKHcGTfkjWj68ZbtLVxPE9hUEL8MhbaCZVekTufJaAu8W8lnEqr6UPWetO75AT3wos
YevqUyacF7/iUWrEm+XCQof8gVqJVxInwuToKQqApAijtXwwP92uWhgoOhgN9YSugpJCyD44PnYo
uNT8BuzVYpvzbbM9xRzUHuzqYS33cHoi7HgsbCTk2v/z+/aFBDxM1lHypOMxWG/bYt9LJw1L4X7x
5A7gLUm3nmAH38AZF2T8oXrxIJkorVWrlvftf9i+/VNlazeS4lPd2saIYerPJzxQe8OYKB7jAtt+
Bk6CqW05Yx+UCDq+aYVa3uyRVsOp4dMte0xVoOkFHSJlklHG14CE73RqUF1dSMVs9vt+DzCJIJbh
MJ7nki/X3jQam1lBen1TL/Jm7EtwsGAIl0kWcIuAEsFEokwifQuR+fLXUMyokMBX4k76x6uN0Zgj
ddgIJ6Zyk+Uxtr8auXvE3FNW336PcLi+TBkBxIculT0Oruk8MHIdpYorgpHOJfPu9Hc2KLsdo6Kv
+d0wn0RKsPBo3lZHe+/Oj0OTBNxUJJ7s5k6SWvhTvp11vTXU54GC6WevQZN4yAhd36l3sUyiKyA9
99v7VWTy5X6Gj8dbA8mWESVpWxQzZj0KBxz9b5dKK3Ab9HGi3GWX1NmC44CNs2P8q72Cf3fm6Vxg
6hmmMm8X7jqUq5VZs1uiyFbfIg/NgA7Y9vg/tOGudK6karf3FfIlNzicCgVcTrmu1wip1Sl6RaOW
4K0flXycoZ2Q0aU/rLpYbzpxwNMSRbznuzbJ25AWM5ZMSuMhnuhJT5FTUi/9vPxzEMCGQVTAEcnK
7fsAefXhuCNlPg/QpIf+1pfP5pZ9o4PzpHqgZ9PbSn8sd/ipSzLOWyaMp5+pmsLbDo4h+qLRKcoZ
86MV/uw5NqEqGFKe3jUZJT6ncM1tzo86s6GLuZT//1/GAcK3g5WWfCT5UYw9bwMY2YI/n6XezZtt
vfCazwhnDCsBfocp2OqzqJNxfrM9AX3dQqWm8ygXcj2iuG1OiOtnSurRPwGt+PFMfBlt1oHJS9z6
buuVTPXechbuXQRKrux/FD4wfl41b9y+7wHlMvrzgHFMKNUVNkP+zpAbmal4RHiI7FNgHzBQCMjK
nBY5nIoYzhVfSJ++HntvFYNEc3akYzic4cfK8+/BDAHLgutyrkJjjo/DALnnxY+taOv2kcqsdQqq
GFxvP+Kq7XSATYyfHi4jQ9CCwQJcJ/FfiJxSAgQUzIFhi/rVAldwxpZZJxlJAuBxLjtM9pABoxVH
edxIboQHXzLUsPn6IL7lHRu0W5OAJcARE7ii3xH6PbcowVBTJW8pwkPTVRld3ug86RXTkDO6EGY2
HXPhjPQsx4QhNFyMa1/vuDFgqrmoPG9V/lGHbm5MyfA6fvQ4A43J1x3YX6pQy2tEIO631UxuMUMb
aNNV2P9UiIp2GnriZ3GCd7uUexRwsxeMsrHvPKNi6jG0rEk41rMqxRhSAu0WvXc/EIHWGOjt4D5R
isJ4PB0O0E9Wrb15KmnvXyG0qy1qZsZLSP1g2dp479qa2zuUEtKWd594nZQOCKCw4sj+JfNETPqO
SPswFvNLZXd5IL5cYg0wCqW3cr4dBACa2N8ZsVbvymLTQSpUpBKCRyHC/ux2PgUfCgKtLTYeSbqi
FQhzvjermQb6EziZWoX342z6E8EanfT2NoqeltbwDJOvEMrzgxgEZnIT0m4AFEXRUSJvzqoa5nKI
idh6oPiaqME4oxljBPIg5h2jR6onWBNeE+7uu8q2nsGw+WszZxT/+e+YL9URV8FKIwWg1GvKjQyu
0JKjlL1144PHnLO2jfShMel1+EOJdzGYfsx8IDXBOebemqoR6+2N+ZDGiJHmshlt/obdeeNbDw0U
I6E7wghmPgK0WrOQIRel7+qU9XB1errot9dKqGDuimeoApEO48lQf1sHRgDVhifKCaAVLGn7+TNb
WS6YmFWoBTG0WNctxA2xqqFxGkPJhxtZtxwSFDPjdR9koMMCR6UMd05sTl+SFIeFUegGAtbXebPS
D/iX1bs2Nsqx5TRORWbGF8vHbiMiS8DUehIHzSgUmZsf/ZD1MET3u4VEphcUgrdr+b18Eowm4lp8
1yV/HSLCBJc5z5HnHSE2ipcB+/zouUw1Suyv9l9RA2VXjiYXfcrmSYqZVN64at+Nq3819RbcTkW9
lppRwsoPZruF49MzoRdYvQJ6TepqhVL/7jec6JT0VuGtcp8/w+/Cf1sS606R3Vq+E8ZQpMOSS+pd
7zAJNx4qCKQbCIcQht2fUEwJwcj7D2QRTj1J7vjYNWwN4+2MadqbuG/iAvB8bQWCF5pZg0ifD8af
pXEeUhg4bE/wozCtKjCDlsrKjFlLvclOpaKzbyDMx+UPa5lkCUw5v5MQakkJ9VpsBhMIP6EBjL5x
elI5/xER8czllfdtBYQsc2D+FHNwHg/p/I7gQEU4+kib6m4MySO4UPzK2dfKTmxTDTlk3DBwtomp
/vYQfJnd0+5/OZT4MpPP9w6pi/80ZmJNfwO34lTK89dwBn/sHS9iYjvdhQUAOXTmrZTDS7eWZKmL
xKF9b4bRQRXzy8Iq7UcNixb0Pt0xaUmZ88b7vdlEhnm2PPNMAAoeEYet+sSPiSYHPs6uiVYYMgnE
dyMuRIrNk99h/ia5A/vK4rIZALcvbxbT2dGxdx64FzodKGO+wTUfL7RTjnMLNij4NGni9mnpJuMh
bTvS/M5DP3Y0wKNdmJUN+Bk0fsWuPKEIkVM+o/ricJUOi9yQO6IeQ0Ng1wk5JcZavumAh05wKjiA
OMvBRN+4V/tJ1y5+rCCGFpEI2JCjE1k4sn5lziMv8ssn/xkas12bFVc+VYQliAcoi099L61aXx3B
yHzLMsl6Dmt3V/mVSRZW64UBCLE+lOPI5yHSYEr9OitPYF04fF1k/nA0LQn+r6P/znBeZztva4VY
a7ayDqma9vDskm2EuNW/4Pszco5Gtu6icvF2h1EJh146qL40w7r6moy+E09vcjm5xAK7Q+R/7SR5
K7HuEKhut4Cj7RYXJc4C6ob5xSYr/Xb3W3eO86ttOMvv0POv/V0//85yThvz4luDv3LCabCVhkT7
Mzdw72vlo7Ct/EGLRV2foiRwX0MjmWLTKiCY1WCo6UNI0FpRpw+QzvcaX4XozbbxpSM6ka87ZGas
OFlsCD52eniNDXWa33JBHs8ag8AkUoU8UtlWTuyTi+8E/sjLmUUIF1TYb2q0aHESM9Krq11NuZ2V
XAA6qKHXhrVwSPcLtyd5cQf6OpRR54n8P166gOhjJ6BtN3sJKf+he1GiuT2P+gKD8ee2UtIOCHbM
604J75TWWwfixvLE1uNBddSiHtmDMz+jqo0tJJ4WDVtjnanjD9A1gQZx4p1ONo5obap/QqEk46yr
SP/xu0Ikl+6CgZ42d8n/y4yjJ+OBhPBq/0F7MRkx1iMPWzB4qgulCrLnGRV6eXwHADcbNWq62UHg
/jHRllrTWCafUEoijnZneLdNc7+2dijH4KVQXNwQxrvBH5Xpr6y+ukzc7WH3qiyYLNh/bMztnLGr
MoYF7n55+d5QgmiAW0+QZXrEzAgTvKahCQKvhDrlcFCy6O+LKOC772cMNLgW2k2QLRt9PXn3uz4X
1rdT2f0xTRWhlhmF911jGN5w1lGGG2LY7vUUaICHGdx47sD1dRCcR0hmI9Aq9xaMb1D1uRfRUeFd
xgaK8vBLlMlnR7p4m9Mjgl0Nbqf5oNHPuoK10Qlbqq+n5tifAJL+MOenUcFhUeKCq8JGoNxWGclw
V+axXKtAiCH8RbFWb9NZtHZklTucj6scDu/4uDsauu2zhZ5YcnltOBvLUriHx56kutdnugyd6MbS
HU7udxklAwT2ZaNouNR6fnnUeEP0os/Kame+XZGGilXTc36Qc659G+A6nZO/Yx0p56M3G+NGYfhM
kLNLsZklVKK9E2PZcudSOg8D1c1Bn+8FhI1SshNyZWkJkA7IdZgfVYXTYKyA0kNOaq19MkwZ3Sc3
rqpKMjbWS9iBFyEEc2FbObo5AbBjQalR0xNTLhNGDGvp8+hcnOsVs5HQkWqgsnDi6GECENmj+0V7
AxUAJaLzpF+t7ctRwnjLNYTnpmtY2ficUWfTMFbSU8HsRJxsRwRlEKJHdLq8gC7a4DyS6I7zqXbZ
qUEb/f/bM5PNEQ2GAFcwS9WlamKhJftVoZO6tTHFbS/waKheM+9DC2wdT+9YCj7QCM0ZnLhRZ9WK
ppNyclxpClimXrVHwYC27PfW8r8dTibhVqTrqO6gAqC5ilDSvVMgN9IpsJQaXAxdzwhrJ9I6vCJ8
tCY38mZ2G/hhRP/1PAP7/TQP/IDR6NwD/QqTEYPGFr3LvsUNxDUp/qOuXQbSVY1g5iXDbr0KmFrL
nIqliq6JyseWg40UfMAqPEaJcGV8dvzI9UXH6BpQ7zz9C4t7tyLZanDk/kZ2xQKiWqWB54GWYySg
PWaTvjBTn6Qoj+k63Xwu+KTQSDbdCYO4i+C3eZolwcPvLjmZhxf/cNwBKiC2YSh5CYW/1wFthbuS
k2M/pWafpYTV2XP/y/2Mu8/xZD1KTaa9Wd2RBEI4lf8GJsK0X6Vgxq5OXVjfqOMVWvTGhPxZZApd
anJ/jkF0oqZ00x075DTNboXQiydv6oeaAU5S3/6qGLkjDvjFzyQiJ1shafaNhehLq+rnjbLpUj1u
AQ1LJDttXQbPkMK48bTfvOxTnpIRnq+9krHTo7ApjJkfv93eJPRg+bbI+hSjr2TpFcjhg6pa2W+H
bRv5zudMWyv0YZRaKKNFePxnE91952V4r/+nr1W6IHRdpcLJTTxd2Gky5Jxh7v7PlNh3QjKn+cq6
3at3DdsiAJzTcImQQL+pc9+r1v9eg69MD+WEg+ipisiusqbzkvYhc00BCQIe/yNUBTepExOdrZdp
HkpiS70JOeFDggeMeE/uO7AUgYYWRyaiKiVM22O0YvvWnBmFY7YncI9ti1SLVQwV5wt4+3swFV6s
RSuivmSr53pKDWqWT66Oy4VEir5t1ItHjJpB4UG7tXEdtFQVb7aYWGZgd2gleCMS92o9efNmiwz5
FUa0qifyylvfNagSW2tRj+VI6hRBV146nLr2BAf1ZAoHFJ7LQ+gQ+dfmrqO7tzCX3OEQwntI4Cb+
4YGFk8POFL3tqqn6m3IVQTFwFDIrlZDf0QwopVwVzXO3F/uDXgmHrrzCq9VmgAjgFXdgowjk3gOh
9ttQOxx229LATT6uc34Eu8nXj+iypUHW3tdZSHXFkj0TYH2kQ7NjiI/g+eRQSl9eE56g5g+TcoXD
uo23jqnMSVqQboVSWBsYmSDIAQCbPo0NgPOXSfSfkNk0wL6+hA+NTwMh0ytIpgX+v2kFI8WLNAN/
mQWDZvoWHpLreEBitBW2nZW0lrPJIsJ2IqO0ql5Lp0jEexC47nyK5fsXz/kSVwV6mj73WI662HzH
KSnVCJyqZeRi5ks/oHTFOAFn0WwK3xmV2U3faQfzeGykcteg8lsK7/Zf2ILJgxhB7YozwDwwnzXr
xNogcsyk7zvEFMPeZ9dAUqohlt4rbrUjhfjEti+zEirYCr9OWgSt2cN0NSGxAe/DD9B/54ZWUKkV
4ZTFmwI7Fpe6YPvmpqlXravm8oFar40vZY1UxOaJezWpFKhCtrY4vIP+gwP7iT81dJbvMufYz/4Q
cAeqLHuqi5w5v/91F8mpzJxSWPzOQBABr7OGXq/IA2dsfYebGngQC5Q6iZAqpjWuLTXjL70gWNis
ilO+WumLRT2wVkAZxRPVNxCaWJfE3iaOeaakxDydzGvAAbXgPpiJZAiXeIu9EREnq3amRDFoj6/F
TS3Y5ng93f8khLc1vG0ihntto13DCbSWQ3dunYHZIoH+BVWV5hXgmlw7OBpy50mU+OMdSd9lfsv9
8a/JpAzvm3r9kIs7edVgJ8Gyr0d5vM0M+gYMeUEAQICCqhGqcALusSwKzh3uxp8j7WwJCBCoLrAY
DlImJ0uIbYLQvskPg7s7ZOxIv/UcDc3ilJZp+hvOW2NQauH1cYsVp8kpwEe+1pDB/3ehqg4bASKz
quZFbPf5TtDlML4D9XVZVZxGXo0Tj6EVin+WWkJFPFJifGkzdgV2MH+FI65/ZAkHAz+ltIHDDn3B
AJ7xafqYh8B6dGwanq4bQW9paDBx9LEukL84QDpykUeSdDoxlYIqAnwCxKFATHfoF2p4qJbSNsuZ
VjqMJP8szhzggLq7lsegviRlgY1JqFSmwgE/MFLvpajNEw+bV2hprdzNeWy+DQbqKF/n9kOpg6mj
5oeLi9RugrKNkmNyR0B2XTTbP//LkcK9BTFlLLATL4LWWw1OvAywiBDwa9S8FW7V+re2w+DEKpIz
Ut4zWqO8aTqlQDODbLRQXiyhnl0EdS7xpd4y7VW6NpvzgAxkC0/L4nmW/DUpn57PyYNOvkyHGKtC
tno/kU9+jCrzXVTQmA4NhVayleo/146F5L3wrcXT4vDeNtvjHmpr8qivm4Sjp788SgX663+bJyDh
/MFtRmabc6Ei+HYOKXH6TBSZ4KWJm/kJmDyFUXKoPSwNmOuoGGWPJXLCJf/TwWmlSAaltBOzGcsW
7O1FcfYO4bQUk0lMpGRRUTSpGyh1EtUAOvrAUDaDkXdRNks3SroZEGS3fBOb7sg+En8nHVwCyctL
5xcdbwhbEmnfYbI1xQ1PC9zLPFlArEod9Ci5PPnirsG3NpGmB8eiOdyi9MtmpFU4MwqY50cUnJxi
gkk3qO3JHycJdlaTi9AMsBCbHeDcPNH9s+bdtDSdJYXyP3iQ9j8zTuQnzF9qT5pd5VGZ0xMi4OQu
UrgydhnTE+Ai1PnYzk+2/ZLKtUmT2loo/hwYb2h7VElcClAbSUk2+Aw1ZK+wut/28ELS61QThSci
Nm8vFeumqVX2SDiuBers1pVavsM3w4bZIBlD0gMl1dkH8Ji9jIJOH+fgpNxGVuCB7y0iJ+zW0KjV
Q5QSCab5jZFtiYg/MZ3wSzE5Fk0LGm7cQf9E+ysJp1TzuKoAbglgDsuHoer8AduXzQNvzy7a4xem
UtLXtiX325woEW6YHhFoQ3xj2nDUhPYvWGc2JY9qQGto14hwn0p3q3+1FYCgSTsRiAhbmnPKtREI
nJNmzCWUlMCaKGf07JAm0moajm6c5v6o3P8aVEty+tuTc65Od6192hcdEr4Ie82HHtf711xsYrWk
atd+JvevgpEW9KYXTLFjOcBcmSlBXpVMNhTZbMhxwnjBAvrWSXYf9pA64L19Z4Fn7YCvTqxk/PDs
Sgi/m/7DysHukTHCr9bzLKimxaW9zjAG3I3ZfBeS7Jw56me1fjNhkmNs8i5G18gRArDcFvDLcjis
J2IduYGWfO81i6o75nKgPJZuzUFMmtVqH4xpTeoFvOFxGPx1JEVFh+ZjjOrQafo9mpEJZ1h1Jgl+
552coK+RiZ1jGLBYxGcxT/2W+AZTsNo6ZbmkhaK+Je80Cs5X8dmbowZcstA5M1MvyIAYRag0PW4V
/sFTzjpEzlz2FRgOHhUCvtyUQ6mFiV0eVt7mw0Vd5G43N+I0Ul3aWZMRE9uH/zFWaZZLbSv7GnwE
8Z9nPKe++d/L88JosfHzgEmGhhnCb3DUQ6yyvAIe9UySOwo2nUsJWI2wS6Oay1QdfkXnn4VJfVF5
+++Ox537psztufgSKNzQ3p2ftCIL1HOFREj3+O5hxCkzlnD4tUSBq3TpMRadN1rBxREnxciHcueP
c96xE2k5oFaeVJZobti61rhRdoBQGDAFvFfaAPGHhspDhMJO9CIJVoKyX84EZZrPQrakBjgi9BD2
UYBs8vegSvfm2/CQkwk/vsub3zBsA0Odd6wdvmJlUJ+hu4aII9VINrzR41nRIgJUhzifIs7D2bVO
067ELxPlLh07qaI/vnT0ZCA4SmJjZtfgdvlVjCA1pFvMNcA1PeImfZO6K1y8xo+rdudWA3Sk0AC3
Sy/GLcywdn4P98TGZt4+2hPkGxJ2nnUNWZYIpwpX+1yzdA1jDZ3W62jGq4SWiNX4glxFCs+vNDWT
g+TsdzRszrM5uj4eYV2n070bpo0fdNu1lLb34eQxK31YEemC8Q/ffv4gD9O/abcz8Xc3gJR/5zNE
fGUOxQu/6jGXM8PW4VUHfSHEmwuWWw6UECshD/DGONvDJbtwNSfUnmygLGeYuyjCysHksjkJNSw8
PQkk5JTbqwg8YL5US7Pgnos2+NXJE4ayglh0wBZMvbNSeR5NG3uhtmlk3HOmO7NbCwh/H7dQqZPy
XUgjsyMrsrNg8astGqLJS7CzG4GFpXzExVt6RlubdaCUhDAzj8/U4dj9DZ8g2FYPlWVEFYUNwM8V
vimq7JJ7NBT3irJvlOOg/BbAQM5RfyH6XWEMNRjdbXan4TxVdtGHkKCTnj0R8HpoHGrHsnO1zALy
pKQfd3Jnij+GEEUFP3v+HYHzn0JK3w4WlGDbO96WSwBvNRoTDTl0DOPGwvMFdPvQcVmMn6jvMAKb
AFNgdkG0egsJA+sPFeZqkCHeimsxKEANWhjMuUvQbafssWo2xJtzpfnK9DkbCPX0hOCNyZWvpFcz
Tytvr0LYExYmj4DBrSAL3Azr9ZKHLc2SwVNXtyAgsdlOfR/KNjp2RdAOF+8nJT7mfuhjP9CQewNm
VolNUNWwy0ooWOfIfFYVoY1JbusvBOffampUNkEOJaP/BST66y63R5Rn0y43zgJ+u/TB/esOkiE8
Ie/LV/egkjVmXC32tPs1YCflE9xGN/hjf9aQHUcWP5mfnSoxGNP9vlogMsnkIbLQ+gcDf8jqf/Nc
OE3omLZQY48PISYRMgcp8h6JDcW+AH6N2Sat7Uegwp/yoW27sI5RJQJUxufrL5gCrvG+0/rYR5ET
tTqbapmG3rklRLxjfXwOwS1EKUJIcEUo67T4PWC4lx9Df+YhyhUsewQP23bxRdCtvaZIwZui9j2X
/cYLQyZUU7QmWTE5MS4tarA2Pzf6larSumiAdUG3az3ScFns6U8JaWfQwWvhOp7QAkLn4KeK7Sqf
A/OIsGLEDkpnBli75vVjzucH40w3LfLKi+1gZmQsDRK0rHesQu56WlvmT01LDigQup1aGtu5cntI
M+8XmaErybYaFSCYFDhcJYGqCDurSLz6d+is4tkJg8lht799cWZnltAmNEpQC26Mg2a7H0QEWv6b
S5u0mPBgcKG7tvSqBEbDeMOmNURdGggnWqk10zdjci07S/ojNxleRS5FUaOCNj6lP50hmcJB1jUg
8eLiexxyXVzgIfZhkADLhyYNFy1AaWRh2V99Sv9IhUgmJyS8NqO54eBtxLR6HhDuRryZY3fpWeig
0Sfi9dTxlw0Sj8Y9kYQvA0zGu2qGq+VOZH5cy4BFNRaI5yGP92Oe5rpUzKzvFDA0CpyrOXcX7U0B
UVLcr72Jem8r7RlsFyNQ6/Ic64rT+OoMQ1hhuBCwBVXFQglU4VIhVOyrcX0LoY7+kIbzqZOvf9bi
r/wzzFxIswoAKuJqgE9mgnp/jzNN+JLLACHnotxGyJ659kQBAFx14kcFgLF5hNhl/7/NI5nhW6BM
ilwVeIYP+j3Gyi5uQfbklPT3DL4hHp4CipARxuC10IIy4BH5mRzQibswHBv+A0sllOk5mOvVaJqK
CboxXegmIV0mUd0Vq1D+OWbhNiwWf36PCQXRcZwQWK7XuAcrFjQ2oInYRoUEEpQk2W1appsxoPRA
OTxYo6P1mIU1iot1XiG98DKcTa44m7LuV4bZFPKTuXfUJi4YsEMh7vAV4Mpm10d0FxjmLW0Mwd5r
Ci0KU5sz8UEDUXS5JuwO2KNK+mMeHPrrAzbg8P3JS2p42s9zpaT7CBNxKq52hGQxpk22i961R6C4
Y1oCnbzhVc7cateo8tiZYx25DKJQ1W02X0VgDCN1Qa4MwFhtNuRJ5ZF3RFpm4BjZMqTwIgOr28nv
OJrnx02wflYr/zo/PjKDce4uQMMA8sMHIv3MY/4VFjCXNdcxKO2HqWd9E6C0HMj2J5UEyL1iqrzw
TfXVb/bI4EveQbdwgwgAoTA9tnqOt5ac77ltMuONDUB6K+PPPubcaQjUwfvTj8/mkd5rICL6kOZo
FjIPyiOj62ACKM7RrmV+NtXZ+3pMHbzVRDSpvegAZ0pJax2mp/wNdC6UXiUPDU83pFE4vBAaw/FO
xMcx9VEjlyNg8Fh1lcfBnyEYB2FKoXjAebecUoAIryTKaS+Op8x5GsNzcC0KVkP9FdcnxzWQZGHi
426D1PiWB+XKYhqBxp6Q7ulSL/K5GOXsh3qEtx02PSETL9PL0OnoWIf08mgclJomqSwfkdpq2fZG
q27Nim2pJthlyxB2/qtCZ9IqDAztjktqGgraNLoVCggeDclBSZ2nNSdc1UBAyee7xQW7CGZ95okI
Dm0SnGEJhmscs2Q4wnoPVmrcYl37enDqk/AVbkUA5+RGWdujHklXCZJr9XiKMchvC8bRDLjZjOAP
8YUMXDcJ5SJe4cBJDSiVSb3YsZx60sVLHSGLhkI8plyyfMmlh9ihond5nw6jiVOunxmtqnSVkojc
NbWpBVTZHTqZONuMnFmWtFiG/ddcTBO6UWKsGO5Jjx2v382LfDKsEFW4tuvoG7PQ9VEqGPuNXhPd
OR1fdaQW+mdaTuaJ+glbK67Qrg21dvqhxtxhO+KCwydjCa7JkkqbkPJYcHjItFWRJm8IzU6YyHd0
dsNAiPCJ/yk2Zhm8dJde3Y0IClB4I40S/JcJLEf6jhzIAIZec8k5cEpu5SLu/bmQxX1J5pTmMyDa
RhDXsswhseAGyVNIp1NhOQaOsMFBYN9Kqd7o/z4P/OF6xMU48qW28efVEDPf4Y7gOqMHN/t3UfHu
yu+HC4wOgSXfaJkhYy0Wa84Z9nBkQbBGsCWLtPEUpDLAI+n1S9H9NFsGjd+oKs1ODjuQXxIgMgCo
9sTWvOVAnQlKn3/2Yatqk+q5pNYzH3YTAwYobCmTehq+Hh2KIl3j0RbWSS7rE3JCj5QN1lLFjtSk
cFUYdhBNRDmamTEoJhu2V6LTFlvjtTJjEsEQMsbc0KgeW5rjP4nEA0omLjjJhg1CjBv1BaoDuDG5
Y5rKtX4vaadWPObS7lWw9TAKweT5tFudieJO8ta0zmCO37X1UIl9N2P7vXOXRy14aTxPCN0fMEMR
V94Yre9S1InKQBxE2blsGPCxUMlfOXEKyRD4WnI/a0foSK0UiUgbjoc3CTxpdItTTJBbi+NNFFti
u2g8cRrXK9NYUId9Wh5KWUMXD+h63V1XyuhQyEmKAEW7b005d6XTVMQ+izW3Lg/QflapmNTLLvDY
LYftdZ5z70DfV7AxdF7X7EgBbwCdXF/u2Xgl8Wx33fgos09bJ34WLtH6TdgRUj1lsJxKUEioc0Ei
s7jL70tOju3WD4DcgNxyHd7VQmnVvowwtX7QLQc3TtKu/4r1CfqR6oGo+oz+6lqiWdtKh5C2tx4k
fqRexjTwYhYcCDry5+OsGwaTBmHKq9laY8HxcMYnYA/bgjNVPLj1mMLR3gMtHjF7lChyc7YuIoYv
lnx32OkxRnShf8Kd9uc4meZzV4ra8CltQJMv0fYLjQ5Mn/v3OWqkhM2ob8HVw3DNzF8gjLVEex5W
dZ8OCf2G1LOBVmmEcQ0+aMmYE5S/AGCO4/eHjDUzRvLmnVIXMzh8Iegv2FHLhsPMxO5u1rYjJhFC
S2IGLoiTdWzxxS/PdCrzMZSCPFE+QfsNDeEnZ6vlm06KvnICvd7i3xyO8Taiu4OvzMMDaG6UKvht
CEwINEXFxkcPeSHH51cAg6mMvCWAAPP2r7TNYSLrkTNCc+hNmu444scOPZhf7pgw48cfycYcOdMs
OtWYmVOvfW1GGS+yAId526NLVtdqFFs5WdCsnnL8QemUXFb6kYfNAZQ21Rn1W12ZD4d52W0xBwaL
HRuLXqtk9UMj6PUUWjZU54dzooEF3vXIRmvwe7qNK3n0Aw+YbvLZ6xJP0o/F55FdcSzoxY1KnaB1
nHAJegmYIvEf6PdJdcijNq3h/UZKoaVkb79AI3fpA0WG2d/6Tui6yEPEoG/RtLCNWnhK+C6bSX/F
rifieJ5QAnGCpjGudTDTMkpZ7AdPGf25QXq9IqUQoObxv/f2amcgTXT3BzO3951lXZPRZZCGrosi
zvG/5NgYbRkk4RUBtxNFmveNKY1MRKA0k3c6DIYh0mYQTwSXhod+arKsdNt76F/0Vtt0hFEFIKGp
Cs1UYbIVbOWRa42CoSNi/gmFn5JULP6GhKxZ6w24mJ8FddcpK6RXNPaObWxDPfld2ZKM9LLuXmAh
xR3nwSX4q9ctgt4/YVUFFlOyxU53BkE7mfI67RmzQY+rH6Hx3Amq0t8Lec88gKrhxREH0nRmWN7K
WZ7ZX9flNzcsWJIZh5ppxtcUMbPpNCsvZ4iRxGE/w3A1hPkOX1tfJeM75S/DiDPs8r23ZzKW02ep
z5TOkBGki09leied4wqy0ySkWQBoGDfa+vb/j6M43jexmWoX+3rX0qovWoBpuRFoMdQODz5mDWzj
N07RbO6dzbpW4fLEHwHjQ+TGHcyoK9M7xreoG5bslXtaddQ53SaSAuIgnd5lPus3VahMTrYP/HmA
bVhe2CFyZlUpedL1c/sXfPTnOPbNUeyh+tUhnPmOEZcyzDKYBxqrMPmmTt8XUlgBQeNBdlqdMzui
JLbnIKmBXO+p28hL7cvQi+KDjA+tgH/vF30nS02ep+/sAdr4qAL2EEu5Zb1ceR1lXSoxLQEnUDca
FZuo4QWB7G+JJZffR0KNqwTfITd6AtZD+HN/8rnkpkFm94bsfeqjzWfhM0wS0pDA+Gy6+n4aoO6d
DNmG8w82HG8PeFMUi6TQzFUOXkOtE88W05iGTXeccD9L2rmfqA1MNXIUgp+fXNpjpUrso4p60M1k
8DAIX5HgYXHWn5/CGKeXEV980YD3BVtmJf6PVz8NM5svcwobuBli248BBz/J4oFPaRR1K1MKaPuk
AFwDtK6nmUw8mTiLeLoe9RTuIQRTvZLetFotBp0g/dOxAGtcXKY/B9q2VFurDIOR1I40fLxIMJQd
tA/oEKYqBZpQbZaYgPEOSpeh/E1/3bu7t1vo/r8iRArXNvOcUJLiRbowjJaAH2iFsSrNfiTx1Exg
+7BIkKX0YgRTvEx2HrrpZ4bPwuLzheZxcbSyiK2sLg7oCPBZYWUkpFYxn8wighoTEuvPOPwPnU9U
32k/rG8s08YrlBuxe3aJqA9Y/Ze5z42wjn7PUVuKbGiWDrO4thKwmq2+DLejlEmvz7gIq0wFv+Bh
ilHUTHlR0dI5w3xRZ9CjiUDqyJLeuuARLRfYRQPk0XXfnOvRdWWtZiD7KDvZOJtaeyEeP+m+M7jE
MRx5j0zI0JpuNS4HOPhfppeiGduV842HPBh2fJPkrVMhMiw+SRRRwOME1tmJKAuri+cIBS/MVRg/
8DtA02msEtyWsWedMhaQM3HEfxINj5vTCktnN51AMLVFnhvqNc9prv7X6/TsjHFL0Ae1mvB4bY3o
f/VjW/iZZazCWaoQHOoIT2s5BlRZ9qMJxl+k7A1oy/vgHmhVbqfPoDUTZnkkc8J6x48KyCJyYQn0
BglqVdkLpgAlBupSGOh+F6rj0vt5RTVg824C/0ZZUSGaNYlD7wai5ZWHFB/+/LTB+SbHUwP0hO8O
TMwNw4C2QPlhs+9JH0xdFJVYQJJi8gevFrORTm24Oz35JTT3X/yjLwqdhmb7PTPEVaXabQRGRrRU
MXTY0kpwz3x5QjijNdk/pkyHxWBdHaLznxaYSdER64Rn4oRGRzbDEiLmL4rJAa/qA/AgFTF5a3qq
LDWJdLF6Ffm8/Z8uaNWPxvXJhAGkVprJuz5VOxrcN1y3foR6xf1H22P1rz96fez/QyOa3yE7UHIB
o+OUxfENC2UsloNEUmpxo4KNZrDhgEFUU2Z/Pe5Ql8B+azysRwWOlpUpft9LlgiRdZHv0Ad9er8P
66BUJfGp+FfUmYxtkGkUvGI4j5JN8+1vkjYUNZ4dYtL7aedvAnzKYSSSvh486uHQnc/W50w5qxeY
RPk2Dw7Mn/W+4Ao9QygyBJingbyzKKi87rmKvxD+ZQsngYuO3Y0H3l1v4+32liCck80yAg14uFX8
SYd4/zeDN7tt47xW5IxLqbQQtlBALa8XZ/aKARSKjmpMFC08ySw89k7iUazxblGOz23yytjNPR4g
KPqSaNatiNLV4o1CS3oUlmz9vLZseMdvzLicmbapMjXsDOWsBKgjvUJ/HEbJ4yX7bBZ/FVkbB5B2
xhL9+cFXhNaNgkK3dru9NzcAErcAq1p6QNUxTwuVePnb8Ilps/VZRFPappe7wzwczm9Ot4OUezby
XJ7ZAVAbWyGWc+xl3H9rpZINGJKO6vHWD3cPUGEzVmHnh/oawA+wmGNvFc/YudLxf4VyKc7iByYW
AkjwUKeqWIYRo8XQuhNcMsgkDB9eQDINy2EA4k4W5C80oowwFN/RY5sYnmTtipPtv72bMoEU29iI
MzJl0p9P/EyIwM/m+3JXu1ezQlwyPrz+hC/QHJJgRcg5BpnMkvh+Tk1QIBT/oNjYAMcyVx/ojxTM
/BuVICKd5k6RxHSnBmZ2bZmuww/84oes/lgq61Seqhp6UM49FUUK80792jTkZETZl1bSHCuxQMQO
Ph/phQ/C0LwcpkYlWAnTPM0TZ4SlIOnXVkWv30dVXIhoP3A2+Hj6Cy9SFIKkMKNjtG1UWcfkAyoy
FxAZpF5y1JR9JH7xMbT3Z2RyjtM2lKscTxlO9ms/p8TP6+T1jbMu8P1rBzmLKrX1m1g67qRWVmYz
eKfQFaImkr00lzrBR+CD7xhtBKezZsQUheva2oTUs5Pste9PpbbQhOSwq4vjEKIHgHqwghazXmO0
DejIIDE7P7Y1H8TY0ms2+2HPUDVyG9MVOM1L3v2CWGMVNs1V8Bxgji/8pRuwGo9hMXw4EZy4esZT
zJ1hc1WkQRHOQ6HRWPEw8wUdmiRhDdY9P+kM/s0mFfpO3GV/txAueXg0kIPqH9ZC3w+JkF2gU12c
EBgCpwr7fUPk8zX3n5xTmvVuHcTHjXVNwvKv8QsgQ6jcw5kfhkSqqgqweYMQCCbsBj125gauMyK/
fYVCwaY+CcC+fNgSrPqCtbBKYeBn7DQgFBFNf9WNMgGUfTrH9hp8exNOm21hFcRxzpPa5/J4RjYM
m98R2X4Ak02TbE2bAEjvftlzDtbrbhOd74GyOvR3gdbr2X3gzQubK/YGnR7dNd+3YvY8qoAKBV8y
u8hy/ktnBwwsZD25vFu113hpEKoPoDsi0Yt8MfrRFyNWHohHmrzhbfik1Kh42UFYLrZEUlZ813O0
76Wz2anCBanRqAplZUv83RQVU3wbQ3ZVONbLHOql1ftRm4qqxHT+LLa9UFebNTzmXS8ioJjZj5hV
XZA75S9x/2quu6oJBVxjdelABgJFGQwb6EbyChTzRJ9smm5qqWZBc+VeCfWnZnXYfAW+NIMRVzu2
cxYuamhHHK6Zj/TiRBjMac7gf8Au6V3HlxkE7EAOptI/IRcN+uug6gOT+FPAmcQf+jfaqw03n4eG
+ZtW8s9Mr4vT0WUPHt/xPOn76lD8hVl9ByIUY4UVsWsNHZQNhfDIBWSX1qSH9p4kb5PAU8p4sXDZ
IUaTDI1VvGCI73JtaARc7vUq1PArA/w+BQMLW7HA6rNC9Rc5/Pdr9ERN4BjZalymJEdmdMCMYL2i
q4OGIqUw/b0AcLotDC1HkE+RVNVOcZ2fOgEugk+CkvjOAFx2PWZWNrO2BbweHghmM/obZdOk45V9
jqd0xMrfc+/tgxagExBEHIlgQLnAZkO732Ymz4U0ihSSc0vOpDzc8wNQuyCwgZ0si3zck2VyqVA7
wVpJnJiiv+qGu6MAx/3pSxebG/Itu1BqoMx6avHwJgRzSQn3wwPvSCpbbHyXCIdesT5LXPnIt02N
pqzdml7k/ZhoYgsM6XGiVD05f4Td2KLNw4jtdk6EemhPJhKcrRFKNTtkunf8+F9vGun3f6asDkfP
i/QkG1naNNvuH3nRPXTSieAgoIPLg35NGV4iZx3PRD5F5CgVWQLOoeMAYVl3cdKI/7Jm7cQ+SqXT
sIyhs+44DKLjhFVzTkoXtKzMNd9UHq2lLoBReA1KXpSU6ACCaw/1iYQSfwTpi7HjWdtjDOgpUXnQ
dbgGUVKFUFX2HSGuLAkWhRUPGRIqf3zVZmEhVgTJrhiGw9XMDx6twmK/mR7V6tNNOncRYZL81CqT
dbR86eYI9JiDMD05C0HcnvWlfKM4krCmdCfiw209XCYsCJh5hyWLF1+sUitoylL9zwUepG4Ogzkl
jKnOfhYGTFI0S0N2QBT5PXgGjWcAqJlDA254qa1S4CUHKuC8C0BMT0XooUocs/4nb3HPT/2t7azz
TSgXQF+dGxyoMO47fVNZf3I8t5xdRMHvWCMiFFGxpNQNybXIsbhljI2W98ojN/ZoWEEQiWKZjNYI
ruuETMOKgmsjSw47IAGZ5TLbDuPROpZYKMTyqknfd7u2xFfiFUoduHUdlsDxPAgGKTNkmg8a1nHg
Xz31Epo4WeKth+x4c42FsRqm1tz/l6txWb1sC4BVAQzP0wTKU4lvouDUEDUwdq/hQzFQAoRmNBiO
IOIZTbCp/srS0DUMKnzQf9YwvbSS5wwsjyWERxKH1P9KwxIN7ZWoOcXHjK+0urnZTvDTaMxCSPf9
o3rbPfwylgTYGx25sUdtj6igGWyCLP3uiU0IRZsKz4blpDjyvWL9TG1d3MihXLs5MR8hxJmhp5+N
4QHzzX0E71iABx9f0aaag6BYZK1FULyXmorP2YZMrxkHdSZ5+tVnFYxNsZYEAuIVSU6YgODBoFaO
CTKjebGr/C7L4zWXArUX56h+Lm+pocwRtWkcSWPQJspD9fXKf7TMYtxeHXYt6jfoWdtOwbrlD5f6
Z07x3i0+RdIZYFmAFzgcf5wb8eD3Js8aOFiecHztc8DiqkiSi8z4jGVMQ+OmISHElch59EEeeAAc
PGHELo0pxnrliADFomdfBLmJpIVbNJ7Un3HmLzOro5SQFjRlZEoHhmI4R14t4xjwgWkLmtKFXTgW
Q3pZeGxrd4XIMO5n+aBxLmdt3pqhM6JznSBtiSLX5QJvJYMgj5YQOd4IUC+j0tua0SaozF7sh8rJ
2CfJyB5ayVejstaSVa+fOu6MH/gqY8cX4y+pyJkVepO5wzL2etGJLcUbAcS9wmOywe6uSzcx11FS
DCplm+WW7/NCZSHj+CLtnwVMn0yUybmXpSORMuKq2tH9iO63oDMNb7WXT1ujbhNt7w9lwXxo3Zbe
9YJtqy8vHgMlfGdqrD1x8dNNaXOPoK10Qhev9L5nsZKk4/ZenQxg6DVxA9n1/1eLbM2PclSFUDn8
aYg5VIdxgtxalXQmFFRb56pAHR9fKq1xeO8VNzpMfBnjOyAysFiXf7EqXG8nx6IWdpFLPPQrA92A
67p4TPXGVrcWAcqCVAuNUKdagq+AWvGSghHGlDJqnErZmsgr1b4oeFc0qBNoog5PQmtmg1T6y9kZ
Ql6OnqL/5hUkWDqXg11Ma+EzQNpE2Hb8eoHnJFxKwgXIYENOKhtdCIwT8BfkMM6InI3vP/7ghMxs
UH3u6o0PnR6yLasgoKlvI9ozUlA8iFmJJX8YnIZiFVP7GxNgznef4yCHTNj/iM7PX5bD9NY/82rE
BDMgA75H1VQZXsUCtpXwa26dnN6JPrIwg+fqSX6wEZh+8tmYntY+jqhTy2gTDASv/Pqcqp5WJhRK
L1vuyH07TpRA+z0TiA56nSo5XH3bhLPCVzmVBZ6YkzdBy2canRC+TE6RGdShhQ3rHYSMILPFf/d7
VvTXOczcohPwr4lZDR4vR9dMXH6dmKY/tikZxu/+PYW6Z5lu31nvHY079zBMozaYdEnlR6lYQw7U
Ay795TncX+msJ52OUhW9yUA8QRypFQxRWiRBN29Hxsy0D0QKdZ8oNDkaQL4CEon2MNRp+v8Tmn31
fH7R0AVFgJ1eXkAxhiWlc8+NCANql0U4Cz5D0FlRTlbSA8MNwZE/CPzAnY+KorqjQXtaaENsLA4g
LoPdmYNXl4fViHbKvWA/pDptTi8I7nPFQjwjjApWwzLEvK2s/XAyDQxaO6ouBpIrf7GufyxbIGYM
LccLnlzGJmPSMqd/7hF8jlsB7sbU2U+o/J3tVmr03u9B9BNINtBFBG26AHrtKKud92bBN0B7j7Dh
vxAHAiG29YOtnhmfSTMP6OiGF5sqnK+2po3XVAS5Ag07DJKKh+g22le6OhtQgIecn+mrT6JST+C5
lCB6M5sR5YgrznxO+R/OvieawwWHE7ouHxeJ4HXSHlfd2Ljew2PiHBSRDGoPaZKp4Gz+u0IK5wdB
GccHUoY3fjx/+XOJpGGrdsz2ovaAKDNConzJXg5mydSpnZfHkQ9RMkSBVwZGgr5QtmdNuTA+HFow
qyT6EQgIzlNJJlKDzRgxua/DkF3akj7BDuJsc4i7upjBgyPDGIxVTwKr9o0LHFqAGpQtgyOMZsGu
dWQFC8F1mSP5jHvOnPKXPZZfIz7Ru8+IZKGxZJytEVvPTLx811aCzYrrRh+bXOCtPzK00UrO1S0L
cSSWuZGEtPr7j8QAyzkyvS9tZkiUJf9NDBQW7/X1TsHQIDS5N+hWEqSnczRmaFftv3FQvy0v8454
ACpHMzEdHqVKicWqY3go/lcWBmg0p05QK2LnOr1h7soMKWHbv3JyROq2zbgRMsgKCTRrHLIp/ta+
xjbuF5azahp0CyMM+sDZiQeoM8xzTJk7AoDpteYzR9JJ1AFDfcqPavLI2yKLl5h4pkzPodcffCFs
Z9SXzvpfhvFrH1ABeOtCUGKYJVWdNDF9yoq9j4KroOL26iF4nvusVkKbFr8cP4DtfuivZ4xL+Tu9
Hm5uf9R64RH8AXxe02Sckc+qb3x4ebKqh6Yje5JacTOA56K3Mu32nM3mVEBX0M06XZ4kusc4NHuC
sDSZyYHN86OHBVw8iGnfEnhoiWasxTVsurpZV0VIwzI1oG8d0ccVt1/MOyTQl3yuCsAXyaZGJUzq
cfrCBmB2xTL3XcAzK9nEZacaduDpzs/+5kyV1MvkM5e5eJuau/X6EKKxCJI1s4DHLjRTWrzaoE/r
O8I560c1xcPNLRtH+UrUQyxWck6h8AMfZ3tMBXsULjkJDPvoiEni33wGQdLoMeUV5HW/3eOoceKY
hI29bcCtY1S5FY7J9CvJjD8jIa71i1Gl6g/twm3DkxI6i9A/V/leCXBt7fbsosoN1toDACjbHd+4
ZdPDclhV4UsGp/NFJwxq66nHk/W7KllM+axRr9xRmRgiwhC+nLmA3b3HOReozGVPm8my8irk2kfy
lQCTCgIklNBW3IBxgHEVWRRoFsOtYkRnRv5pV+kEPNG5ADWpzojBSTAfQflvLnbOS/25J3qufdMq
Xxdczvde3z//vG+JDUnyw88P3LymS0A2xFY+aCMC544Xrf7JxdoaLfl9QWUq6wvNZNPc2o8lh+R+
txtPSEBBpPpgL+2TSVGcRBoGLyJSjNM0nexmFUdDT4StwtYb9kxFU7CnObx2R0tZy4LrTOlNL9o3
Viudh+1YSTeVuZHxdbrMh0WlMYv6+Xm6wt8iVNBoBiDVnUbcIfemgULnY3ENsEvt11g3sfiCeT6N
OcDQ7pXvAY3GdZFIMqlPufGoiDpDg6rsvX373v8RDujCfJuwlRJ8zR7mNQeqX+dw6jJfu2h9aSqD
IK4H0nAWYWREZqUiqQIlckV4/6tYsTa4PAwe5XNbmsk3cG+FIyHRJHxLUHsQVnGa0x+IJmQ+xtLv
lJFlgajXHqHK1nGQoKxHQO5zOoQr2mLVqs+cE55YfYzD8bi5SnVq268qMHp0K6HrbLxwNPkvxu+S
CF/st2KXw5tAr0kp3BmkutWx5AHWpVSBHCp9iTvmOJfGZYID6lSCE9OzuJgu2cbgKYAf9FLXkUCy
hyXg2YwGNWxN9pXzC/O0eIgt2dGQJrh9QKY9CPlmAdaqywoEOkeHJ11mOUQBRd2zfJi6GgQJMhB6
1YlSJUOsbhuUoRxFfqr6UUApxlLjcaXMiDQDbh7TCdi8tqnBazK8BQ1NIe+x8/+bSiWZmcS9KTex
3aSU976az7hInsEQbd2w1XCO5k19LjHyIEvd7PdoJuY/qWDATJK7zqOslszLyznbUfWKu/pEVmQc
ir2FaytKCTAsmi+s4e3tGknsvohwkecwCrGtSkwi7iK3zuUTEhkdQuZTBVkbZHDEelErGKP2nJUN
GrMnUGOuo7hbmQcXdHgZ2F3BxFKa/SmE/K0H7BD0BdccZEOlnsboykAEVJbclf9vUluutQvS4hO+
5jdcTFcRdlZyshoLz8croprRzz3p/ig373kSvoeQ5lsD4AolBRaBYWfmd/O557axkgbYnk8wqQLI
s9jBhIues23cdRekJZfprL4XLiGp1k0DPSL7MUaPjnvHCgI5j+coT7lUgpvhcM6hgGMe4aAhyONy
UbjtDQT9AxEB79GneGW/b4LXyYwlGoQWB2mkJC0fgpzj9sc7H4SnVznmM0HlHyCv9jYUp8GjJYY6
T92AYQQfJruCrmSJoi94YuJ0tpK9XI6N8tI5NFUxjGGGFOaJ00eS9YQKMilQ7t5ero/jEPuvr7OU
TdllmnUZMEnHtx8kbDb5DtGqZipx+JCad2l0/uvD5cH+qt70S2A+lDuRilwPvdPc/Z+8HqEbPU+q
iKa26C8a1VQiM52mxq5W0vJiNiMiA4jQuaIEZ3lO5RFXL9mwTweGwtnBubny1REsKhMiUVftaxq7
yGGjR+9/YmLQnaItJuKjNvFZNjERO0fN1QLe1vi5LGwZjsd+r8jzw5ql0CCzJvSqtaTRn+KAZNM4
SLEH929F0D3+P51aJhdairepqOt0fJEotb6DygTWSnEFYoLUBqjPbLF51Q8szqYo/D7nA4jMiKBH
d4PXWMh3tjkQf8cXVEozzOZl043apRrNC8fatXUQuAcSqVzsJeTwfzkG+lE9kmaRjm30OIFztlmr
+w6olb2FB4LOrMIT607fUbZqvQkeC7s8Cww6767r5SpcldiLrnMnGE41kDGyiO2oOs0OFMUqw+Js
uaaCKDttGmIuU/mvFx/2k65f67itW21MxFIe2exzfa74yh9WoQv/SfqGuiFU4Qf2or3ZMxgoKLh/
5NIB5xgnVfZ2jTgTq/JytgPD5EeJrgX6ZTpjUufvDs/0ogY7TDHkokR3x6759SdmL2LtwWjxCbid
f0weVN1LwQ1BP4aGCY5m3Yi1Am2lYvDe/G4pcAO2PEEj+q080NmDTmrFEbS496gVeaApXGsCY6LL
chp9mEnbqQwraSfgS4t/rMmqjV1y1+GUbsRaJAyA+S+iJNqP3O6kYBA7razf34Df8XRI64K3YjBT
RFHjeFDB3q4zBF7YiAYMlJGw07h1NckQXGKBGM3PGxo5UEZH3YSxREyaYljoHnayfVfq3wF9b7ll
ITWFP5fwfCUiqRVEiAiqnNdvOMNlTIzR7HdS4jiAdsVuRG3pxJhlJ8RtJuPnJFuewynYUEAMH3A6
/+umBLhLKFJD7wsHXx/OcdLZLipSVho1j8xN0K0/s3v7OWqOzeg+8nV1M+igbVYS5zt/LTmUbXfm
rPMN4PpdezHXkrNnDHrEcDWqBxDonvd3nfAG3zqomjM/mDvo3z0C1qrzd73igN9yFE2CBsII57td
SBRD66XJ0aF4TYjxhubE+nSzfGZmXV/Jh3YIDVUjh9zGeAye/D6XlNTAmrR5niNlJ/39PwetmKPq
ueAd9iAfAUMmf6AkhloWDtlUd45SS/+9OJ86F/KKnAQgM3Ed9l+BjslZYRYpaPSRFcSyloZpW34Q
z+lOk4ZttqbQ2H18s6Oc6kHSQmEc5UwMSifZEHsdlTWYA59ItGqtC+ztUJLL5M6jcGYtwzQBcdzU
rC41ut3ZHMxwLFW4BMe1vZxxUViKEslTxkSJHm2pGxkkzDdZTPBxSoluS1YpLZ84wVJOsnTvQ9VE
lGo0yAUtMLfZ2p9aUvscwH/2GIKKYWii77Tf1w8cl3bm011XSsuv4TXqRZuOd6jEMGY3vrQ8W5fA
iHnnn8eTXSDCWcs9eyUEjPp/Q9GeXAH36u39OQJZYVBgJ5CdGc+YvjczOEt02V7yPFN4wV3Ep/pv
DHIV3sV5Y9/F0PiInK8EJZMrUXSjo9VlUHr0+0TXj+b2QVd6P3ZJUtT91UAcHJyMpzd0kC8TIpAx
w0UQwjDITZpnvWVEURURSqWEMvNSZnkLjZX2mFd7+BvsU/JbXevxHr29g441chbeWjiRzc+fCJ3A
Rj/TuQIFrM24e9NUhpEzQlWq8d136xGnnmPHZvqu1Hslv8FHqt13/W4tH/EHrhzL5w6vK9Vwc+2n
BJtmsxZFZontJ/EYBcQvm4DR754PD/IEwUvHwQ5xKo+pd9wZ1F7hrhAnsTDIfwZPDGXGhlT/gxey
2G9bDS0ks5yjEZl7W9K1bgdgKF3mfsLOlMowcrGJE3xlFJEJb/SabY56XVWFAorZeTeZhNs6Jgqr
gCcWrwzpu+07/Z6IL11rbYRzllYlX6TA2szPVxZUm8DHM9LAW76UR4Urr6gYAjS3nsG8/yxxcL9u
EDH/SrYA+5tvtBFBdgINSJnm7RZCsJF7kEXuyG32v6Sd+0mNDuxtoP+6k88ZRXh5zCR4nyqWXyah
eYL/CRHJjE64WPoVk0Ijmc/rquEAMWyOMAJdjHocvx5KdOIU0ZdMUywsoNTN50fVnjfCF5Q+slgh
E7wgFZAi4igRlkf+j1/4sWn63hgWCmTr5hsyDHuGD24+VuBFmg7Vn8YW84IoXYENODZBTaQWkNd9
bfipYW8z7VNH5FrKdm7Mq0bEe9oS1wWWkQ4aIwKwb6r49HcqLvkuhIdvf+LwR31I6vNgq5Bwc5DH
Y8p5MNPTce8S+l4VKzy+Gpzm9sFtPg5DUjmSUF/Au5GRKH59nvKfbCGVLDW5yThiihIJ4lRYQX2k
rXd3HLKnmjQwfuv4AFPDB56StsmPi8acQqTQVCIxY/UW1v7kKA+5iFJ4CUxXfvm6DRMySTYEmyj8
HC0j/bS3sV7bYKP6K85MIKg1RvbH9R/TszbCBgyHCohsoueo1MSE4qW21pbnN5KrjXwZJ67orDBS
5zq0bAdfkWI61aPCOhbGiH4dygSMbi7tQUsMLl3fPpwImSY8VPlVAqLBw6S3k4CKM5eSOreIL5Wv
1We9idKRI+bdPDbUeC12hm4lFzE5APX7uyIwq0izq9GDj//cWmw4LUYpRllC5WISYKMuElA7/PKS
KjJlczyDRPEeh+m7WbM/MZEFVfViG7zkO33YrSnm9CbQkQUkklviMSocQEdHmr0epqiFzQfXL+oE
sfvO0CJ30ug3mRzkqGprYG5yFOGYsGRzTUG0YRko3RG9MD/hoOJ8QkIF36UZEBbDJpumfvrXhJYz
OX9RNvuuLpuuwR2hnGxGI/hD2nwc2+OfT+Ch31ndIIjqNFBsbgT6nDHCqPcnvBHhEyZSI2DYjrZ/
r4xESKjZUVZSyaRHuCJaHLjyDA1mFzpvqZqJEvLtnAuwXjJs0s8y680eQvaUNJa1gCt8URr2QHIo
niP4FZVMWmOl4afcX/1eCYLZZKnCwWxo4sGmzacZBdsVQE5PHi6AOMcBFQn7KRLinxF7TvfikyRh
0/76mt2iFuUzi+PUCmqrY5kUqhVo1co7zX58ONkB0FIB2q2fUOgSnyQXhgI93yUIzDs+tZOn9t1H
oZRTkmYkV4iCiMwXe1rFFAjOnmnGBUiNboiPm1kQOWtPlYe89fwY3qUW6Lsw67WzV12rz3QFAE42
HQDlg3aV29iLM+K+vIABHQeSenMN2zccykLGm/kO1KyhX+7Bwjelj9BgReyViHpqK8eRwgnxeBBT
OH0p8aJA1/hypvirkGIkyplz1lf1IC/HOl9G7ZPDgNAMk6vda9lZ7ybHuMssTW48GixXJzZBWPoQ
oYkF/vWb5BSyBro46FdYpHzmbQWTOS4zWdc4dEmUzMhaLqiFiVHRxp6mFMFGzDz1n1A+vRpmbeJh
sPn+9PwV31nur7outMcC1wASfxNcecLoA3WaAunA7m21QrttbY+SYK2kZJTCmjJE+lZcZ3VHLtUV
XEOpBJu6k1jl2doP30CGwTNlbHzgFVuS56xXhnTq86PpEhG6CqvdWDj2YWoMltxu4oibzsy3pkFL
UAHBkuN6YEmKqGQrDYf+mYYeHQ48AF1UXuD+XuXTqJcc8+MM9qwTzgI/c2N+JHawUBp2ct0HjXTs
P2ZJbpUfZlGFayt67Q49ne/1jsh0gZ0WT29UWng0uKKELXGPK4se3WLxT5qkFeCOJnwBC6BC/1L6
X4fY+T3OX3uVeWHp2fZdIKEOmgVJoJVn7c/B8m7f49zYPlHSivVOBcJw6R8haHZj5fUq19HstHQZ
Guu3ykLOXn1zOOJ0T3aBxuv5y/oRkLEW8POlN/fPtLYavxJtAxC+Ll37yu0A+qzyHjtDgLbaQVtX
Gmviw6hpiS+uwdkJlIPu6s7RHaLFxm9b0ZNwruOZfcK6vlDhgAwGX2bQVM/m7IEbU4C7K9PgybdH
gR1bMOXIsK3v3UZ+e8q256WjfESa3mfNCsnxWwAU5UuzaRpi4YcC6h2vYYsiUWT0IGSeSc7yeqJv
DD13zJmRDMmQDaAsobG0ysA4DmKKsEDg1bO8BeoDvGUJomYm7mZZl9gwgSpCw0Ee0bcfeDcX7CUV
psWsQ3vgtdooIc4E9ce3PoKsqMIjUk/we8jraDco/WSm+5fIY9sAg5R331q0pt0YR8r59aX8R4Du
y2fYYiLni3P6OjO2c6rAF9LkFiEubxSZc7KMy1eNKHi4tXm62DQtXWPSFDnZP2VAHRzUFpLqcpVe
Y7nhcyRaw5WNgyDMQWVDIFbjmopSLoVY8elY2zyuW2kdDrE/FfRy43lkjvlQ+e6yaC1va5yopqgT
qXrHddbFiqPSikTe6rY7vG9AMuvKlSEZeudJPfggMEwS6NLnu0P15Qs7k4ls5c6dKbBV0k7KM/EQ
nkfzhTX5xwY7hCw4JYFak8lCyb4lFXwI1Fn1WjD1YstirUoMJnCVg57Ysevc9LnO7OK6k9KE/S7Y
U55LCrUhh9zPZUkqAiTas80+FV+DLArlHKZSyB5gqt22fZeiPJSDy6qFtHNRxfstil3BSFFadBnx
SDGlMBOkMqRQqZ8Aiv9MfTR5zoJjtvXgTahgPIzgLZz+YepSb+dee/ooMX973pLO3wA/cayTK/t5
3db11xYY1022EwWuAbyq7TlC5o+3MNu9GfllEq1LopGRKs3Gz+eFGyOycSQrwDNAwnPsXRdzFZ8O
hPpOzV0PLQBCI7a6yIIkgezjeh0QMtudDkgPJNqukbMdmKjYV6tMGM6YlJvSQnPr8iSMzJgxGFtP
MiLIO2dNpIjevv3GD6PygHDgS9BPm99jJ4M6KknF4Ba6rB/HMBpL8rjG/6mI4u/r0NIZA+cV0PHL
fJPSrXNIviIm429KTEMoWF2ujqOO231gcfbQ1gtmXRKa6+pgxrr6IIM30vuFZNjurTcDJZzEL9yx
VggCmwWtednqHxCJos3+IxYd/bLu/Ja7wdSnk7+NyAKw0a41VQBmU1q0yefuC98OCrGJS6zOUCQa
hp8xiG5X9fCIWuAXmuzJ4M3rSFa3SiADSTS9v1NiLPmSYFRwZb7hn0tsmgOXJ66YDBKi13a4fj9k
1/7uvgG+loLVhgErUllHTmYUEL1ADPBsK3R9RSOi6E9fS3WgVyY3ZbOdS6KgermUlgSLBRpO3/cM
A/zOOthaeaEtdDs8Q/m77jEyqeSjfAFic/h0iV4zI1QEDdrc6cvVmiWPp6L2NvpXdlXsnnNwv8kc
6twquLMxAfxzYGBIGupJISG2AGOwRzxjaqIcxAhgFvnM1D66pKP2eK5/abaxfLHUdyFlZsjAfDUK
aKODNadD8FW3rghOdw0aN6pNN8n1toz8lzx8SB859/CQvD0iPl7l8Zt9exChTAudSpuMgNhVGMqY
t2t30V9sn4gjO9aQue9/ZNAa22tbxllgUmKzgWsnbPxQgICum90gU10EZtgU+3Nr0OxYNEEpF6/L
9AhPci+kb5Fx/6eh8+UPinAOjUe8p7oojja8T/oqCsH7oHVzwD5yoBzd/8Z51/fcJioz7/migkzD
HoV6eJB4KfgysJbV4jcjeKuw4FgyTQVdLJsihDLVLtzeSUhaj5vFNilfIR6dSKfi7W4ytQfSehDB
EcUr92Id2A5ZtH0rol4/cCg9HMbJQcLLrA+8VJJ3z0yfkvziiD8CaAgwAgFSjLMRN4OLfgM4BmL3
iYVsE4cIGaHiXmWeWZQMuDamBrTxPXD+LI2RoaurW1/7dlBpOTKpR9WZw+XP4i13k3wTaolEYprm
DwhCeHC40+WOCzeSXKcWk9Tch29Y6jek5+GC4r08u/ZkKDjn8Xpu+7xmCzE/9JLOhSMZlnLpnozE
IPr9CsHYxrwlndN8S71kGV/5cbHxfHxoWyse4p5vdbl/SriLTR5V6mLb8WwKbEj+dsqVEpXcsgl2
Odxa5HsA6cX/Z39ZQJOaw4BYBlMQLXQ4B7kSh72qtQX1ljIL79nQA59gUlyaaQ3J4Bpa8LdHrjgj
FIi/H91PD6eZk6JZhGLb1LKl6Ex92niUiOUkWhN5C5TbpdAzk5PUxdMBsXFlUvaukoxN8t45wpYe
Ip0zQg4pPdodIEoPKLZKK93CZ0UyuobuR8fzDokkt2wGjnKnqB5zJH+ig84OQuaLi/Z9M2klqGLs
jHPbMTBw3iZbzh5tIo2iH5OVV7yNDZ73AbSjMG2IZep6inE7OGSsq/dqAfjFF/bpJa7/AAuLH63D
UORZdwxjeZGoH4nAek0qWl3k4lJh4VfmOW0cNDeegb6V8jhtetkMfC88kUBGDNZrXCfrrazkhIrk
JifIwBQ4rVPey8d6WgMpRj08Tfk/DFem7T88yOECWsdNjZmbny7KEMdI/p6GzLSG6N5f9SXeZ0uH
iENhxqR5GJ1QEW3iPHmqTFTv8G7EWTsoHakbXNd4Hb+coXcTOhYRULKoX1m3ex6a3eMuJc1PvKpq
7uz3FoQxI4avapoOpKdQDF3sz6gX6r+tCrG8VfJ/RmsxyguYcY28RwBljvAD/heCPKs7CMKGRhoB
pfxN+UM6QWQJ4pcHTKA2IRmRpW4NQl7qdAyipEdZbLhsDLYqLAqTo1Nk/Sz8mDRKfNoRLbglhVsC
rmd/HOo7H9f06LWU8j/4e5iHBuSL/czQw3ji3SZnmWLqEoDYEUNWVwz5X7eMBien1YERppYjXXZf
9RxV7FCuWXDb4uyLBxhPgZvCNwyFpsIskw6NRpjiLhJYlqYy2ymKIXhFglw7jqlrEqnM60+riz4N
MZJQJ9/cSkbiCmx2ExmCyhcSNpLwTA4llMyPXLzm23CxkWhA478zVYcL1HCqQW6APcrP9r3EPKlL
7tId2yISgHEJXZIOLU5hLG2kR0puvDau8TCzhI4baiN/I5uub7lzC4P1Nv/tuVBFjYjv56oilMh3
QjxGZOHmLRpP7hiolY0JhNN/yU8a5804K1fxub9gzNtDwwGdoKJkuBePUR7kK11//H2QyV6h4j8L
bErsy2+1fMPsJ3ZidXbscIKcklnYZNOjtTlPygOmK0aMPNm6KMCWRgdjc9yhfZWeTknzgmHcQIyW
INeDkhuPKwg+Wo/coKlIBgkrAWeBJMmjzKYE1NGTGq93asQtXFAQyGYjb++ZPFHRr77MNONfPT8X
5JF8vnbYaFATqvvH3Ocg6qlYTVmZIUsOdqdX5sUB7uIaREFBV3hRI5CHVUnyDGMg8DLtxvXkCXXG
9pO0+k0YiidxSginr9ym/IgAuzC+A69yVfk9JUqLZV1CrE0TrO3JjqBSvbbHSvYO8OiNapzB8fhc
WtkINitDGf6G/0ojc87Emsqp0h/nECab4xT9BB8O8a6rqq68N7EHYG0ibaLr08xWRcm5a/cpF9kM
62gJKETfGbCxyZK89x3phlHWzERX7vFmkRBHCmUrP366aPubkNNJ2f05EqEFhJuOb1Ev9VEdf6Uf
fx/g67oPg6ldlJO+lKzImplW3P0ztMEOYCFNElafVxWeHJ2NyGC9DD+Ecj0oZfwv3t9PYHVQJTff
zep9FUmSUgOUrwHRMY16+Yk94kFhCu6/ZEuG7isyAjqpoYwIyChegl2FF3/rPJL8+YlzLTriPJN5
qYsP5/iyvYDGxHOZpz93AKD78jDSn4lScVyAkU81L6z/ue8zzgAEIuTL61LVCNG+yiEfCBP0t1eu
qKu0k+MKWaQmBrrTOxmJ+ZFaGldBcvnO66GrZ5qYQ/P9ds7UUHe7o+PWk4OGiAegVJyPSN087jW7
Xlb/NLHh/w/L/OEO2zFXoXYBmvz3bD5+o1y36NSl0cYJQAvfn2EAzwOyL0+QzcO8H6FA8vU3+CZl
umbMsuGF03/GHe+5cwiMc17r1RXXWpUzTYT1JS+s9n3CQtYhFco/UW7PMrGR0ohYaaXbrp+wiy1c
UI1Cb0woJIUyHRIK4wVF1TKhit/KfwwAol0IdenctEX7fGWr/xJdccJPAsyf9DYRFbuXazdJgZSD
pvYhiN1McexDwdsgyXH1wgxQy4LSlVsrweZ22bkE5Xubvo6tzTFd8faPR4nWLWVAAKJOTHbZHT1d
4YBJg9nBj26XMLyIIYSdj+1EDFqXHRyYGnctdAnsn90OnUfTA1ZY4Fj9nl0qN9j2wNfRloyarG+U
xDR/I+mq/RPG2coErBytXFKsahhyBtpJjAg17lO3GB3/gND/oCF1TLfKOWxIsWofj10SuD29YCJO
W1AvN4U9jbdEGGNpLQaOT457MpaWbuAOKLoLj8aNh9QAxkKM/yd08aji4K/jkknBDnbBqAcBSE7l
JdsqS/pE+RVXp1PEV1rLKiUHv4X8yxgF7Zh4QfgWxcq8Hdlc779hPn6Q+X35jeQpEXZUJiazWfpN
lXaX6ovDd5ZrBVyEgZbqdTu+qSxX9TlPU0BKnRaibbtbYo414beimCme7Rbes/N/S/oWLVsaW2Kp
+gmz6NSZtIE3sKpBJTqt+D2jSJk5WeSgLyRygX3iWz7Yb84qV65WhE5yGAqyVKzsJN9aSMjsnvAs
NWj5+foDEs/gng/uqXgUyS+XDqmugPTx9HV06NWliLPn3kHNDFD8ospqmJ2k8telepZAhUdsL0Ow
4ldUT8vnGzzuYtC0LBsedqnqEPrR19UYSBVd7plo4mcPwd8ScNrueui0UuykTQnyqmTabmM65WH0
XOKaDReyAIzZwa9DxvbzK4pQ92EXjV+N0ZKLZBawwT8hJ2DVev55FcsZJ49KM59hXdwZGXKDGlPV
y7oflTSNe8MGfQrkikoNB/DLMR7mOOkXhzQ/rErztaa06PD+cx6T9Q3utviBQ3802wz8bCpXT4sw
KZcupCcJZfItIg1Vx0JWChL5SyZgQTHDfxJWDK6waXLKIUwfaSAI/Il+hzAZ+BAXKQDKDPzttwNo
SPg93CsLCCYL/D21whKJfYWd14XLXwfWTb2CAvL0JwVlMLZuBMmv4sVwWz7VM0ugm0a1DgAOQuJn
H79HZBWrjHERTZRjOrEYeX+fuQkVWdljn9X9OAVmY3spr3YKykHvV/u4/T/F1bW9Iq421Qhs1CVX
9AFOfWhirEBaW0LaXvdfQ/mespE7bY28PG3vPPwGeqOL5qfRvRGYzwSWYq9qWY86GA6BD7uqr13I
8TxmNN/5vQuAHqs6db7jl+5qAYaNnDO1RwVjce3rEUl5DnRoalGnHdiO/VFEf3oY4SIfzP2oVBOb
J4dTNN4RMX+RF3FEgNHFwCGbJjcVL0+ujF9l+xB5py5c8MunYeM/22DOTCTJNijILvOKYUI2J83/
AJYgOmR/+8VmRkZAvGhSXamhMvg3FDrQdAHBqR/T1E0GqeMCeQ9Sb2jyq4kC8QcIcRf514m6YZ/F
CBtbWaGzsXcfLi6Scp/CRZQaYoZ8aJ6kaeGBVtf7J5MOrooAQVcg7QX96wtbQjllxpL4I4ylKoQe
igdckwEVAIF4CcDKNvNOJBkTpN562hpn468HhLeeAHJle9wGo9FunrrBSowlI30hj188t0V/RUQ9
MtQQCFycEDBOO6/3NSyQH/wIgVcjUa84AAlJNBINb53ZI+0oYcQjwJxfepjFKIRqtArhV//7cGcq
Ao6sD5Z7OqLWUtJh5xBDm5EWH2THZbERlAagj1nms9JVWsV9ugCmEKWQ4a4npGxJIT7PIQF+ZqwS
q2sDa0N+M+XZQ9fRu8U4GSEwb0PEtNujLVS0FLUTiMaNKrBFOcQatuaK4eip1+3LQV1vUkIuanUu
jLWjv9HJgDB3canSWRgyLWIWahr6cDwmhlJsOW7oLcMhNO3/O6UBtbiNK51pc39bOssr2GaMvZWT
nM0W5JzkxtSg7dg4PpJ7LdqIN95fzP7JKvvFVSxZ6uFWFayeRWuhSPbN2jYDH/psFcSDw8A93mIw
g2yJgC+uHzb5j4EhAy68W+3+ZyvTMDP7UKaMlbJ1kjTRVPq1N7UrRXGJnuuAcvRq/SNd88Vw6bo6
opksK8XR0DhYubz+W/cAxyJy+gopoUJVIv267jHF3C1u5hggfyoKAisLych1A/Cs2+r5aVgWFRVr
nXGYg688yzoIOYZynOXW8vSpY6XXJX9Zaae27AO0TZy2aQqu+AiC1L4DQB9UFsHFIBfXUrx86Tf5
YHpLiLP2JPKc1/wfnKrlqJuUJy0wT/uk6wc7E4aYYuEVrigIzrreFIONg2M6YJwsXGpWTOcd1c+g
1nR4f1ONBGe6AZrJahpLjmh/xW5yepp+DNcqgA6IKdKfRJDhQ7uKVSdRLECtngEmT8iGfZdcTcLA
xc9y04BWIpIxPXMUQNtpzRjKVslGylE6YHMPkNphqu/gc6No2alcv9hWvAzqROECRb5NvgNVUraV
xBKsEKOwWRLLXznRI3SUjHGfDDhy7mtUoZt8v0dGxdzeX6GuK+j+BBzkaneqU3DaTWoNyybPhnh3
f0VVdI4U7GdQ0lpep0GHaESrZL7DUA8NPs6WBrQQ/Wy6GdTAV4jEQXPDhOFCjVVtBDGt8Sp9Bi0+
v301okZ4312J/U2/8qpgW/iiBU4Qtbv/dMGCQ6xyRu4yE/XrxlWDHVOeNgAD4THXxiX4t0DBqP4+
oLgQ0N1Pwh4/nBNHz5Nn3IQjqObuqYRu6EkLRqifOZEHyaGTIriIl8RNrWKcwZ0bhVZhFh9Ca70Q
b6tv83qYk3y13nzIYTLyCakCoNRn2apbMFNgdHG9Z5pdihcAFOFI8VsPOxSNfNxK7vCHj3NivIqk
qc9LlQQLu2dkn/AqqgqBK9tpDA5i/v7eZJ38E+Ms9MQtPiT6nNbudq5MI8JVxUwgjrT3q/8mDYEJ
3G79tkeX8ZEl5XDgWkMkbpSo9DhKgmNioEdZhNKqYRjEm0M1kvT+yHoXbzjbGBvhhu+KVXr3V+mw
COxScex2ZLertormda4hWcM7wE21w9Dm8fs98qWs+USrnJTfS5DB2TiAKX4fOpRQJ8mrMVAbtxfK
xhBHI72Rh+H+5tFd95SSDPJ3+To7OWvTbAErjTOjshBqTQtfLIs0X5j0t9S5tuK7zfcuIl0atRL4
ia0KZkTh8s8JyBTQ8ziejf7tE8rWK3weMEiJllhgLgKDmUyTpW3LEWTylzWBR5RunOTN0/rKN+Mx
TOJtrgOYj+MsyaAyOh50cd9OIMwF/bWAGy5+RQdmePc0ZolKFOlmr26LIFbMqlqeR8LAKNT3fAA8
vAquHauP+lZwEp9jURGLty+jbeE4RHdaWbFuLrj4TpI5U2faHoxz7q1rzlOfEXYmuvM4tTbMHjqX
al1jvYJMcXAMIjPSTbYX7cK+Y0OfWIDRjQtE/BtMuyrJFFXVYCm8uxfu+/mgH6WsWimSDoI7fWpN
mO6PoL99F7sBj2LvXRX4FUJI7DwGWhTvse2siYKG2tqRu9M/9DfvZIFLUf1ovfh7gGb4to/GuTAq
NzXlaG3BBOOe0mUtA2uo3QPiJBy3a6dnj0WC4SYCROH+As+hDMzam2vDZOBWUt1gjLzEfOBxASKQ
mCIFUCT2VXl6D35ndqYtp7KcoDadbKedBbHnlzDHaHHUyIEZ+/9B/Waq4JhG7TEWjYWBdhGj3rtH
V5Jp2voh0gzIVRR9b/WFAtQkgE4B6fh/jB3tcVZGMGTc49gBH6Vd1wiJ+xJcjc77llWbc+pC1JFw
bGwr3brRPzdwHzmA25f5WIP9QPPfzZaviL34S4yS6QKD+8y7lTGZhuVrl+r+j+5J4e7c/XsifXY4
uHLCEIyENxjOWTlu3RE+klfLA9Lbm/eo9s4Q/fj3gZytuiH7peJN/TzQUE37UxYaTa2K+Yzmv/PO
YDMZF9HFZ3RnxzCo233EeYm+VYQ3ethLaC4/wX1S8mXo5P80s5MudphX+KXZIjhGqowtYUfvGwYr
7STt0yFvrcuc+XUv5+yKckYxgJzbfESZvPsEKi/DezBKGSG6DS1Jpn2DWMU7w0g0FeYF4mNLztAG
WFDEuWl43VFinT1aFBX15eG3pi2u/u2BsQitSNNM3/V03m/D05iohFWrSwsMTBsAqGMmrhn5psXO
ZGwwMTyyC1h8FB36m90L4B1wGQIYOYSd0SzUHbF3jUcKg4hM7pJRiRGK/CxmYa8w5O17OCgXesmi
Xuj6Jjv4of/xLlSVLZRl+G6ACxj5i0r2Lb8/xmT/4cJg2vRJEdSkGCoKAKfiF6Tr4S8ZpSmQkRRs
nWl6f/D3gq90NloMa3PZSoZLw5pCGsdVv0t9qd6fuLZSE4P1gOHLkdTpX/lTMV0mo57LPQP1RneW
H2A8ltkHvMyNmfBGK3EXh900xrWSX2m3OonSPQfkQF9T71IYjBNFhrrKWosRrheq2SgDL6gzPHRW
G/6n18x5YXKCIUrQ2f8klWdhgmLLhVjf2njr+W0dp7hJ5y32m1vb2hSmoZmOUgWlGXWe3lhviz0t
yP8FpAPmOEiMhI8YOIuoeajHcXdMdjV5xNshuWMS5azIyVo6NaDPlNSEDxMXsWmyy+hnA/cewuea
1rLr0wMi3pNhOhNaUZVrF137oCwSKbM+Z+uPCE6S/UsXKfaM8PnCFkAw4BoxlKy3jzMZu9soij2n
v2jZlMEHhL760bCoCKtod3zdgn7nhwM+HRMdigyLkat27kohGpokIFrwBmABg0EfCvwkOs5KWjHP
IZ6k1Mffg2JeNdXQ8ei/2TedJ6viS39dPha+S8qhCbnQuG+f2zRGC+eVQgFj+3BAA0BuixS1l/Ye
0OsojmeTefIiH0suDfZraoS1MxZugxZopDnhX1iX3eWUnG9hsJj35x9cZ2kvgnaSPbprpt0UvUjD
S7bctfkj7VXx8Cfi22LUBRo0HGLuGLPhuhJqybL7iZjVxOU6rokqTIhVmNLQRjydPpw+xwZVNlwX
4MSXzt3eW18v7icQaUWDb98y0BUj/U7ZEwcFkx+mhTKoG0gQERv2tPVVoEQmYLsddPafXJ6ANI7W
2HFgpQHA9QrCnU5r2bm9cyt1mb6jXfM8/kQSIOXMa1oM7/e11sRpyOviYotsCr23U+a+IFhrmjN0
OSkkCjZwUu2nK8nY6iAgMMDTqjsKTiz3+sHtqPzcduYda5iAMnorG4h7u3uj8V070rVbJUDtTRad
t3CAoS66gpIxRlxlEXu68mVacPAixBGQLf14Gcjk7FIfaYNEDW499nDryytVVvQDoSzQqSGi0A8L
anTqbUlfOJdxXWLGyp7Ln9IU8cwop4SRRAinoKn9NNfChjuDTUJzhyERnaaATRB2OhMt59bvV3D3
pz3qg6lswSgnJGh/wTEH1AAX7izVGJaPhpFA2CtXew52NNk+4XGXtB7i4Sj/Utq6JSSJuP6HT0G3
/ssdn8/LS0wFnwTtjIc/jTiFXZN7yOIArX/i57/LQEIrkbgAC0tt/Nd4iiz6AabJXHjU6Z7CoPB7
Ly/xLyzz6wnzcJdpzMVjBogCVQxLnNvWnEZy6CwJGVVVce03IHxtQEVaT/DTdlak193shR9mcp9T
i13rE9UTYqS29O0SUul5/VJT3xQetRS2v8i9ZygLlZShlxkHysc88h5vOFlgR2Mxf70ss+4435ug
iek3unxEExGpICe4OXRhw1f3Phl90CbeJfEgpyi/G5a5T8gDMc7/KnxB955u+5YgH1z54NT2zyQ2
MCwuzioSmIi9szTjU2CyL9VNcaTuX1PPrj/NKiszbVXNFL7DDBU7S9EQDvNgUxZc8iTEA6tHHlVw
qZw2fTk2QBN31UPEzpc4KMz8OyhDVxV0eaURI1laj85UP99X1rBz0KDarqOLHiKtM3e5OBr8+Aja
ZmQlZqy1LmApMVqgBjgvUW3O9KwTi7UmbnY3XGwXUqKTBmeoPVIUqKQXasG80FnL/Di+4zW+qe2B
nZW/kYj0YvGR2dNQMLJPcREaQEJjCHJWRh4/0ff79otEIR63uh7j0WfW2iMeJF5CbBaELLuaXbHa
0VOsWVrvAue/sHoUE5OIoF5n3ZS46EQpIBkUydjxd8oR9T+x+aH+T/3wsJsuOC1lgPYzd7pX45h8
RXOXJrsWU668qP/WrsHuNGnIKlbJE1hN2b9kS77CD+/E6sFaLQQPVYE2n2gP20qQKDRXdT45GdgA
DlY9hzB+PEJuFl+ZedTabolAYda8y0ZEDON0/Y7F3/SRB8LTNqQa1nmAc72RFu5hh7JOZ5bWyA/X
ZPx4jE2LMbl2zmkg/09F79X14U504QbQYpv7WvHzrzbITyj1fa06r9kSpTz7V/tJ/6tfFDnohL+i
UqiMucoqWt8EoNvCQfyrCK0WkQJ8VLTagnaSyAg48va+oR3RgUVscA4Oe99v8nUW1wt+JIDUrN38
o66Q3l6UTES3ulvW8cyBHL+IH6e3NPNLdSoGuBAtUyWX2F1EBCniLVYtF2ZWM/oZfSUIgh+1X4t1
GBWj/54YOTBeuthAv1O5gu1yYHtlT/MNh5LSBYiE/t7DKpYu9PP4NFKfu85iKbb/BYz5Q250gM74
NyhJ0N9xTmODyQamr9FqV+DLt5P/tXa3ZquBUuwDPlCKY1/e/HOsqDq3RM/I2qVbJZtfUN/jPB7X
DNQ6RsJWjEE7L1hEFbRVlW7RBDE6G+cyP7VoAO00NZwKIIxSZoX9HaI7U9p1El3B1YW5Xo6XEdnh
C1ytAc8wsM9qY6n/d5icjiB0i9HyNS0dmxLWZHURmAxjI/f4KCbj+1JKeb/cnCF/TmfeFApx+aOE
dM4vPf3DDWetdBzxdt70y2tkChAMYmy+gqhQSQcsIUekaR0c4UhvggYucMVOq9OvZ+r/K20z6wC7
fnp2Sb4Qv2FKOK7UBlIxGF4l9rL4Umh0XEXNqEaOPpBmT07RQZT+VzbzBNWta2IFCqmrkF7Jljz9
xuVKJuYnzyE6JzNdNjf9uzxTj/QZLSREwLa0LeZ7qyJ8Ij5fcRhxvVWqK3X5CnLVVf9D5nsZTC7N
MQzrHClsytc6XBrjQVl4lnAulxsbibxJzZmO65TaWH+HCjtAxtfAFd7dUSqagM+HpTfEZ/alZeBE
l03MT8K9rCO7C7F8AkWJiPZOFimFhlBhvWygeh+eeG1oTKWOZ5O9HY/n8zqjqckYQ0RZMKKAcZYM
PLJptQYlsZ4YARa4IVpgP/Wm5CpfU0m4F+VIRh/WM2UjRZ2RCFcQ2GumZzs4oOS0Ts987B+bKeus
koeA80+//rPiptMNP8MpGjby9VjlYaZhyp6mqj6nMq/DrVyWmAine+2gN/YZTDp16gKiGkvdtc4K
qxefvcMcZPJRgt5+x/HS+NZQ7/Nb0ozapQR+6Sld84e9Ku0YvhuKWNVi9rXKjO35hwj2G40VDwoF
mRsYP01BqUds/zzGHwcXjWTwNcCHriqwpXR492W5v6tBwN4XMGn2boQGU23sNqE9n7YQ4y5idRpB
qY6yfrGUXkTtNVTqyoZjNbfP58mYu1yAQNxZnDi5hR6s7JO6yL3yFjw9IlIoPMvNzgdbPL7XxYKN
+95RxoYnQD15z6Z4odH/5SoyJGyfOl4Y/5Y9pBArOoMw7uuwuRarNIXmuH2PJejydSwtEkcaIWIV
rTFdP/bgSZJekqcLnX0z7VNehYdqq48jkCuPZ0lyGGJl4m6VoXGXNydcCl5uwMWhWwSUIoitYrg2
TouB/IK1TMtveVaAuhYncwCf/OdyHl1PUnuYe3D8knI/7J5o+IMszPgLAp9tksjAcCQmGjLU5/9F
jh3arDz6ef5sgsIYNicOeTGOvGwRIVA43Eu/6EadwY1j99tI9058xLRSJ/9TDhZwUs1BUWuA/+cZ
p48oPqB+AFP3b+Saz3P4PoYvzDy65PrSMb0bxvRuJtfB5aXeBhkhVCJEM6gkGWOoia3rzVGxPwZf
MvrYlXnKOY6ujH46hLLQUPgt+Pn90WTu5k9GACTncGSU8fnNrhog8lpPPwskaYP2Y5ghkhNKARfI
Ll7dVFEKXYJkhwf0SFGJe54Hq8LCk8524PfsRi1lTyqR5W2ap3xnnuVJM7EDni7Lb5AFwmn4n1xR
i6cz47pmbL6QvwB+FzCuzYvgoQEMhxiXfSHjhVKkksB1fWrPKXE9v94qgySWqRV1VTRwhuXlilzo
J/QDNur2vZTaCBh4AUxBB8zCYzka+9dDXAPi385JRXcTDdbyCkcIeSYrSah5zPCn58f18Z2lRTld
iso2BhKqgJNDn/u4ImEnzr4GCALQ6DnVywXkuf6geBD/N1hCsZdTGh/PqlTXKpJtrhBxWXaN9+MN
Io5Vug+irolHi9jENkqVioO3F6BfRem2wTaP3fCCqGXGWny4MWOTWm2Vqs9hDNhNScxKZ6HbnXP/
fQE3Udqgokx/b6sIo3urNwlOZTHRqEMTr4oDPN1JKH+dO2E2P2tFaPeXvhZwEePSS3DVlUZIUJrF
ePkDpBVRGkcqptAgLrbTHTEm0Lq3GtriA9HT/GlTzRMG1EMQvVrH2U1TkgbPbwIFKB/xl/oIW3XE
xl2qPR36QEPqzmPAvklENx01EFhhSJag0Lq4/iVQPDJbZ5ofed0L6b/nwH36bn5F7yhIrV+StvOp
SPtGJHP5wNvgeE/5v4X0KyWCC6XDOltQsRHYjfoirY3yaLkF5y4jA5fYRglaXF96VWgKWT/pj3HT
H6CCN3A4EsNdlHB2h0yM0+kGi5vvUJIGjUY0dp0GzT0264gEnE0kqo/bC9Xzm3SGNTX1emq87aCD
A/2wz7cVecj4S65MEViIuDsmIJeitCKP1JJrmpwN+4uwK9i79iSZxWVOB/GPJCkZZl3pYqD0WrO0
eLopBogIVD4DWDTlLmL7LlsNQfBGcr3D2MAIjmefCYR3aZC5Tx6SN9by84NmymNlTfqYG4l5Qunu
nvhzoHrF+Vjx2RpaiCHmjz3ZlYQIFF9vO2IEPpUc+tu0CN04cWTvspRkYJFDWGx+9bQEpYFWYlMj
JKuazVkOjdwjqTPMhcJSR/s/RjopaU2KOzal1xwJzveRmjJM5IrTGQwiEdXtiOldkPMLB7rT0jIp
jz9fB4pWwiIugPmv+LF9HCMVgc2ijlpIws0iA0JeqFQMi7PKLbx2Ofbf0mazfJRd61fz2+hX8dt0
4aj0PpeHC2lrOJbax5TYScQPpoorBccJNl0OHmpbhEabsmOQggi37JzPuYuUkdUi9GJBZVss7kEV
fPkO7aOjomrK/2y/GQKOIOuU0S6oV2I326JLgULvJZaR7m7tq2OX2pNv3NMV5sA0Y9zlSMYNWOU0
3Pvcek0bH+AnWe+KHpln2XEv2OYVWLoBaawD2da/vIJYGzjaqQ1XY+X34XSwx+2Xap6ExHz93P/b
NGMa9fjnx2CJn+PbMYmrZ6mA4HBx1lgkfeETiD3x19clJsYtFdkh/iWkMZo8PgOHwanhhHOvaVTO
OH/arvbZjrFlCbEPW4fSNNf68sA+DyM2khNwd3xrFxYKet+REewJ9Nlq8AnPtdR+/yvL/+5m1KPT
umrNxjNocQnUoDBp5sLRaAnvVHs0KyH0OwzNGn07MO2Wjjah1pR7BCKj+FGJl5jFtEFkcd2AixtX
sYCcBviYeSohdTJVhwvr61ITOqRtaWsYvl/GmC8fprwx4PbhQh3egrJSObNxdhqYk9/pwrC3eI9X
Xh02LQCCUoB52rNG0NW5sJJ+ug9EfKGTYPoEQujfNL1zFeIg9t0QNXop5Y+YuCZUCu99qozPL3f+
1ANyXl+RK1PDkCx0vbc1RRHX9fXR5t9sP2dTHrmxJlThX5IPOv2iXtVJ4c6kpF6BWvDykBnFLA9x
axg5Jm5R3DE34PbEb10pouCEysk7lZ9sPXKs80q+1MoAp8rE6t9fTg4KstbQr78NeAYDYXbUjuBx
pYa3vW8Egi6uhO9WCTKLBgqTSOixoNKIHLJphCio2/8xbmOI/mzoZAKVbGtYqypsIJa+xY2fdiCc
T5W6Kf5+YC2qJfZAZK+2ka2+h7NUGE35//+qH5vqPSXXGc3st1/ZkLHxGXslOdXiB136r/GJejYM
3j/qeeDIs69RB+TEazELWFKIZZ382Kf2FIV2m/FfvbYFIw+dHoh7oKRV/sEavISKYrpOAd7u2/TJ
9Ykh3jtKc3iM+vfcJzFKAh7ry0HhS1gc/1yHBJxhth4VqSE8VW4GkKWkHY1KbMR7CH/2qiuzF0OZ
NKJ1ctvGtRGRrfEy8iEvQMHBM2Z8gdYhH6eTCisFe1hsruDfozPwCUdDQr9TY+ofU3Svjz9paEPP
9YDOFesV22HWzpoetvX72q5NKw9r2VuCx0HmqHYSIGV1q9ix23wGxQSWCNgEF+1CUQqsLsISSnpQ
bMbyJIDqqEHODASkB4d5KRpXBpOP90wxAvXzu0Ia5hX+cQYCvh4MmXAaISck2lcUxDA+Q2sV17xk
s7ANT5w9Co+Cpm+EQ8n2K1oXMzow2OSk3ZcfilYjH/SFVNobl/397g6CMW6iJpMXijeKDAY60Wiv
hJPw6rTZ10hBHgtF3z3OTPB8Ujv3+8+4oBhRR0q9sWY1GkD0qG/kLI3rFGgGe5DxxCLn+FSNHsM9
pFAU2xHD64iSPVou/eF4gK6zqgnKFoTBQu7/khzPvZ6qfJ/rw252rQy8AB6Oq4hj7dw0Rljj9BkO
lJNICMoDrBp6CrzpmNSVbG1SfiLhCZrcWYardWfwgpsSJJ0GpLmrlCHV9Q2QNTesaX/m1XOHmw+P
8E3zkI0gYizTO31bVU7gmWv6Wymx7u7EnTJLw+qOtLRid1EYdZqMoWpkr4U+L9YtV9uOhXII+lO0
LZeilWR6Mm9tsxBWHRAdVy0hV04y7XC2dD+9eYQ8mWMOaVsh7mII1rwxPm6okWGyhXeV0ME/IyHY
qNmpW4v+0lhP/tqOABc9g2n/SD1YULX8WOwle1Fpp8rGz4C9usWdIToBX0Qzzv6n6DfVPFh4rlpK
sE+5kgo6eIrNpwemVPj6rgejMOkhh166VE9osKilZEFaeIAwcH8JaYI7PxBEImvg2BZ6PGiADMTd
YNFzfmXlfMxtocVZsUfAyDKzIWD/m8LeaxcyGbO5SeIdHg6Do15Uhu/jh4cXvrh6pUHUWR5r8Yva
I2ADs0MO2MdelzqMn6ZgC+izg2ppjSDH7vTiwDKGjMBXPSzKa0sI1+PylRJAH6mBkNAZB9q23hsn
HFkkPOD3HILHEBXq1imJ0U/jwm43J5iaep9craZAnHk7iNH+hsvLFSDAJDajWjseZkmRRHMSTiPG
oCCftM0Jp46WclLcx5Rb/ihmhc+AV4z01fYrHLhGIfZO4DNrYgXM5OD0qsG86KKaO1AV6yPR1kYS
gWo7l32S6NaqMHblPKzpmONOtaqnaxIBW7aa+PIB8fATWYy4CVjuORSem9RPLOeGoiJmLwFWvDOW
bUFRz91snDD9bGSUqQjJehuczRdVabvRvemRFHRfj8HgGazbNNk2vI9QtP+Ay3TUJHv5BZvyoZvN
JBaTE3lsKAuDm62BXFY615sQQELs/Co5tkSoauekjTZVUG9bKMb2zHofMSp7ZjgqcTfFA05ENVnw
lDdA2jW8vzl45Wuj7xfuV8Bh9o9ykYNcU3iBwQ2SlxgnPmOQ++n4FOdudiSeHIDfEu1V2SrwNQPX
gsCdrUY5der+UPYdHk4YEWlKGe4GPMkfU5A7mK1NHUCqlkvpdEGnWjJETMhrBdc3W3ndpt2FhB3M
uPzlRemmr4ijiQkxFCeGl+KHGmEDggW6iaNfdF1JYpR67zdPWHLyFC7FxvGlfer8PtWvlJXgt5Yr
nhecaCUo+TNhcMOdxM9iDbeNnbsfj9VZpAG0NOJ/+npD5RNuaATyZlZ3L3ophwbOdbq7N9GL9ShJ
MIR4lGisXYSEsvzAmtVVM82ao+KGOiLwlHXEP5W+mIBpAzpkZKvy7l7ARpVmJwVETy4udHMf+Nn0
VLOGDj5GZ0PZ6yXpHIJaGdBfWmdwQVMm7Bgci8qdSmxBBrrW4CM15DvV/ZIPx6yxCsKq3+lgADyi
hz16r4oeIgXoE9Jt46bO9Sja2OOezISUU4LMQNyJbS0f735/7PXTFq62ugsJSUTpQT5meJtwUXWf
oEYXRAdzUz/fqV6SnERPFK6M9God1UDRM+7OcRoRbQKWXubowFJ0p4TPn1kHR/A9vlX8SpUW8jaB
B1XMSQASAL+q+kA3prfTIjFaBn4u1HULe/1wOs55pofMaAKE7Gpz04gT1o7sym/4BHVbxsQuVuz8
U6ikQ3PImJIFLMVJsXAIQEf7dDNgl/cHLCQspNteKXVsuIaaf9pxNulHCJgSC8+1JkCq/dB27EcR
gp+usENfBJamPmY5FiD8T/r6Uj0TsmdX4dTc9KUcwocXAFtmnbXbV+331dSVT1aCwkcOucEhcZzJ
QquqK5r7qPjhw0hmtbyxibFWvyu6FDFgO87CdwkotMeOlDMbSZijMfRDcHOEN4tHG539ZkFCtUnU
kPrZdokri66QwA+EF+IpK7waDHcvURfPLlJhvL2mCtCacxjgcVDZkjWb8supTgj9eclxOHJvTXtT
FL3TAGO3d7aLSgIv5GOKCtPhMA6IrFNG1Zg4ndZLIW7SNoFpPT+BHh2QdEnNEXgL2PkcDgLpmylE
JQfWq2l9j6LEgbVAyKkYIItYykfLMxJWGFI1fr9wt0NxZFk9tQgwnIurCCdRQh6xBLA4A9oRJymJ
1P501e5sgCTdtj4AWHY9M3miWngRPTUH27XMyvvrArZXX8FhjowAg9OoUWjwlY3ioMxy0b2xl9Tr
KVIO+RuMN3hFsOqfcjmYj+r2C6vsSUWclOFeKq1SV0p4byq5qZ6S2p3rkywybDn6G1p1OP8l3XSF
G3PGvglClVPY4NF3dAX9sossyuM3glsMSXw0K0KSmoGr7+iJzfFFjoMKxxVChsG2J8qS9/GaI4SN
VJ8vvk9gq3R0rx/27tqja1onZZ1e6bPIO9Vmwl2derREld7qF/Doo2bL9/MIwkBV0nEMdECPB+uw
umJTfemSSFLxvKzAD3vN/009sVKAh4OTlAnev9Vff7P7/0gzfb1SutWRA55XvG6TiLKimBji4Emt
aUaThDwjyeQZZ5ku23POC0D0Q7l8KvmhFQ6U41uTK0th+QCzB20U4KLm4B5laMfq1RYr7SVf8eyC
x+vfNZ7QmiZjd8lBEHRbMasETNZ/5d6Loal04fgweSuhuR9xadJDYZaKeXFgzRxOUjPEcAVYp3gV
seau2xGIw1YwsVa7swojj5rXFKpIjmuXsHayMzUEra2pSTAmcc0weKKN3OaH/O8g3M/ZKYu+CohT
0n+RQgw/9N5Fp4zr6vrrSbhBOFfbOVvxNi2/Oh9DBRHTtcu3l4Ibp3qMQI+cpnMYxnDY0DFlhzLM
rUY+wWSsAkXsJfOHRyqdC8qWx9eC2ZJlbeIOmBOBA7JjEgUHeqMk4zPdH1mVgo+KhDZTndJVgkYY
KtiAXDYqsuaC1qXly2SKiR8XuuYd4dOrE9vIC9domHRxjSVdgLVKjB3uIwIC/4nNiNXKkdZy2Fai
Y80AK/dTp1ax+aGUEfCT780QSrXjRmdBI/+u1n4N6Gv0hKP4Ul8JS4OYj3H5XIdcq82JX7NhwdJH
P1V6J/SSdS1BxxlXeGdyfG0ZbydTwYp+JYwBRmKLCSUT6WscsFM8qGMhWjZ3NoaPZiLtvRMcIIKH
SynL+hcdCK44wSOiOrVaVz5nx6TjMxvruNwtck/n5yqa0VkNhOIA5/3kEdj/TpjNMu/q5i1nZnWx
AHxw+qxZtWvvjvchq6Q6SolnAGNe0w1/6jt76vQhIlcVz5yIa3X1cGf1qRPlOxCb8eKxGf6UmrdD
OWIYzb/muqk+kzmLfKklyNIVofNsRC0uQrilzJ1tQKgPwUDXkd4U/5GbhNOwwNxzHPmVje0tYCTO
u3aIUR3CT2GmGYlTEs4h5iGvsarHJ+wV+Zav9wSZHqJwljuYwd9piQ0LiqozXGnpjS55cDwB+CUn
3nuZWgz86KLTZHhZySoU7wkiIfbSt5fFVd5lj3/eftIFRn8gjTJEQeG7xHlOaNBym2YbizGR4r9v
NLXjSFTglx4PjR3u1wDm47cVAUGZHaPIVEkaNJ9Yl93wJzhOgAs29o2Q+iL9c8CiN5Ev/e3k+Qzz
7HGXFf1OGAVkaIfrFVS36anaUcMLsoMhzWBktrAxEkAnFOszXmF49lU994xd9eP55EOcYZ3zf9LW
vo0iydq+2yxZcBrXK7GcSunGaxn3nUUeAJIsHGEy3XWZNd0/9aGrr3XNx5/9YBVYXoqNTt+848f/
xQpT51Bd5V9Bz9GS6WqfNgB8O3qb74lpLcH3P38JrI0nK2GmmXnzmUpsCkH57mFRFc5AfDIUGPkG
gyqB6rnvBYgJe3ubFqE5FfTuuogw1mp7sAvzTwACvdU7rNiKvmWdoPoP11OGYF7hjsTlhR+66YYL
g7b9ttE+LfbszzkLUISuJVrWeGFgG9XvSZy2nqqa1JG3JR//H4dIu2xFfWVC/YrDTXVeSF8svwEq
r5bFOZUs1lUeUiDRz1jRkqvsZyykhC3hIvWo+Bxb/OY3u4J25FKhlH9CPxplNDXtCKrzPLGpUWBl
nwww2TlDjb301znBXq2TmcuQ5T4bHywEpkf04NOB2mI4hj5aN1k18CT1W7Bf4vyGbAvAHU90cTTI
4dNYdNmUIPHPkQ90IqGdRLo+CZNZG81WH6N5oU0htrJuLC54YV1iZM7Ceqdp7wxy92gSaFtQHmpD
Sqk1HV3Md5i4d5icr2Nx961LvNXXwSToKKxTzng4Rqvi6xx37bM0a3y2kcMH9UIGpDSin1TRI2Lk
MiPqipJUqc/mOLYK4waTBuGRs6z798NBFmbV04NXuycCpzGCdz1rWZ22vmyZRYvNPBegieDufj6h
xpzw6BldtbUJVoUNn8met2J9vRkJzWtdiwodEO5yr8p98RQ09VdsfG+rwXBt+2C7e/wXZvptFzY5
nTK/vBS0qTQO5eJ5ySzmvu7jAFQFwL6EXGA8rWPD38Z1nhZ31iZlaiZxruDozvxb2cEjrE45f73O
omxjQ/iunFK3jaLLPZqjeSFSqbtt2H8Bk/s7+yszd2Kmq1Or9X5wxbEBtO+SNmZyvPhTJ1fBRuS/
IB23RMNAz9j0JOkrufnrGWyJHloYcc6pvZz8OqYrBkVXuchJEu5UST4IvR1UhcGNsNd0Pzaq6rTY
lW3L1u5HzanygOZo2KgzlaY/HW1L2SbQLMnLMS2IZoVIFf6wbkKTeJop8rleWsXkcKG7Epzh3/ZE
Hj4JumB6cOzD1/t0HpN2Ccf+UEd7Ag3Zt2UP/3zx9BQwgcJXH+zAdjovHiFUYK1HlYaAYQoReE5N
z28j1oltTkBIgeMEkNxr9CGCFez+H2ur0zuCg6Jk0LlP1wEIxIohsmS25KEXdp6ktRp8ieqjiOiQ
mEsIS8M0cBFbwIhyZLHiAG5U0epJmmVlSOI/xznvAFQN/keO3kkzST1LPnJ/T1oT2mxOa+Glbvi4
kKSFPKNZlIAKH5c92pLXWTRH8ycLNcPOacgG4s64kx/doZdQ5Xkptd9601AlF6kY1/y+3HGKp3rm
zuSAKs/Y26txB/qppw39SVZHLvXlOS/1UKDsyOS9WDFzDSfnRbHhve8IEbnWwDKJv8HWI3mvc1io
oDl2GjXRi5xASBNKlYhW6ENFAsYZEImipR8wLe1MLe2DXUUhFmfNXI8ci3MG1TsRPArLAymhjlxe
F6h6lpEOhowftGTI+b2+SCA6QZRD273JKXFXONKqruDPssXrgM/3xFWG3a5+0rEPv8FTVzXwqdNC
HxEo7sks2bm5noVZCPhYu+9ZimKrP/wKwPQKLpIOPXf8Ip0Np6bPwi1QrWi96Ac5dgxDCAZWpDxA
iczkKao1mqzG8ZF7lj8gYsltw63WReygyYYH9riPWAHd7ITAwQ8+wDI+3nYxqvZBdeLVefcwkKf8
cHU/IBXrkxIvl1mk/maxv5SGoQHy50QBWiDPSL+bmA07bZ6EIj3SIibxXqNRio990AYAEtHUx6nh
nlYH7fuWvr+D36R5pvYfIhntMwl+b0Q6PByK/WQXfhE+gxOzMw6Te8FxZ+hX6p3+aN2qO7ufG9yH
YABqzSsmgBTA8NoVF7lsGk/lgUdFH93zIAqXu3Va46qwXpmAVgrpU+0uBldnVrI4El4jUBwhHgNI
oWX1peMYRANcXroO/0Wh35eUV/Qk4chTEIxcZzRosz+YtF3tUPw9ucr3tYKeuMATbsKk5eRBwz9z
jSXCETIino9WT8+H65+DGW5wbJSpP0egs39YfHLrlNhpPRZ22juyqQD2VuHIw4QGYn+SxoYc1vxG
Yep/UrqNsfIi3eP1jVj9WPsd18aGFxOmRVFwQ4rMHdR1yuLDXnrBWP0jCHMCbDLBFEcD1OKIu0Er
dxI8cXueINPzZdALwIMFNtf4WqCVhf1dsPNDORTGoNGDhl0KdGSKbMuAQOzn+djPOY6cLYc3czwI
nhnRb71KoS9CiawYxDzMEhNgbGFRvEnkd7reNOwFay9zYvOqTodKmzzRw7c7PrceATdn+qb2QsXd
wQpbPAXpNhakmN9GI4rWNp8Or01xATXddPteWpQavu4+FmFlDpidD0rIk/VvdxzPY581gxb7GePR
5Ekg6NW8KYJOyuhat75iGsD4Too6hil7U4k+7cR63a1awEm2zlnJSh2Cv85SsBewMjtJp25v7Fx1
YVnKZjIn3ns0e/MZ+GxA6MdNZKhvZdO4SZDDD9ZSSQegxch0a7em4BxcWKm7f8A9fdHGgyrsb9zv
Yj0VRQKHHnFWQywG773TXm8d3xz0mzeVSjkKcvnSrmJtY8waYZoiRLjqaGnHC3CYdSd89n0coK8R
rjmQxvm2io7vveRuQ/Ov9+LLC523Pi7cRUwgEBOuIt4mHCuQsrlG4PMBWFy48DStav5rVMDOPABT
hW4Unlkb2oYQCAay04+mqKCo/Jld0yK/R3LxwHzUIJjoxilNGcP2CZgjW/8nGQ0IDak9wJpc4qOV
W2JzUWMtpPAIzu9QOlIxedaaD65WEydXSLlxgWayX06Xb6vdpVJDfeRw5KbAmoAwvRtZfeAKhFKg
Vp1jwlH4vU7M5Uhd3MIp2Hngi33OAJX9LHoN/uOOlHFumtmBTaO7dWvalkX1IWCSQxHfXG8mEtTG
7KP0YxDD4CweTg+RwtBZRjvbep5/fIHa/w7bED0J/bZ8j4mR7ATYDZER2uJd6pB6rhFrldbOIZER
Cd8gSJAETJh1n4XG94YIX/YWOO8nLnfz11OvyR2n4tcRbOYfQ7VExArf6rW4JQdwdVm/mV1V9bMP
fLJeb0KRqdOKiwRRtN+ZFYyFY29hcJTyZ/1RzUacsTolsYcPG/bvY/ny2WsChNNS3mp4+J0BuiCY
yLYeZH+ht9Xbwo6TOwCVL7pMgIyUnzVOHogI1X2bdMAr9GiQFztjLT5WWhIXdnqHR0aM23r30fer
dHIRa3c39+/kCcZx+rHmzlFJqEli+ZcsZ6M3H83IdsWaMl6e7EVyHx2o0/PCdLTKSD0TlZCAeMZF
DAshhIYlME6aBwK2Kf5l/8/tViVP5yIX/0ndxX3NklV2FMRivpfiLFTFd2hOMOddRcCvC2NcJ819
Y4ODhjBtztXeWebVW8Fg0DjH3Njawu9oTooXjl1yfpGXJTzSe32icI3Pr6Bdu/XsXOyUE29FZJac
ik5DHKqeqxlKqELhG75CFMlFSlSdlZEoYIcPVSW2hPNMN83PIb4AB/Zys8Ypno+ENTr51OiB2bsi
ya2o4M4WjI53mcy4XMF+BPTYbOEIehxUb2V5tFyR8fkptm2mpmWfuSz+k6bq1T3jKCgBZA5zRwL1
EQt471oxuI46Kcj27vctoqcDbVfKOxcShrOTVWDpqhC/p2f+4m5cw+Pd6m8qrOUqD4iswVBcgeYu
X580sO0+J52VOryl5ZQm6O9LoZSiXYqQBvuDMP/HxsxmCd/7MniE8giSKv2Fr15DiqQe7OSEqwMk
qPLaMj9KPQcSCFiegHdGYliATuUl241QndUHIGUIBdSYw9lCvTSl9wF/3i9mET0fvvxeNbgqLR3D
LNoeGifXzGp+9SARKukIGBOjKQjGqZZSJV9yGvJAwChyPftf+9Z59yFUFTWtSP3Zdfxv/JjsKEEj
0dEDNrRIPNXVHNAaN7RpUzfDcTnVZZ/+kFRw0qbtWGkDf/XT8A6O2OZQfoY1LEv4g8ENZUvOz1S0
JrqH9hGIMnLDNcvFMSxEE7CVDuwgrKrDROulQwa5ojHwHwBMfYqLTrpw15skkw4wq3KtvC9FXvio
WVdUP4MvHS0520/y6+IMzo8JWeZB/0cQGhzhpL1BnumwZJpC/PObjPaaywj3gw2QZof5hmcbtEG1
ommKq7VDunZMnwU9IjE+VcTmSEAmFvu+RZACqkPJkKKDAwEvzCpZ3MBHFc/XeSrK5ipFwnQoxWmZ
MX/N4aTNY5BZ3gH4Dox+LhkvooNsJrq2kG9G8KiaFgAAAClZfEOkmYALyI0jFmsKOxWTOHsSCmME
zIfW/cEiLDhXGpscxwDVncqgeotH1b6d3mmHLefUIxXuNlBel6xHbRAi7LqRIW0PgSB+oKYLVA6r
85MCkccxfYxr4zRh8lpyDCJJT0KAJY0MdkUp75866lyrDBnN4vciYBBedYdX2JlgR0UZ0hoMaTbE
Pg5WUZ0ScdZ2msGTzz6jbjeXUt4KsqUbypSoGUNbodKGeqXKiKNdMUtx0T/H1YWWdC8NpXsZINA/
ucXxpEBpBdn3x0iWs1M+qh8eilRpCZYdxShkNjRdJ3FOkevJELY3ikSNhyNhcmdCpuCR7FZJSHrj
400ZQyhxiSVMXj1LlhawSVQjntuktdlQCVbOzuMRaIP2SQFIjLMMVmPFVV2e6sb7XyrMrjwsJeVg
g9EUCl7/ytv+RjJRGuSL3AGatkVE4q5ObgssfFfgv6+ue+3a0ai3mR5Wx5054Fp31IF8CBBIn1WD
b5UXozCAhzEG7evOfi9rNfS6jAelNJm0cI39r7G7UTT3Q0+DGo6mIbeVciIWtoeQLAEhe+Om0bmr
zVAyornGrsdD4HlOI+IxWLnNFuQPX8GPGKvsNrsV8WTHNsr21eCxr7HKEfSikmm7lMbfVW3PjJUq
EHY1pfhZLyPR+GHnNEwPHAwD7uOLLvJMNr96Fe+pKux4MJIyvRhV8oS+9XKuXlhvevKqobl+vhsP
GPbPwLJSSYZM0A+CoRZSCKVE7NYloWy/Yzba3wiUD53ZUhxlUPIj7mfa+8u0V9LcvuGCx1+qT38B
k+SsKml+Vl3V8O62kXGsrYjwNoRW5hWdtTJLKeZ9FE7jrLoJuUtRQzxPC3q96d1lo1gbBR35hThN
Z/qBa+281j+EECluc2My4H4A45JNWj/zHvlHj8OiLs4eNvxAkGnS0wpYj0zquC0uUE7ull9Odlwi
Z0AnS/1eKar58BU8hAvgEzyCXdHIEiZsh/cuxlgjSkYJwmdwpswVGCZ12pVMe/kjU6NvSpuxA6dV
l8BjW1zB7sfCL7h8VVUfjhXb+etpCgH3bfEp9nR1Sy1k9TLB/EchtlaYkqzcL4hh4LE5bsihBpiG
ywjV0qaTKEkRX9kFkhh49DNb5K5ktGQvxYbwi01CO2NUqFyh6bgXncj6cejmChM+tnd56CUBr6v9
m8N3NTTR+Dig+d6j7NgdJtxuJ+l39u/r0ZhZPxoseJJ1ImwfrTL7i7UDrgy7paP2c1R8yuJgn73i
+7LLfdiQQHP0a47xryzB1txzZkagJxhGW1xwJ19a4NbyqmHNOWHeLhyxypUl5nm1sVyV+JC9pEUj
+tSp37hyanIIIUpUo6i9pGDiTy+26nLnyC3K9Yd9l4OHWYoa7UXL6Pvm5Uv/8buWX7ssupBPd9j2
A8Gxt3h3y+Ctdc871VS6w3WMbkPwiUcMj7sTf0OXqb3xrhW2FWvRWodN6lD4TL9xGlLKwrqHLlnx
mxbuc2/As2J0NAKsFOiwuZVz7VZ/ke001anH9gDNDwcBZEGswe5Q4ot5sVTfREuLrQRpRYIWg7av
7x/BD08UHDoNSYxf1D4VPIgCmnka4nSJKFlrCDaOhozRMF7J3HKFt3R20lKmCxpNXuccCTgPY4EG
eE9FOwJYx9QGhPVY4/HYvDR6iJkfr0HKXbFUjCH7d2wwtPp45f4npOJdIwPEP4yMDrB0OCJb8Ash
yGFBhRKkL8hGIjgT08UY1FuYkbYpVYZAF8pVioQ6A0ooxAr2WxX3G059MvZajAK4YBq9tvnzM4pg
NFKhRuhXd0AmicYxCh1SJf1yqMdZYqQOyEQyB79alJeMLPsnbSkkHnGbDzU0tTs3KcNVCqUpbNTa
1fZDdLAXkV68Ay0n+keyV4BbpHbSxgLesqLlDUr7BGdyitV4Eg4zZ/nMcP12cQLxxBlOIIxWIme7
7YN0UrPN3R4iy/YIzXzrtPAwu+NqW6J6ufWMuUKcDv/IXJXpaD1yeOXywner6PMHscHxwdRJhwJx
uo09sb/GNGwu4dAg+6gm12L5xfGEN1EKoEdQRav+i1JI9XI5xvUSlriWY7voBbd7Aq+pQAEDXwn2
9Qc7RUYzbClf0NhYAySpK5g9KFCeKsHO3MkWSO427Pa5NvtegstM3jIj3Zoh4YNWzJEs0r7KXw0I
hDW01HJCAwFHG6QrqyAo95SRAHWg8d0KIoXkTNEgAqA+KZGnNlx2nF6JsVrxKZpRpfamIW6KT3Ah
bzGMihHXFXDoRkEDH1mHim13B9OPdCO403IKf5DqQXUucQZkevaEHdLSLKc1RJ3ukU0StTtrbz2g
ko8QOJ1D3Dk7kOKLZehUkctQqKPWSlk2H8HZefMndGiyrcQmy+dqARVyWxPjQ9beg5Gp+L9ZP/q/
H0YocXdOlOEFCgb94GplDV6+ZGQA3ngIl1YhodFx1GDBsZAWfui7Vh3bsKYVjnimiTP2ekKDAbDq
+yZPEKj5AFoLE/ewOcdq4Fr2YEQVJgJCHK70p7Uwiwp/re3iGVuBl305ve40loCITVzECyJ207Bt
SHNHl+erl3pef/XH6EjDVEmOf/InLtulsaxUlqQSZm1VhRLWtkQ6zNZ50KkphrHuHWczKr/jhkra
JW5Ehuv0n9vrfEuJpqsi396EFA1E1tYU4lUq0c7K99sneVuwWSJzCPtZZVG5xmGE25ijdwa9FW8z
FAUt/r1qpj3SsRiSrOTxWGlr8AiVR0LI8GdjgIDHbdNBfWmOtsmetnv+sv5PglO7U3G7ljlGvCBq
Ub30SxfrEC2aBE5/7p64YI1njOYKEr+klbAXzxd+DCUbNjyLMQ6yXZn+x9punrwXtxYuoune9fYL
JGlQgTEVaGTWiTO0lJb8RBqPNxWUR4oVnL9MubJQcyvk9scSVDVA2Q9IxNhW+ZOQO2HncrbBn0kf
w60HSfOxp0WJGvK0oWElaC/srgmmNUmKKvIVBvL9xas8poygmrc5r0CuAijY4MO4Y1SFapOyaKce
ivbNijrAEHRUp5VndESdaSxAD6QEqvvDnde/HbHLfQvBVPrhyH8fCS/nSyG07rNeUlMm5xIOOZlH
7Fz1zrECgtD3cnr+Jd+uzLPf8XUNqyyIjjODAQMhmIhWLp6C+e2a9d24+MmdhRVCB1L7XtS/6dcK
6Ya/tbj+De4VmLik/4knC5V9U5QBjQGhxKYVpJz0aavvVlANe24ajAro/HI789tPqRu18lF8C1wv
5OqZ+jXWZnDsleJedzWdG+iqTkolJvksbu+v6m+w1DZjv+hlWNW/uyJTjHhdQrPj2Jh1q6HiS3as
d9vRFSTMlYJeqXX4BFSpd5hDcYjfdT57Jq3eKx8wxpLXzF9YCg/o+HAslxrbvTzcSR2eM2aWORLC
jStCuG7fjI8nB/NL8UVgKBsoY5bQoy8RnIMDmPck9N/kHHIETDS7i2MJC7WzmeAhYTl+XgbeaUOz
ZUhVADmQUUNoKaqlOX2fSaJlZwIcAMa56MS8y1albLfEbmExKIUuZ7ySMWqJyDdPTs9c46a8Nqaq
t6trnLLOTNbVts8kUCHL3XKx0aTxMHGeQyEst0/bubgSWZYVkqV0jP12Ri5kVEK0Zc+oo2x0dHVA
cgAS/gwjOnSEyOiN54d3+x5g0MGcR3YoLQbkZ0DoM2ePopVsjUUdwhMPUl3MNpXDNwGD0Aev5SCI
m4mVpuh8QWTWBbrGLjn2INXIloc8ZcYrlWMtT56ADIat2/SMgWkpN9sN7ikstAgl1qnhf58l97ee
GY1NO56YPZsxANuF9bxreU+Ykdi8C21Hf1NEji+bHS3Rhx4u+utOHfgLKbp+tBWL3ebFjXRJRrwY
TmwQDIygSNQZ2Wlm0jIg046ksQ2oEdJMUoHj2m1LKhNegbK+OmwbPZ4RwhZaYI4YQJOTypkyE7vY
w9kTFR+biInVVyfz9cxAXF2BUHObgPd8Qq4HfGHaTwbo3gu0tGbqeHBM0M5ZaD4ks938AoYMJ7Ro
kyG8aJexifILCqLAQjXiYeKERhx0xnD4wVie5dwdxftWc9+lhcF2har9Yw/eSLZHvD877UYsuHmg
EDaC7EPUt48u9iwsZl9tHDflWo5J4rFQoWdJooyEzuzLZXM+i5T5uASfjXHVsKaFvH0QZRfD6SBy
k/JwBrGS/yK6OZshj92Yj9jFC+L1Wya0IA5awL/8OHwgQ0SLu03KN5a0sLXxmd3M5IXInmjQ2koi
cchugZeZgzjhPhv+Acd6cyN5o7VeNIfRHO+GcPJW/rdcELqdS0e8j2gnZoqLrMawhCcVSgnULGd+
uGcOrf/mf/vK59Ok57QQXLh+nEjjaKoHk8ctcEb016EoH1OAlWOHJtk0YwA1qKBSUbsWYOTF/4ao
IhDzk3WZiOsiQlZU/vqkj3atnLKqx/sy66JXlF/0IK+Nxa6wwtZ8zPc7snuWaC8sgb2TEtk7GYla
h2sWJ5PxlBVQD0+LQtsZIVCqK0OJdzG4L6mOcSsGpFhg1FlHqYZCe6Bpisy8MnxGUGT+UdFgzltv
QDA3Un4inxCVFadm5Jslkovq/iA9h7YWKtfxZFi9r6ZgGDXfdsjytFzgI2ysa+FWOqPotsNEz0bT
7+YBzxEgNgS2epbxkEnG6ryvxT1fIXHp9k3CCrwgQ5iicTLzADyhWxLeOrM4mzeiQ+yJQjLiaCz9
NP69FnCsfWDCA50idt5ijkntjfUaLMeH2T2ttfKavWsnniMzUpr7PY7yrzn36bXZZFvbz55oekHP
HQvHT6iSGwBpyU5exNUjq5tSX4oaA8bR4G5UvioyLHRl2mpPGUKNzsxmxUBgQ6KHc1dvxiWyRxXJ
TC9njhg/cKp7XfvDar/FDdzphTsKwCbcFq7yA4cLVJvyKin3PsmXCja2wmRTzxXMw4ib9INGZeYg
CfioHcnE25UarTPQUURfByoNeXfAsI2m6KuOU2LRuFTHBICzWKVCOxoxICtHCxK9WV91SEGaLH3Q
oV1BYr4oP8CTs739KUalsroRW1eqajU5EJHbZb3ZQlyygkXhYPTIDlNndIEYKSFzs3I0FVcdgWjf
dBA+LKsQDLntJeYIyPbD3GRuGo35qdNPSFmvasDTwOcZPMJu8J3mEYJLmVpJPxX5zMnJrikSpSWi
5/P6LtPU0UJez2tfKlvjjmUCmRi7dhCP/ALn49NUoxYu4i+9dyRvyYet5eQv2p4lqdZzZGLCCC3S
iJITTED1y4NvMK0IR0zxUMitgY3uDSvf+gWlmzruVCotXud+70BnMsfowqEJQBPzgvKOxAWgC+dt
+DNuPz6iZF/zWuoGGTZtFb626Sv+GR+doqa9qcMjJMXuDVx7It209CWcBOUN+j/KAdOABYxVgmSa
fIscW/wZqfXKOdQyzP0qKsePGh1ipIWt/DKFbbKG02Sj+a4OPoW42vXbI/B7GzGd22KjkeduG8Uw
ldoWO3TZrNGbcSFn2TrRRoPuKrknUIXecpRhCLzu4bfGlneG6eZ/iO64vI4W18zMYxModJxNoa/T
nJcWxwiCcm1Gd3MH7KBuDoFD9tObc654Ehkr3IXIPbqR3xIQ78Xufj3fA9rOvUiJ8Tvy30Fsnqyv
HT5Ma2ZbgVPzlPstOaszAbUKlEa76MW8l5/zysoFx4w/i01q67eGA3a3XNw5gQKJBQRgFcdTlKjZ
6hXaNAm3qG7SRQnv3xVowrlsH4NXicZxRHCxBlK2H1fCScx3HB1bjg1GCvQrAtnqxWvg9chaq7RA
5woC2oPHJbxBObpWEBIsVGvOWYtjp/RvQov30VE/Qe7b8QkpKZCrBtqmus+xlH2e2Lo8Pc3x4rhA
nQbFMzpwqyP42Zs3BHFWP4wtuYz5e/tpyz4P6NiIDZswAj01sI6+e2ohsnbl4yN915QvGxq0q73v
lvVwPxum8MpKel0MaqDwi5LtxRYAPYTc+fuPpwXMm9GSGfJlIENadfxFp+HZ938TfaYYxHcsF/jg
8xy3GttuPGz3xwTz5N/hms2x1z5LfydRIIZPnHDME6tP1ijE2toPCsulRnCuYLVxZvtlOhiRK7l0
utbqF0CivZXGqZYayeNcXr3BX35quSciKahNFBr+B9RorakUKSNRedwFgUy/m3e9fHEGJw+Jh5Np
c9QlFtcZl15S4AXMgh1ITciUelG5UPQYZNA+vMCJCcbBnGxRf2ILUCrH5QKd3OpU1U+rBx7Vpybm
8iw79ZVxafHGiZ7w6Dls2GrA48uSsLynAKq7u6/zkdkheWANHmSbFYV8yg6hBEqC9O50UJgQS6FN
6ILSVF7GbhxQA+rt+3lxq7dxrTI+BAWrg0t1lYUZuKfN2WAbqA3Ob66g5T5IiutkyOo8hbmu1KWk
kvMhSaCHSFeomJuuuRgt0cyUPMT/8/dj2C1NfxCGMHf5ZFhWSb8Ikbq/mjZVFMSOZ9O8Y8jbEwRN
Q20QRkckgp/luV1DV7togx5W0PvfQDU3svQyuRpgGvHBz8/Y2V4Gk85uH2wk1RC3u6rbBE6qSmaH
20SHnJaOC/kUbKDJKhF46NFJvwWfo/VpEcpx5Yx4irCS/nYZ3JQRnjUtumzUGWSm7QFXaP3vStem
CkkDHyn9865FcIdsbSpRV+3S7lWzHK7newnPdPTOV++69ps4g69EEvP+rFwUUyC6MeZYNqger3V8
lZE9bilRyV8yefoejTw3FbnSJagDPnCuqtIHcwE2o0I7S+auTng2utmJZhN310A4mYqKBv5SGBDM
Qb5ipWu9cWnetadzwjLj+HP8njVaReRHp8wdWFNOTzcDXvFCcMmFOjqiVNn4hKHk7nkmKRuJvp1E
qSDanUWsb15Q86uTPxIieDw343e8iKiUfDuygNXtPDx/x09WgiFoo7reO7Eo1bThcfzcUvJ9rbxz
KPMeAwanHfft0FS8V2e+knkprfnb/E3N80kx7RP5NXEjggbejkM4bCYhhCrBpQII8MGt6QNLR9Bb
Of/YSjOt3tfwwMGP+fDvipPHkMO4VsvHOI7byjCJSoHRqTtCwdO4fWEZijwuT1H+jNnqnQpURAUI
YvbLD5AeqcVuq2bOAcxI/cFuZ852ae61b9lPvyoasPBQaZUhJmKVRP8M4A02pUG7V++jdIkEaWvY
F0+Cgt5jEuxtldMfCT1mOTO+YpCYdRAWkcLm80LncV1uOp2BzgROWnlDWpSwXRcLC4q6Ku+i/rGl
HHneX8KLF8ABYZB5rTIOgyNMT5+T0gagZHBJIw3+4Cf6e/QWZQmYgC35AeN1InX313JEOQm/3z8Z
/DK5DPRwvualJ1EGE/5W2irY+wJ6I9xCqrT3YHC7QLaPDUDDhnLrJ5V40KWUo04jB2m3HabIoikv
TsQZ4e1xIN54YOg4ueKRMU4LEjf/2KzjlggyJanANWJMpLU+5na9PLUeat9LGLcwr+PEZyKOeV3f
hKMr3RfrgkzuBNh0fboddfAwg53w6P5yAHHPTNJ0QfbsqptOEqGH2Y3j7+fyVk2lYaEjBgTwX0/d
KB2Cf6wUdCab66nHJ591yCUmWVHjyuwbdOjPFYgh6CXlSv04KGf9xivsBbOcDd0B4W6MmqojTUgc
34t3+6P9rJEFe04CyoipGUhYD6G7vR7JIMj5Xyej00n85pKX29Y06U1PxV0fyr+1zW4YM84FamXB
oxq2wpw+amB04W6tkP/KMOREJE87ljh7rIt2PJakpA66tYmOdmjH456Xh6zbQmfgd4uQrqLO2+L2
U6IqERf3+1Ew/aElFj3L7utqBCdeZnr1dwYtArHLiMepPmzv7D5/g7QMpiwGgvi5r1VMExaRLgLg
tzhCf18PoXFJhPJj5P0/P3FnbAj0BGlzuxLPi4EBiEY+u2B5mOYJ5Cx4PoDUx9mvG7iytWoX5+jT
vK+vJ1o0feG5GHXDIQaSZ5NRA/o0JwE8Qlvxp7RA+fKepL7oNli/vR+AGtA3B/jFpDovpOLF9u+a
zm8awDBBpbCw8GTL3xk3V7nzDm4VgP8K986YoFb2OA1EgAqElaYqeHQXw8NSvH8jn9BrZssK3x2/
d7mXFO7nGIkN6nyEPACu2DqCPQ4OApD9AyhLtdlbgKsdgx5KuMJATJklmJ9zHG5u2NOJ8Ia+eSzF
VWimzTasfSlppg3FhdzFIZBG3/Q66BHbT/cHKM7oHJK9LDIr6p4wlHAhGfykEByxppXPVtPmsDK9
Kl0SQJti+MznKryfrS4MJlYDo/IVwty30UXzxRTZ1CGssFCVYnYY7eEjPpVfX/M8Kt1Ji5rHbYdB
v7xfG5v+hGmpdKnOgppoDdsNrn8RZWn6eTpu44/k3e8KffHH/cgKrlN0Lb7K+slUYOEWAqdoHIRz
DCs882ztV0Zl7tnr3fvu5lB+GFyZjuKzJo76D2INrRc/TmeyFsLEms9jiaAad9uA6iWq9+Iz2fyp
h74N0PZ/DFAPMhshdSWLvPSt5N9gCzMK2HgYDk16RboEcDg6dv0y5GehllsDxf7XGGidVU1ohmBO
42C4Ilh9ND6Lmt+5m83/T7VOgmJZxY+N0oKujPqR3oqmJwHRadQVyfREWT6r4cawOAhyqaNDE0R4
2w1X48c+dXx78w/Z/OR6qCPjLOxAMvI32a24LUKEVbgWgI7jPbey2UY5gNVmspsVQorgQfjmjLOC
8mMEnsK+/c43yj2ZCZdA5hbZg6wCHMvExUTA52uAjt1XP6yrLwpdijd63sYeC+6KpyY/qQvh6E//
ZTb/L4bxySVa56iYmIA/cKCtiianIn+VoCZR8G0LU0Rgdtamon+Vgxs39+cPV80Rm4PoUga7VJay
vNFkn6nrPeEkLsNsf4l2nrjvs1qJc6cDNspoXIdSXTLm4KbeuQG6Yii4FMXhc6KeQUPmOROcl6lc
EF4UrRqZu4p7Oenufuqe3n5Nm3JsoRva1MfSf8a9YMQdwDkpvHKqCOt8YOC3IbdqYDlbLnfGtV5x
Y2OxyN293ez1rlPJZ5qgnWgdPYUsfESioGGC6WlTN9qZHRN3uaf+voAzegcvteEHl48BxT/goLqC
HsI3TQBhrKmDKFiM7WF2Ji7s71gSnsRmdiKjri2UZFIg0QjR9DUFn7mQsmcG4VEvRhsHQc/PBngI
myREaLeVe7booBDgn/m099vbeKigeG3mwErx47Z7DgpOrTO8gB3Cl775XZF/F/A72gEyX2wks3sg
CCFWABBmW4UoTSGbp8bHI61tFODRiq+6gNbM/0oB+S/YISJE8D0LNH2b6To2IiNiKnTTo73D3QA5
r3L8P49C7kinm7TFXgh8UeFw9KoizP6Jf411v4e1relyvjf3X2rPueTYqOU4hKa69/hSM3bIb2RX
s7nLENc70Aq3h/J2rRCMvXNe8kN8Mt7L26QkrHzjxZo5mecD6/HG76RZkiLl6csEJ4uWRF8P8P/j
Ms+q4hnyb2TAekstJWh6U76zzihaxZwEgT6pZdaQtkOViYQzZPhG3lW33ktX6GUU9O9u8jy+vpHm
4UUa4cstxL/UqrlITy7CeQxTUnWa4+/Pn7wt1WWsAXJITGQDQyMsHUQhElXTX56fNJnsdI7iCzYY
w7d6IUmSiH+ykeYg25wM3C746tbdeS/XLHJjZeVKCQAuOWDqlrRL16isf3mr+yrvgpcY8a6tcGab
G5rwj99KGled0LnmRFxrKldHGv1WwZOqVrZFS8bub7YffYppFmQu9KzkbIcQYsTeUYxLuZQ7Uxuh
nm6LSNCWDb2Jr16qjTtbd/Wfp2UCe1n/5MvQot/gacxB5/sJIYhXAt76E5DEtUMq55ejtGzpkHFP
UbjPQ2OrD5I9bK1uzod3BrOqoDFBKXHfRglg8Hwt0FXMuximgwCswG/SxKObZ15m7EBedXz4pvMY
fKqhrHltEuXO8R5mTjF+cQe7Fm74c+sFmofotcw2hIhed27BmfoMc+fxg71zbVZJDazWY0ptM3/b
73H895d8UK2EuX52/L9zIrm4NMtwBZIzyZbUPwBGbLfS36gAIuZgYkG14Kp1O59NlPUurUdtRX2J
WURcc19eQlsx85opX8d25h+XuNR/a5Y92WzZHrDjuEet7su2IsXoYtuACVX0HlO2apotJ6hDcVwA
6Q/y7mRTj1Xb6P4093OSyXhGwpqh8lKunMQtGz/T0EkswA12Ckt+KtAg08ksoHCnIkAqyrSrcc4Y
xi5anU9GgzQkxNh8PmaCAvj4nf0b4ZC5zfOi0Jq7n2f/fRisB6Tob3JVm1fqY+uM9Nv7TEPk6QS/
UJweXekOS5ujN3DbE18EVznmQAJYSOm1TUcGIPqKC7WfTWIrYqDQgca6XKrsgamfC83PJMtR7vwo
lOt1WHhnkjb8DlEv3Keof1W1ySVN03MSLHhZnOjBW4inmRvkvEIT7OhUcClP1ewApq/0gRkHK6i6
92MC8CGbONBqo9wid0WetuWEkKl/Z7HqiuP62srPm6/SXNjtAz31hdSNgimb72todUcU/4jeMzCc
VUN1449vY7CRBv2tG0LHzYEzO++jLJ4jvSxf6PrkVRUis+1TaJKSzf48BaH9FRUkCDEexeEHuUd7
XUxyVwm+kKdTqhxzN5Z+fG1qPZU4PpZBadrwyZYuCJJIKhxWsM2FVT5JtFpVVkf93EgVx3mqOLeP
1mqxGItB/NZRZ0iqy2zdkPXNimadXu5q6B/elSfdYcdY6QP3E4pCOtplw5sb3d3xds1dfEeK3Y+Y
nebZaftftza/75UxYWorlVpQNudMDQ9HPRtTS5wB33wtpYvO3tA4/Z7A3Iy/Q90Uyp9tSi3lMaB3
hZKixwOsreNiOIC5FyJiRNIjoIP0okOl+y0YMTH2DVGdEuhZNI7BsSi5TYukg0DiFfKVomMNa69u
DIp3FMSsQJv/CjZjtM7Jb/ifjsoVg/qM5HjtnuNuYHMd0kaOnlOX8KzYGrzNuNnr1mENDQLYooDY
7BKbXXpQaHdTAJky4spcaUlnkl7iOAbmo3Mj8nHhjZs+DH1c+64UIPkMj1b0RfuCmLptVlYyBbF3
N/E4nd9OuFaFlQzrzzUXjelTTd8au5PVJa8/qjmE81mIO43ylHJUYkxOYpPD4VMlBEJhkiqjmLOK
jYav0cvy27OKA5aZGA5mS4L181v3Q9M6hcT7qp43l0noYphxZg9bZ3nwWXMo3uw0Hwazc14qP4VA
Dm5Kpk20vop6AS6codFqRJiOFqSut9VS9mBR32TK17hMLsMPgHjqKxAJ1rFxK9k8gnEwQIWoZY8E
huKczRQ9RnXqzdIMZqevmAn72ei9TvPvQrbiJcxlXzNAEj114XVat5phCbBEl/ySLuiT7WQBBpJq
i+oMRz+29InRLAJ9EHN17kJErHEJvfjbjCYVsSeTHx0x+Vn/D2wjaSdipXLbztiUQqiZb9Oecloc
PGF9xHD0H1wSt/vS+cRHcohUtgslUhgC52/07rpf6Yy5XuqUAfjEaRdsviQfNv9AD1gPEGrlkR5B
G4AY+/dsua+hMVR014Gyf7b61QrdAGkDz+33PgUQLutMz6ScTZxUoh+pk/NzvjKEprJndyIHO3yx
xaxzOWxkXmTpHngOcu5OfcgtA++RHRPAZAbSauflYcFPdyPV2sY5OKOJUjQCUOYN7mwI+KT5KbZX
HREMAC76S+zBoNXIg+Dl2rQ2OHVkcs0YCSoQTw1Mnvu72Z0JpwMKPR3nPy0UyEtj39BJb14kQ9+5
WLJ5eUXcDVWyZ4AwQWqXFdx2+F1WjkYgeAOaaKOC5obVq5Z3Gcdlkqp38vrMYPNn7pi99sRrwLSj
JzADRBHWObHZQMtGQkqmWyzwAKkkkptpBrE5RmzsH7u9IN5WjHJsZftbAQo6c0N9b1nyM3JLxLBc
Q2aaQqvoDGMY5Bzi+RBg6OBrIM8c8yciizZ94pKWMMNJzZUPAe1wnAH+i7631gqlCK2FsX4/9hsT
O/uGAFFIaQw2VeQ4KUdzweCMqMq2DPzqdeXA0X5eF1pd7GlA3BbePblUo5f7YZQy4MGnQr6Mgbup
OjdIQ7IT2fdSSZCVddByqB2yqI5C+jOvGl0pSOMeFzGbzUShuOTLfSvuW8sjtppVDEN0YHxrg30k
/2Ujaddc/gSBDCThaR2kqjxMgYEDFjx0OwQyzj9ytIQ0zfUadVhzKbRlBpnjAgsD6jWXJ7bRWdMY
wVRFw57u2e428HLMmwsg/1gS+khACHROEfGg3DNr5u+FT/Ju24wLBTpRBhbmYS4wndREykE7sjwI
LnsQqrpaqb6jf4O69pCatIqMfJfMYbR/en715u1b3yKgVZNNGxDtWEYAyDqOY+ONpD+WD3M3sfcS
X/HF3o+5+6ihg6G2qGMfEQW59DPCmRAwpE9lZ1CGK9gWE+BAgBvP2nwRNMdNrP8gGrzyhchJ1QVK
d/WbQwf7+8+oKMbDzcOosoGJrlcK6lbe+jGJ/7BA2OAt6Lci5ldKQw5X0T9uPDM0rCmguFQwn6Qm
J00FzSe0ljWXFVhkhnPI4/x8sOiPP0QGHi+JxjZvUkMHKpztZegvidg1x69cWzS2OfpCMDb+9r2q
y7LFnIpvaixvHNir68sB2MOe5WDcz+1QBiIecZ0royLUInsdq/cM1P7TzQtxYnXXoOUGarQYv+tK
XCFvLEgGu0A+6AnrcwLarZpuRb+Q/yPg34MXVy/IWIz9bYLAmInerpKH5yf1tXL1l6Ai2aOXm6k7
2hQRtQIlYMVtqnTqE4scLHxJqw0nsqkqxJ9nsNuX9+gIbF2N8vGl/QCCUJRNokt/HgK+SV8+WNQl
8jUs7gPk1mEEdca+NqFiVZV1srHqdYpUtdaTFJ+/0/M3fapzqA7q8gjMS17BLA5QU13LrZigVSI8
MbVE+YXE5YM0rE5YJNnsMoMO0fGQLy7r1rJcruxGkMw6XEMwuh/LPEXL4FhyHehUJS+byAh1vk0H
N+gk02zNGX43KOlrW/GKoEyo+T4acGK4fJ4J/XjZcllJlsCdTNz+o7kinvCJydyc9ac4kkFbuh7D
tzCYwm7ETtDzeeJBt1UZp8Zv0KVC3GJPUXeR5n5Z8doakx46XqaRkADUY0Urdpf/j1Vw4SLd2ZxU
dRNRrYS1fvdD/HieSHHu0QXLVZdz8pbZjd2bnjhYbzkoTFRZkWK6edaV1guDKxZTjZsnwfzFTUPY
L54SyQDWFUwAV46KzPn7L7lHl0srX9FWWceWukgT6qr5AMWmqnh3127PLbWpcl25uwyFKDHguQFr
NRVdckYFpDvK19sv26ALzA0qYlQ0SURUo77+o8weqsO8Q3JH5rPQPSLwEO0oImLWRB3G0dHY4dWB
7X3LWX0xag05V+xaBOJo+gw+Xl1O5IhjqPlZfsCC8u3ZiONMwI/+h4YIyUl3AoAWYY3EEpxjiD9R
iJKC3jb9+47lqqstxzNu9iylj/EG/lvnLwJjBQ+t1x1a+LftppoybTsTv/I4UETa4DwVqPiguWEt
DAtJqcvOhbiD687UwlZtPNS47OcB93B0WghFtMtIN7dh/fl8nUbpjdHqOYoAR1hytwNHB2OIpK4P
fVFYspqQQHhE6b101nySquMTclmbbuOTtf3HgvRZF44fxAAcHOMyUyRwhD3R/T+uS+8NTjN4zMlm
Kwu7ATnnLJKD0ivRwij6N2dpdj8ic0J7BmdQViXBQ8HCHCbvoMk5DKYsxP8OC+i4PmE7n6DHtVVy
uN6Mv+EeHhgDuWGXPeqDftWQiXwPL7tRcHicyjOro6+xKT1fe2UP/ujXXaBOqGr5+Ijh3GI/01l8
RWdgDncQlRFOho7K5Vc94cZuE5vS++0mWPkidO44TjQfHQbzupYqOxJgW24eceVplgzDe3LUlEHU
KzC1JD2xlAVohqcmP5JUXmjHMG2WxJcvjVNFxpOxxROFFnSToqSZTYlaHPgqu/6/FpEBLc9cu4Up
t9JKoBTevsrcpVIn2QXjxneUQuO1Cw/yLnPi5O8uaqm66dAIPUNyrp8JUIYbz+oeZ5wmyc5olUeA
gPbj4Hm86n5lmzAm+XjVeIjY17rIDoyZnQUTsgSfwxQbZ+Ueg1djh9gkh1oqOzXw1H410nTHu/OM
0bX/gJMwR+goFd6HfTdy5tzCK8fcUqeIiITISzz/FyT6JCTbGm3FVVwcmzaBUEQChB4jaKyTRx4f
Bo5HEgLR7MhSXGAoVjIdnZkdylC/ShF+Tppz01j4fzKbaAEa24DrkrkkmbMenIuUXCZCsXEM8Y4Z
8f7UwwNNAMMtIhhxAxPDivFviuDHDOD6fc0VzIi9PGNFgZKnHAKYpAQhXG1fwYsmDFb402dILudq
teCeH0DFVxuHQS4OOiz+TeaK/jlyGowaQTchaop2rIQtjjar/6Xsdjnz86aHLzOA14Td/QoGejZq
TGwKvkWXBzr/q9O2657qpGkQ0paEPaBVhCeLVdhLLdqR3eyQM8jeVQ75qKsdv42AT/2f9HbR58SR
1sbVyA7mpPuEKxTh8STyi0u7RFvSUq9qsLQ8gHWBgIVjDPRNif+7Oe8AdXcdk80aFJYaCRcxN7ME
Ja6YlJlor9j4iDRfhx4WXsF+rmWErWO3StO+8TwurHC8UXDqwck6uXtVCkne6L+EeFGYhZ0yiQFR
eMVwvGmefZMdYTxgyfY6jal5QqJXJHmUJ/VmT95ob3DYjev6f7o/GoX9Ev/lI1KjRWUDNtd2mHNv
8PqSELaDVd2PSCqNOwI+rb6cGachxodVT/RbfvJ53HegVWv07FA2x94I6YeAzeQi8DbRJgd8bc0z
m2hi6qzHzRVPupHSY8AiQJXryjIrc3B7qZYxaPQZ9lf9M3iwUrr2vAhe3LyVx3UTM4j0vbbLQedy
tIj16tumri5UEqu/2r5NiUfm6b4XoXTmHkQ594RUD3uXly2PVRJqUrtJ+JBpNPG0+7LYB8vl6vVo
8bkxwNkcIIyH34Ifhdt/wrzy7SsiyyxQelvrOuF1TLEfnGcKR9/hTokprPliJxeR0N9V114e6ZCS
3yM0Y8tO80z96jgXFItpFrGte1P5i0+TcCAXq/aiKQHOc3uS182Xfpn6xacB4FcV1CsKGhtwji0d
wCYoaETxqCRCClM6Zou400o1QvZky4MyuwV5SfXYuvbo6zZuLxTYbqO+wqbmD7v0e7scwMXBvh1B
KRDostvT1zhoTNUl2/FPpUNBOAYUwIcs2hGjQi2gfXEG61vvvmSk/r8xmozqp0j4QGghO7FZWzkj
4nh3yjKwwovwWCIrYHPoP7cpz7Mqfa6v8AHu4KUqfx34pz6TF205AJBEGVk88vXzKXpjWPgQ7l0r
Lf4sbqJu+4sxylVfMxnNeScPyScquZrpAy5rN5U49y2G+xyGhhR97/+1qi/4NS1kHHYflSBBBosf
+1nTjXc8VOMuFhT10rGz4P+qBQHFCxUiAvBw709HJfYRCMt+FD8K3bYPuOMUpck1A7/y7wdFNgU9
0Ur4zUQTcVgBNCQSrLyBM2o+u50/JVEUjrKeLBuNGsxzG8s4xMHNhTTwH0C6ElPURyBT5fQguDU2
AZPGv3BtUnJlHVEopXefVNrSXkIRIp+2GqMyGNuW4q7AhK8HgUAFo5RAL+epReTWs3qx4YkhUP7q
eSbrafVsXZ9E6hXr19I5BneC86shF/B1HYR4x4OPOAPgXuhZvSU9E3lZIeELVhMG8d08YQmUjo10
FrxEhS60dW4Cl7eLTv/I6VLUW865BII6ATiCZ1d7VjARi5nwDgZK1BIqKoE+ZifA0CuAoQ+0NF0c
/juHw9HZLCbNSKg2hGvsxz2PQA39wJa3vbTu4AoNOX8Hn+tHMjhmAChaP/NBB8VcCDKnLCCf44TQ
IPjZx41LPRsNFQk8gRWHPxXMLD5nCjWK0dQ+3jL9IWwk875m86YbtqpmIhPqdFh99HUqd8kKW/cz
SS+7xvw5EezzVAUhUk9Tl6UsCOlVX0/+zW82vo/rjB/BIcgtrFQOa61ECjldmBmZ+xrU1Q0XV9W9
yw9on69n2hzI2+J93/EI7xztzZKZZZ1jkraOdtIpPE4ubpgRVDmQVW7X+RkvcGWbzQr7mQqOplRo
YuJfHecO8ovB+m3k8Ram5XU+EHNi6J260fFjgwrtAK4YH8iUHizLgIyNMGHeV/bLfFYeHAfccay9
J4sf36dsa/rmLPH+5vM1jKoaccLuC6M6gqbHMMfP7NWSKENiWDAxP0QIdTjtt7+LrVBmkpKrSrsj
QiKMzNQ1KOSB9Gu6e7MRduC7K3fgqdr724hcIqcuRXbeDq5ArBc7waRqIa3TuPieGhqSvXSjM5qy
USMugpvHJXU/T1eJY786a1In/fyBvvbPxhdjxb24c55syDUqQOMYarGDUhdTUPiFXr9Oti1iA+7Q
5S29sbGbF7o1nbXGIlzQt6tysfZ6ZiucBFRGTPz47y7HsaXyBJVcThtZ4tvW8x3r84afL9nSud/S
kuwfIl+suUZ5P43JpkBsNRRYRAoiYA4gyhGtSs4k2woHlZ++I547h5IL8Xiu+LlCyvcI3T0MI+/O
CcGUMFVve6XhhysQTkDWgNQvwODHMiOeUb3ZZAht6M+U7AFfHNNFdF7kFZWvLLH/u4pfTrmlqgUw
XAV/2UXYZ2OJhjB0Glh3khwP8bDf7Ne0IE5z+aVbUtJEBRdRXkDqiuFPBqaAx98KpLsh6+H9NE3x
naf7Nd2ZG3YGvVk610uVmVaoA6utn8UtUruYUJfSEAGnICDBlEn8r1kMxecsX2RHvLOP/2proRwK
0ji8gpKTt+pX0qb76aog0vVrsUgEAd5wFNWJ3tt9vQWrQhm/V5o2gsHHYL3SyWpQ+o0dHXVh3Og+
/bDyPCM9F8M8uQDRRGKEpdKtEoquB1JXbLuZcgA1RpvdZrYPtbCA8u0FkdXK56vqIHfqkQbg3HzS
vPQ2LDKEmfD3ZOSYAU7RKHpMoi9reBcwMia7ucI4lhsQKE9OHoXQcnoUFO0q5FNMUaFnB9GrwKqg
SFkk5Z6O2yGDIXHVmyGP/a/X2AhcbEAR1e9NmrN8eHi+m5V/uVv3h+hBf/kMoxBjPZdEjRGySG7r
Yp+akdcnjtHNWJkKrKBmUcyho/9hOusLe4wG6TwyLeHSoPH6Kw+SIjj0D1gMhT8DcSSFiOroX9r6
Yohe6si1J5DeIs7feyrMCio+v6qJ4V98BMDqo4c0dea8VpvpCgUUZR/v9XGY1KwuxQmlyQ15NMO3
eXDi6Qa09XOZuY+Ybh/VKWH/d7SF1jA1dcVW6XtNkxT80G/c7RqPqOVCi8KINNS/03A7s8iweU65
61GCXCR1eB4NvzsN+Qq/22V7XtvGJNcW+vJwMO3KMiaCcs/n4ihYFgvdI0gKfRiY7hp+g73MVWr/
hTbeS2oS7Ch3PtRmllpFZDiCQvAdTUzOMniH15Gs+WqaBsej/aCx8prslaMClsQmbHODeJAqQSg6
HECS8gX1Cd22REJNIFaAKokF41jvL6FeUodJh5yqgAClgXmPumgWMwT4jGZuOhQjl4mlHr2ysUbO
o0OFPJujZfwplozAVRYcdwYni7tZlMNBlvieafpxsAJD4jF8q4g9f/VTb64BiWZdwKlfWk4jFKSY
ScIXC7GMvctphEKHlB5luohMrNJH2q/t+msSTezZpmCiermLXBklDS7xfg6ulFWPD1z5wTuusOo4
XrwNc6TEqy2ZqNUH2c8cuwiNtvEZK3RrjtVLGJo6J9vCVE/b1Eb4eNuWp+1aKGWjx6eHZEYf8ua3
mu7uPtG/DblthXQyz6MnqI7uXxTYVlPZgdKgSR9HRAaYy8MFnq2VvJMR3qMrsW/LxaaHC/knHwcz
Hakrk8rNdRnwjeoujsKAUXV9V9DgTYy2p85umyCCCtAp+d9ktMvwfHbYHEEOm8A/oiHX1J2VGTNX
8z8cbbLkdZjyYlVkYmNuFvYux7U+nnaTx2gC+TsO0btUi83A+lfoF/b0AeHEdx1EIm8zcOy4SAHM
HKOiVyYQA2k+bxpmMnbHflVo3YMcdattVCwcgSqDd3KXM/zR5xjVNA3Im5i1qdNjdxY4BTplS8mm
vs7cOYyk7kTUjHJejqPEGtNqdTeE80/7/KSVz1zK9Kk8hrk1qihtG13Vyn+QQxrsyP2BRKtVbqnA
uNV5x8bTYZdkzJfnqgnW+GOkwBaD/snqHQ0VForAbmP9600pknlZZUcuEbKfFdBmrmF76L8eWWX7
s858mtBHpqjKS+pKjJ/X9TzKL8IgaQBAO1lPKwecUNjBPpxhC75AAzHt0a+F7kag0n2Y86qBHxW6
y6WIf3khW3wVodBDNzgq23Q8rKZGJtEdmmD/cavL/AkSQUiI6O6hfsBW9sOehAduBWGLKIWTCkXg
Gkc+TTJXeWtAOUxcetdpAc5Ko0ht9hjvKHZG7wYXX5PBxvCFSHpzFEilF4UjO4wH3cmkc/oEbJF8
6KpAt9XPGJcDru2z8W4NvxpCn4sDZP0JEQVxxmGrw3F6IO28nAY//sg8YlSH7OXCgkEyw2mjTMqd
LDuDvCl+wrjh2cB7Qa7TPOyztoEHDhDknwRBg7ouAqTV1EUR/ed7d6MPspfP4dgZIZ46H+KT+24w
eS/2qES4PlnwfQ4LDXUIRe9G3zsscghKiGSot3DNVWD0zJU83iHos208vIXxPOpX2KvuBERQz3uU
KkHiQAn6tbnIZP0aV+Ka9JifKpTeuveiqDI6uT82IHVK82dUOWTAA5thXRj/r7jkJgQyaZ0oDVWN
4DjEf/pEsZYyCKjgQG653i5fWvwN0p+U4tXoHzlAPyj8Xl2Ai2yIkwzo9tXrgWk38PflLvmTKRIy
fCBjqR7UI7i11oFIYzhtFkY5eB5uySmeOLxxxY3yhfy5+fExBbFYuZADKJcsjJMOyz2eFml1A5aI
kjq8NHXTant+1kEDolf+STPr5wuGbrRmQ9ma+hWF3sh/8wUTpgdhw8BFgKLBrkRxhBdp9LlF5Kkf
3Lw/A8yZgtOWrRoWS8Q6uK9kMOhjASQ0YmCh2GAKwHYc3S64OZAo5wNLlSkeBpCrRXs6Ui7g/3KI
PQARsnSGVmhZnsAqY/Ovpvh6aJm4RPlSLz6pmlTpKn5LQ1fD+vINN8lTIbQwy0ZmGeUEOEAavM0o
VZJvUYTlm7IOoryCEu1ClLjgUWH/SvDpL6gCgup06GB/Zbr27h83lOMf75IXThYfXQhum4fMMMVW
bG0n4vP2DFxPN71nYYOWQAwdbwYIbLl1CcYSAkrCsYbGS5EXrlUoErP0u3NQ4NEn75dqfe/y6Egm
Bwkq02V1nWd7MGQROtoqGOIbm5h2BZbREvmuZ6RM+p++stEGAEO5A6q3nZsa1xc3x+N4hQWaGRJ1
FD9i1Fx+zvV/H2yWG7k2bkh0GKir+wiSwXIwJMmUqabnK3Q9WlIIFdy2+eEn2n+xpAgyB2z1Wq1f
7szHdwWy1GNze8P4Dh7scw14bcKxivbkA/CAfCOVz1pxPxBfdi/XfQmT0KW51QjXNM2+QjmeZJ9o
8R01bnr/vCQ0nr4gLCS2oo5aWI06TPdACHxoO7SRsrR2Gc2ZunmrNZ8iNmG33mK4P69095JUNHBR
LDlcKSBaq+6MgN9k0l+OjTLKdezqm6hZG2qy8dlqKWmKMeNSaEOi+lIw5Qhi6fHUxQSoPt05QAwA
iXuMv1ed0wLonMNxMuMdIonmrww1wFSveddQTQEXlsy8dOf0zSlExYAOpjGtUJA+WULNnnJSI3AX
onDezKhzDDoBVIkZPkqTOQDLdJ3DxBf/puoYZveMZ3p1kK7xW2yeYwp3OeaDbrn6+q2bdr+Evf1S
jFWKragMgeaF3qh/8ttQ3Ga6NR5Otre8JckXsrIuDl8u5rbkHjVQLLQUPVg0mOZzA4bkxnniHsoH
I7ppZC3w0dBKxowi6TaQFu0B8aCnmOREzi/WxHxYrFDdMWHhur4/fxjDQ/c2a5kkeFii1YevZwhW
MyDVY76vw+TDl5TE/xDKuQc8ANrU3sTjeHL3uJ3wIRR55YV+DBOXarGZVCcc1dH5vmqM/buXuOic
GO+QUHfGoCxLKBDP8A0gEsqxGH4Sf21PJhQLf6mfwUstZkuZsW0f9jCGVeGu1n2tnjH/Hd3N0yXs
Vf0U5tY9kgtFEueBNL6B/mKL+/IRbVSKEAaamYdFcQgxyOfk4wMq/TSlaXnRMqS0AXC3ifsZeziM
Z2dxuIL04ppjMVHg7SIK0eYzMpbIbAvfYwW6Svm6bs/C+F6Be2cIQkilUDNQ7Q76fVFEkn0OmA1q
O3y5rKHOgBLVitopQOs4LEpomTbP2Ldj1m/3IJyZQDmJAjNAltEi50jYlfZgGtZDSCdcLqabI0dI
NkASFp4K1b6x9U+zcUxd7lfMOc9aEX3DbIw9ySuVSqRsiX8XdRDzDw7uvQvS3vq2WovTALy0Pc2b
h9RAJTvBAk9BpkzyzAcKmx4xwiK4brL2xV+f5JPBMmXb+r9tsWDQzXVx86nIy8QZx9eAa/nuykCC
fOM5qQqzd8Fj4h7n+3JErDe7w8yfl5b5cAompQwK1Vya03OYkiychPUzsYsAScwYGookuNxRZOuC
I70nNWBlqJeNBVmnhre3L083uIfeNEyGmG26zefy6TPcBxhts92VBSB3TBTLjoS6KHgiLUxKwF/a
It8Eo1Vb8FYaA+t3b4yZDiSteZNff05gPn/kczQj8N0Btb3eCIdeDSa4K7IYyS9amLDhlSdoQqpx
APZrf83zdEM8VwlWY7dTj/5TqfbJfxzfErJE/pBH+ZRpBAUb0Zw1B2zees30b/z0O02On9kNYlRN
gF00cAJ1jW9Czk6axCKwmHRvLNWuIE3YyWeIyCOvewdyalz5i1K3Awt80tVFA/RiHmFeFbDbI6Nb
gCL2HqkB/KzQAAoNQzWaDRJy0wJSpa4Lrq7GSrm6niArD56BE24pI0xoCbxchjoAFrgrIG4eIMK4
OtVptDudSDyfaF+Alnl2EhKqJn7wjcVIUwplNQC3Rj/bcERDBvzBMZK15H6/LV9aBASDKaMR/jZP
wGPAXLV9vPZSyI7aDYE3CkdHL1bqaNVY2sOp8NltjqZ/ZjoMQQ9YOINflZxmdxCVAa+IZkVhUAGn
Hy7ZQqjRFjxOX9FWV4BhjEul38SKUYMegizlRVcHwSPhXfnZBdDFp0vuT1T3OunHL7v1FM7tSF23
hFeSCwSN9CJwvyZkFhH+PBZzUznq0XckH4UJ5KJDqB4vp9Wqq/1b/xkR9lwfMlU8tTGusYsqT4qK
90q5aRl4pZXdwKc+I3O/0iwFWFJrt7BLP/Kxb+WbUn2H6y60jInQz544RrFDLSaY4NU517M+MGsd
Ze0vRdaRVr/aEXPDLHG9YRUMnDNN7pOSs1bNa81d9b/DInu5ctpFTFSJVwZ14zIsUJvtGWx7NQBt
jm7cUVPSPWydWq2BWeWM4qkIzyfjHCNxZY3Gr8fRJyuGg7etbpXDt32lnBExYs34CA5FvlIRDo7T
f/flzauAnIfFlORZlJSKFwNG/7l5AOJocCEzQRgqN1EuMlgv23T1gNA2pcfMDDMN/FfJEvFpnNWJ
apLVY1Jjx4Ou8zE+zs4WRlG+vmrOZrrrRMnz5roh0Sgqx93Aoqs/oKe/055kMemx+jBjGyvqzJ37
AkeGMts6O9oB60ELyalyhR1bwmb8bd3Tfxrsfc02w7MrJAyCRpVEMxbr2ZS2fFgTk+feH9TIKGkh
p/zQkh90gwZNoh82zWCAYOgujUl8L5Y7/dLV1Pbj5YZIF7ICdA5LPOoWa6rdjsde3yS45y5d4rIB
RxMMmM29+x5S8yLs3/tVY8R5bv2+HomX1fvwmc8+Fy5tbNKH4G6Xw3vT+Fq+1H+OX0rUSCZNearP
4wOvkDbmviF7JcJYjQKMQZRY1hGraI+5UkCtQspqkmacwX0EhhRnI5pdsOZXF4rADW/RoiDFRxUx
MRWZaun2RHtOsUTA7NBgIS2YaI1WvVzcnCIH9RWqVcLHNkEBvnUV7UiouXu9Q4BnuNoXhuHmPOeG
zuHyqgc6fJE7eXUJFrlOCpxw4ZrZA4SLnZsjs2mFwlnuKUONf/23VHalrgLiNXaM53nFXAht+9qG
TwtjFv1+IRSBNc/AhBk2S9fpMTSfgKlxiGtG1adtA53M87xr7BYlcW6SWvJ9qtignmA0TyCfMb+g
Wpdi19DJziJocoLapPV45jM8GGooUg/ProGO4JAVSsagHgSUyBLCxcytg1FGo7JW5quXP6W7OJFt
trdoOQx8wnyLNDtxYnsbAvk4OjHpY2egQXY3gftDLslnhKz0DdviQXLufUjDqTnDQBroaNx0BnBC
Q/ADMylEfQlXUoOKdisGzlE+vSZcxpwgkq+3M33+bb8eeg4vPrZ+AmY1Ox7eaGFBz7ZzDJMZwi1K
PVHmP9UeyvNXEDeEBAn/e3urkmtjmtT37Dw4oy6F7b0gNHwpap+y/NavXfapfy6r2NdfWCCVIuW7
GSn7fBKvMLC8Orv1zmOFJFY1yFA3+T51uHDqKt9NbpjvyKWMQ0yBWpxTu8G0ov/6bJNB6Lzc2ORH
VwlAuSn4mZCFBhkOVSHTcXRbrKKT4Mq66bCUcQyI/XiPvvy5FC69rVyDUoMe40cmGX8Do2QIlfMQ
6H9fsThqr2hyAf4r/yJyUTd5wTtsk+do99HSA4psyaazu5BJ31jJfY6GR1EBXy97Hxd1NIhd1bZY
kylDyEQIhRNak+sU2l8LGvUMBAgcnCq/NjwqHjOMEBsu1MSO8M4uejAzQSs7chEGi6fFHcwaeic7
+ja19ln0k6wH4L3vPOgzzmphAU/xy2KmcCLcnpJ7MrJApEjVgjNiIYWn/AI6QQSUayYw/DtOR8Ls
sJYbThUX43ipc22aqCBJMtda2VBBWpZ3kxXLEnX1wkzVlDd+hXl6Hoy+9eald6wCvmeMbzlQ3KWF
ZhsFvvIbZJ0wjkavNBvJ/DJGRXfn+vQO0U0i/X8Kry6g+tFvzgAa+HDyVpjSgUmcDjUttTK1dSyk
WacZKSn0xlFngW2vHP58Va/scXk3aQKUf1bNJq4g2vr2v89tuF0RvD51panWWi8Kcu1LRd+mfCGc
q0BRVeU27U7kKPS7uTDtqZJjzB7VhNGNsg6hOh9VTg+qK2t4AhoA1Vk3aWUsNLMOW33Gp3f6NXsi
DwfPy6iJssuplchAIpZ9bbFbcjQcLxdvQVhe4K/SqYBdgemriDCs0xM3psyopB2SN2REkOimvySa
q0GRzblu6IarM+7BAgj0gIY2RCGAuMpIJRbh/Pnx7zL3rdBc8URiam4X+FFjcDNYozIEW9WzElrM
SW6Byl98JsIyrwnutlOPioK4jJ8CTTYzrNZiGQbqg9ip1FM02notGEWuoFgRFDvG+i/c7ktu/J9x
p34oRHigV0Vw/1ZsIoh7HXXLlWTZa/paGVeEJodAWB1gzUh2FiD/A62dSXTvATjgt4jKcAsIeBhE
h5aOVmTyakIiFx+loDrti9fDXwHTvJQHidzTKQQGtbudEFyd0hARRhQsTGSEGNDsubFfTVmDzC3g
1mrDW5qTvvJEFT1FqdZ9J20T69SHIs954+2evQfcXWq/TJEJHNRzh5Vv4FZaKqeQ7PLkhLAlawMV
VTpxNGub+JM96NnT3sUhueBgbSc/b9/hb0wBin4/hdhuWQCJIbFWF9NsAC9Wj6DG0U+38z6Zzd1P
e2ydXIOuOchzJSF4CgSkcrEE/DEYl/ELaGzorVAYpsQgp6R/IVDlcEmCKzeJQk7WxRNoQWD2/Kwk
hAT3P7Zs5EIGSHL76mAyty0Z39pxzETbB6kqYsm3RLW0Av1LgehB7oS1ecWNueWgy9I51wyT0/ig
l7q4IoNlVCLwb4SzblGYud59eqYwr+2tJNKJkSPRQcsEQQnEZdcD1FXVjBrMdEFd2JrFJlkIe8vH
lCQpKDIlOddD4eqfvziMNrlucSfI2Veqez4aWDysEd94L07A6qMSEi2RU75bXgYCSeB5oEvN4QEb
YYUzCVCQPbnuZK5qX9l9AO4CsTl1PltL9dCy4kgs6ER32tLzKf5YAnmhNkTKbLYTaIHAgYWD7qQ7
43R8o196kNuU53f1zqBcrOE1P0Jx+IAnvP7qkolkgwKSo0oBbdeQIl1sxybG+fqjsmZt5lsavGIj
rkE+chC1knaYIoHl7OhnnQPatpr9Pfw5/8tqCX7GWIPG7Hje1i2yNO+0DuOYpIxIIBZ3ztv6yP0t
REp7ZR1IpaemPu2LwTf3x4/kKVaB0HbXcdbNHvU/+fNwSbft2kIuQlo0Cb9iVTcPWhFCAH6m0bxT
5mNtp+5vpqs0VNfbRVeP7z6wk82CzbVxcJ1eZVUM/ElIHjvM0SeQWkhVTn57OODvc1gDsjTuSWUT
HTSZG9WyFLi+lmirnRZV8A3cx3G7dUPIh7nYcfEd0yLDuyAQToEdZpZFXFrykOFWylpTXJz6zLxo
GV/WVj0y+XtqE7LmyoQdMCJ2PZlf5/ceOt00JFBwdUHxzJrWDFJX+d8G0yt4WKOgG18AT/IgkGHn
2qjjrGjD6gFPGX0neQ6ABaGqZkbR7JM5HLRecj4dk3RKQ4eJqeAyGSf42zQAZuNOIpNDf7SeQHzp
E6LyKW1z/15luIpsqaYj4h93BwTtLJAk86WNqYyU4tW/JTnOnI4m9cSxljAf8YmHBptErqsy/NNH
NJ81uo8zfEOWuG6+nE6PIdP/Drh2O4P08k7jlmypF1CXP40pN6GA1WO8117dqnpAQpyLmVyGWZo4
pVCcFX3MFr3rOXpMOhhwe8+irZV6gI7wwP2Wa6BMI/vgVcQ/pwu220c/0q9XXLfRRsVOSeEHO5Cj
qrCPBopgVe3oY1Y1ITKR7cz1iesuvQe/yBnI/hnEIHkxrEr0MceKZqwSDviwh+ugwV3mQSQX047Q
eJEHdgc4v3u1nnd6cJXSzpO324kAheMvKUn8X7jsxOWLA618vE7CFNebizZSo6KYeXGLmvHLpCS9
pNYqmlBTIQvM6R3w3ec+YXy62sf/O5pjAxG5KvQUq4k9aUOunqB20SWHZcaaKiMAYK+RMqVSuyxv
T6Kvldqf42ppKcYQzB81jf5TbM+TaY2mwkjqSLSqAgSpt1WIlKAW6ngcsJl5Hau0Y0remqy7cVRK
zHNv1swVzxUxRlK1WmhAyGv97NxcEK7Dzj7C8v/5fyNo8p2VKp+x1qVH3TdYLW96qC4XB/JG6uAm
mcOcH9bYL2ijjyA5x53yrr49md48xm3/MuQ+WGzZR5u9biqyyBf6zio/w3uCUTg4eM2lecyNFVF2
jpn0xC45VvsNETXK26qLDJUs/4dF9X+uxrnyiYyVGph5C6PPAInz51fLGW4gID40jFMEr1hC4XQQ
75w3TQwYgI+NW0rRNcj4zBvf+oaV3gRExZWH6WS8AaSeL8Ib/Q86A46IBfO+5eXTI3iBfAd4/xuo
GxoRLtrCLMkORUi/W/hsg26cyKU2UurZ7YZgg7VOi6RcXGITIyigkNWdHCSGgLuvdrHD/3hkHaaM
FW8zCqWNP5IS9goALCvwWeZZt5pI9AgBp1TYVvRbggXPnFDvgAnmV9M1EU3qCAMjT+0IqtUSu5uo
UOFjQEiptAeRgvOzB7oDUbgnpSa/dHPAraPgAwLcDqfcHMjxto7b60qZmc45IwOaMPmMkG4yoeZ9
l3/0OqIlI0ksXxZmN4VWcIsgeSp5N3Jxl53q6RrqwpGlczBqYxDsDWF2+iCejqZeoo8bEGoHSV5b
Y152EW5MExeGjIqBkrO9Gg+5wVY1wF/vzOkkJ+zWLoOKj5XP3AWL7VafGFq/7SQK908JqT4oCtnI
lkzZwn9/bwmun1UXYHXPi8xR3oZu5fjoIvVNmb7+l1X3Q0JvEm7dTk41SCJcBOQjrPB5I0qvfi9j
egBeVEflOnfrpWgColezyMbC1m2Qu/Vkr7r72QdKrRx8MA38EE1khCx2tTGSuQP33ginys8mXF7J
PoQRWELvkgRFp0wS6PQjXa513AHYug+mq/9+cOcegHSrUcXAjfTqsnQLVWyG5ZD/LtUM7yOFCoGB
xXgeBN9MWluUuhR1vIBuYHbWbeauv8fiD/xz1KgcjfFWpmYDF4T+MsHfnk2c6P+srCGzVUQ9/f3K
PGHKNcKx8Uk64/1FkUmz0NPO7FH96T4bK6dRQ51LxLt+K5bpp/y7sre1Kue5J0L2TzTIZsbPbXN1
D6hnzUprW7HzNKcisv24RRKKrMFlIIoIlFFZl+e9bAhu8W+IqfK2aZf5r4kyquFbem2PylyMJuiZ
jnKgS8xi0RaQ31ttXGK6OlTANoPyGgXJkDGGFqsV9rYwfWnf33p5YZOtmZ7vhn/atWVBK2wtvM+f
Gw7IRLIWrEts+rgUYZGEEYeAKFWZoM4gpQk6N/EPtK4V6GwH7ufLawEdjdZQ9c9dwxlxD03ig52n
niire+Xv/uXjy6A9tK2B/ohi7dXrnYxPfRmQifOMGZHJTcu5dzCHRkyuUlm48AFwBeIRM7EIks3+
HD6Uq+3dK1ACLhGhegzjTxKdlG8LdpPzbH2zUcZSKtoiW1iljwPPv6szaOG6b1Xoy5e1Is/Rhqlj
s+YZpKjOwQHs8iCuFYkrp80PWnlmZ6f5QGj6BqsWA7HlLex5/8Gbwqc4F5THGdpPL6amXoTNt7+m
AsKyEvpJR9dTm64uSKJrCppuahH1Rn+v27d1aXcEagx6geBesCNWUzmVsruEMmvu/neJ6UjGMXF3
XLwY+ykAlr+C0n4szkj3RIH5zmouGAMKA+ojZAObu+Wf5/OYlE+pPibQ2EEZzYcrNm9mkLL9z9qc
prwkkHrRs+wnL5u4F7/XEaZHU6qZ/yb5ji7FxTbzykfFTK7inRiNrHW4X5ra+GdiyzNV/HIeqY8c
8qll7zZXFGwRTFMKhkAz60GrMYpVftWNMO6yte2EOS6/2TzJv1EWw8XFWTCU03UgZn2SrEwF7j7U
FPh5cDAaHbs8Nh2p1gyJrcGMqjoMde9oMe0ofDXLlCMmQoTK3lLnhAfd01RqHrImlDDiXcrcYAzA
wUWbOtZKSNciDd0DScUUKCOq/Y/BY9f4IzHclddltlC48QmL4bg4fsTrz/Be7DyrIWnMtUtqwmoo
+aKA+LIbz6g+ry82lONtRb2lV1ku6l0t7iO0rj0DIZyEqEUqiSkEUnxbdJdkH1HN3c/dan7IFdNE
SqQnuicaJnmBS8k41Rb/RsEP2lg9RxboiaD0yHaq/dbrJpBPPDRKce4HI8slF5rnAFmfL2lR4YKf
+39ewzEYQJXZL/QfxbR1CS3aaboBu2QW/yn2uMMlP5uo6zlwTDKr66oAt2JxIgMi6pGUPm3blr3V
iAmZC2zWG0eSFeK26JpT3ZFlMmdICIpzMLUwXpXmrhUFDs8IjJpvwtfUtWFwgVjfEj00ULZV+GVG
MmH6qvIgXlTeE2k+jRl+RfQzqgBI5KVweAhmr7gsJz5MojZtSpw/iZtxlJZVU02c7XMxqaqeFli0
sh88ENJ7L2/AuPs+GPmEZk29Ft+bIPtvFst+RLtC+XA8K14ncfRKkrnFMh6g+yeMRKzrJ/+npFDX
DM8NMAZIElWp/17iUf7jsDFhIQkbM4h5usNO05o7c0Ivx2aZ2w2CX1pFqRJXySMpaBdZYsw2qr4f
1glEVixegbBRnkKxiFUI12VmsV6EFb9KbQrwxFSOHCp540D1plSGJJHV/Q/nnzMhI30EoHudPQXc
C1TIGkMHazCXgdCSoYQ/783kgFe9yRbO3Hv6+wW6n49etgnPh+cBxJANxVT6iwF/qgWDutZhIeCg
CsiOkcLPqyM5cknGhXxv9uvg/e5NUgtvk7EbQLRPiS/8cKqXoI+Sg1Sz6Rlqdsi3VUSikhahbJ4g
tzn3Hoc46MwrSTHRdW/XSe5JjS64AJ2hmRtwNjkZ+1UFPuNQiinem1RUt1ab56Nj6C45GH5jhhRm
QfxWpV+nXzdl9YmYKwUKNNT7lXZQITEHNACj+muf+c0jZAZVc+3T/fVLuq3AWJ890gxa2ge/sXcG
nUuUmktVO9NKtmV1FOGp1HTIiIS1smNU9/TMXURUSGXF+6fEvxJOU+8stGxJNx2Iw9Aw+4lB6mBj
F4WSereTKQNSEfGmp8RA0EGN3pRwNVcuDb4GzAzFcp+Ut7CzhOE60DCw+ydY3OhGbeCSQM32+kM6
uBX/VYaRH75FcyV9pQ2LhRE1NGePG3oWvbkitvE/jorlXUkczHGUoyERJgTD9xlStZSanJd6vopi
JO5NSQS+benyDsn7AWmGSYftPoazdJ3d+T4j2YnwwyIek7Rq2zfp8Sfjk9BIPxphUX5GmVhwanYs
FwmXA3NHgrQ6QHyTEcKESrNlHrkk+nuDZKvgYO3F6qWdXK8PpEuUKNeTCUlqzvJB6POkUCp7UcMY
Y4CnDvSZDhAAbxsbhgv6LsECtbjPm6AMumwNEQf6oUjCB2QniuaSU2CqjnqMd0j6CinbFdrPB9N3
RNwucO1twWdW/QuwlsNit/RHjcPNLUcuxg71Gq8qUYvTI+JjKClABm5eSPfZkqLqZ/AQOy8Gp72X
8inXhPPXAB0PxWpZz+HZRmyqVQMu8gUxiV78t3Xy32Z3XZWWOE29ICxccCsYvV6uTp3sgv+faemv
cxutFsk8ZrMNUURMPG1Cqo8adBLjYmOfBpraFECYO0Xbusj3FEtu003/Z5cItoHIRrbKXo+0zAbd
3c2a7hAil8NQCfyE5BE/rlj3rp8lsYcx8jPiLleakc/cSFXO8EqllRCzoYxv/2BKghXhyJU70JZY
zb2xHXpeMvKoNbpL2PzK3e1Fo7pZBzT4xGb+kTwUlrv3/CZ/MBKBfic/CGuOhzhK2as+2itaStfO
80duRuxLeEC+8KbOnLQftPxNhU2sIiEOR2LV352bo5GRJD0fvPub9F4lk9aRjTkd+rwpLYqh8Qk+
QmBAxRWRXQojbvmnY3QmylxKtUoD5HVTpiYTfXcQ7Wz+GXtefd3IWCJH2GLPyii4deWJ/Lmvc5cL
2zBliOwLXROEhbWwpdNx2DvhjMAOgUW8fNueD09NUuyJUH9gFErM/LumlICu5cPihzXfS8XIl3rI
NUbgvlh7H8ZxL2j+V8u3jAL+byL00p+Pt6sIaD2fSiM0woQq+z+oRfBib9P4bLAINJMUsYBKlqjl
HOGvHeA6lKxa8bm3CnB7sjh+gu3rHzsmxZCNo/bctY0u0SuhmdOlVMt1qQmBRKSSMiCeIroBsHSW
nEmGCfhPXN0xIS59SzyMVpPCIqDzJFCMb4tIyzeiMfTy5m+DnNdbdVixWkPpU3lBXW7toJHmRH33
GtaWrauyWfEjLLp1qiFM29GlpK8I0jnsY5p91BTSrxKp3GBu2N8TxnSfNYDyBGdyhdMMeXQOI8S+
qefU4aQFlei+fGH4CPTZuXGkScDyCsPIKJ+gfBewzyhfexu8bUZAxsCdxwmV5rxdlGBjXCnA27U9
TlaheRSVpbBpLp+2nO39SlDtP6LQErdAY+BMJwACQp/bN4vkTJMriIhZ78PxcO85CCEClBX21N99
Yp+XBjcSFuAVcrpodjv3wS3mX0YJReF1Z85uZsVrHMJ82A+xr4gGN5cfO1FnmaAHVjfyi+7+QEIb
2W38CV2dn4cUTZ/ctHCZosc75ud7aCAbCpQvjOgvD+NrbSa7mQMipyLhC6/co7hP45HCUknu9NaW
hpfBesjdThfp4akezux78H46SQ4rbuUIe2JQ++CIQDAcfyRLQ0BVEMdHLxxQFAcuvDNPFul958en
HtJZdBgxDZbRyVSEFmnm/POMTRR55ry+kORI6SaMPN58fL6QTXXKj0Mn2MBz5CGJmuIh3PNhAsGP
lKtxFXzmbmV5JuoghjC+GKWJbrInr4gEzomUy30jY8Jubmt/D+87CkI9buEsa5OJFdm69qFXegn5
5LXocMrIs0YVkuc4bFa0LGJyV2+xZ5MIiiq6mBJWMJiasz74vjWQhAhtxw7eL//VSmi0xzRw0PpN
3OjBmPYwnPjLmYsOFZiueQ2g0UdbD4OaLyrYe/MP/UJ/aUEQEhD6z7iHJ+GyhiwXfniVzqd7udqg
Eou0EvQRMTtApoU9f+2n4tMuLA1kT5uePoSHGbnlWQcfclxGBUK+RCtq0Ran0XWQwlL95Fh/1KUy
XMvTqfEdLaG5fXiF0B8g/CbZSpR2AJxEvr670HUmyzv68uCKiVh/KlB3QNtiLKtuydndMVIRr3v0
Yk5qYSaC91Mn9FBGnCXhTw6U2dpmL34ReEhk2CjN0xmvu1Uwb86jisPvJvGu3Qug/HwAYePROVO9
3CqiBgoktSvpO1qp3iV3SLXyQOYfXTJV7FmbXnOyS6ppJnLqtZoXbmZLIPTDtxcaHRo68UTvBP6s
oNSiZlYzbAWNOV/4ki39wirRTcKIe01wRAxa14fX1e5+Lra/naAVtcs70NTH2DhxDJBvGOHD04Ji
g86w4wJBsuIddGLrM/yq2iK2usZkrlJI9VbDT5IrP5Daj/TBxa/5eoVP+swWHpwnIr5DYjb/16Hh
DKtm2+hhslTUej54oDIdeFiZWz+4+KuW2G3d+8kzz0r88vvuKdTuy5vM25xpvtJ71HZVYSP4Bc3b
TSWDgkWD1w0KrAixwsug/T6osEDqhJlfFstF2DRlnaqTWf/Zc/cOSln+kXKrYCDFn0r6+bYqwWQa
ZgI0JCmq5SExaTQuTbos03in87xRfUqzvrQUUsqHLFTvGzgpZ6it12ca52s8aSxmZg9dJd6LlkJ+
KKxDYVmrPRYXXizn0HvuAWqFBioLDSKIYke99L0wqo0cLwTyfgWRkx0xNAeecnP1fJTHavxeuBYJ
jXsi/SYh/dcTBnLyssk7g/SK0cZ9/JIsoEq+l4Zq8OMQAAbqgja6ErRhXgOMqNwO67uJ/N7REBUi
F5NVSTTMfa0mHGpFHbn3tu5warWp211l15n1YwLrI3eub4pNS4L+kXFmKI4TcaQiDc5G+DMT4uGp
Gq5c4kVIOuqPuzR2nRYa5hhVYUohqTc6EDPPzfuKOLW92L8LkW+rpVwNyhRytSojGpHE15FgXWtn
S6t0kZfKQpdRSwBayssF8ocx7MHAk6DLgvgxUDbvNw6fJcwMBJbHFmh2eQJhaPI9afSEl0ymnRIp
3Bq7B5OYbr7ih1FPBZiYlx0/nOm1A2evQzK9jppndCdvp3UrJxQRh6MUmTYs/cQ58Jy7CqIV/BBi
Hyhe8q7D2BC/u2OOD/oy0zYk5PejTmlA9QFc8NFpDUA4mUIEioGVxCmqQCerQGA7H58/JriQYTFY
CyFgnxjTLXwisJT8oemWSr8bzy5JN8iLypJ9vZsQp231h0WCyqF7RKurk4wNNZTPZ5ZlLxNvyPak
M0ODYavRhCrxAvIgCprhIkuSHeZE0UCeIyI7SO1Agd4XF6kYTBq00h5Xvt0ck56kk5roj0i8CTBn
eTVcCTUKVIBe6xjhYlKcSLPbsvBXoJRbPma0IN8FQB6849WxTSS9cXJ+cQPYM+DiDlXY6/5asr4A
+XLK1TlLAr3iw/8skd1xkz+4R0nxxsCfUEgjFIsjuHGLxVm7tVEz/Ut5pElR5SehcafekF4ieJNd
YVIEmTixt98R1dphZ/lzElbTm0O17R3JuOBf6Q883G991W4jmAYUrWeIsWfVizlP6m/Ac9RIdJBu
9fwKLjcap/5BFvlf036O6mwapVe0mXglG0rDBrYUPP4gzHMpMhEERuKZvAOScKjoGT1chfz5KYUV
HuIELzPTqlVtim1mUeJLipQtbHcKwUBXvc+B7BRRQ3gbAbtpOZRY74FE7gKiQce77nNj6/voE+vq
s6hFEymPAMfoTDwqeTZd2eo45obmDCaSIG63Aouar3RA1E1UDZ6T7OufUn3JXItCZQsu6cBVazZ1
5vw/QkglBgMxliD8nmy/1wmMwndUcIP/6GAOPFBMcAE3JL4SNGvkJi2ao1bUpgnTniXcezrR6Jlh
rlBE96S5W9W4fhmvOx6rABvrT4GB0elu11RyqlD3RDJYnOwLX2GzxTWH4+P6KU/XN/2CypntmAdy
agsdXM8aQhlKS/f72fhNimursVt5gMg1g1vwPvKii2m7B5MwacXE/IRpmiE6/fvm94Rsa5pyrwKL
+3vpuT5rtGwPzoPap7aFYY4cqvmhzos0XZ0uFKsOloykyCjrXurgA4AsXuT/ZFIY7ICslk8CvcaQ
pJSJdgd0Hx4Dar/2A5oXMzTCynfNUqAOOAdun2SV1QjltGsnemwLITkpXhNEobgZytWJTXVGl+n9
jfVaYdJyGQ6rslrOZVXXe2jXLQRJxnpWZPxtO3tb8fh4t5t1S4OAsdqLQtUtZSSgvRM3oobwEj4u
vpur2Bi0oGn2sgUNdWb5+M54Q5+RF2y2Y7M1SCIPaGOhhrf4goVyRypHMRmNsjNwT/sKaHFAuM62
sSaCSMzXF70mDRZ9m07gazG2+s/p7pziYS/FM8WvmqvLjfZVAtWnIUIt2SbhhyTplBHhs54l5a+y
lK2U7hqIqDUCAamZVK2lUFvvpknwnGwTd52Zv0MYBnVvjNatEBGIQgB9sTiTar9DLs81UDMns5Qa
+s2Qcoj+frtwCfhKpblR3MpwS7NQ5QSntPMMvjDclMKMnlynFzhOaNofM/S/XLgCag74ECsiMdOi
ERdWpIR8ZvLgZLqy0Devwv6ZaeIQ9fR5A55wcY/yIlmah4bulooPfCFZBrtIAn6NEHhUyfVsU/Fu
0loXqxHT189+urJxeir/YgYYoYUIueAAQ82EX4fOWySeUld3nkSF/rtj7xlYuuZGBNCW51kcf2ub
mmLwTAode/2k+F9whxXLa4JA+DM77CFt9MxqTVBYafedhh7BgLSegZM56SCqIgAVBPmZJp8pPJyj
zCLrTx3FBSP59hm2jBoYZqu/pdvwf4iLQcrk3Ixr78cB1FSnOhxxrZfDKXrqlmRXJevJ0ZFhNPbR
1UtInJrLNoyqeZC5vSQsK5C9ZTmAT2KGkZ64VnDI+YJ57g65IqwNSu50bjPZkd9jYEUy2j+Uoeyp
BMXCU+qVcOaJRMNMkNrIqIPa7ZR6V5c25AngnVTz5sO5i3YWGfM+Ncyo3MOeEHJBnSqwOZD0mmU3
X2XBHdKrFmrdaM/PyygPQipA1dD0Zv909+CCzOKpJVqmRcqdAsfFKTH2p01uk7W21RKlEYapvMyR
BY3Mw48aM+k/bncq1BKAQteyFqrUGWlbuKCQVEaDI70rmFwO0H5UZjt8IoXabBn8/WUaHJhbVNlZ
ZEIO5s6/ZOfTV3N8xdoNBPFq1FYyUYTstT7gd6fy077OrBme06Sspcv4oV7TUXt+7knDHoWzhVYT
fpYumDRThSTnF7jByS3nwg0COSp0hylL1yF9aDn8UO8o5G092bOrB5EhIrxaz7gmqh1TPc7syYTg
GUDMHOjRoex5fb2+P5+XZE+R9wzZ8CTiJg560MxYtvQm/GxdmA9OSKTBJ5Y4m5GlIX0ncRGaxvvL
t6ksrmNP+n0/MDP9uvj8DmainvdwR1Ulp85PVHjAjLYngmwC/JUd2cT/X44OHdBbGJxQpo2ElAPq
36ycSvi3lavldM02hVfz1UiO8uhGl/cRCbZhRktbtwUFElShPEAszJZapu2aXkasVQz6KyJqd7VN
GcWV589UZu/1B76rdfZpkGvp8MwRha0xXvcQz4nUQWsqeoeIoKXZYvXkV4E1ReP+UnjKzz5ZN4H5
gYnYxAwK5wC1wsptzECUXGYYI8KxLqqOSJwDzdajBBvQ4hAMGQk8UBs1AQDYLSquPokCjM/BH1W9
R7ihInupfQudj/7POtm78xmRYpyx4gh8uCIcv4fQ3anIzJ+/cjz9OgrgGMAArImJ/MG52CRGh5dv
QFG9woL1pz0J3fBJCtN6zc6Dw9VjjRFd7dD/JVddEJlJwSvz2UQ77F6XJ6ccgVFgR0lHVnaFZZKp
ajQnB5+uTdM0JDm100/vuAJQYML/PccoqUXN7saTMtMA+ZRMCP7OTgY82BlfMJ3cdVlXJLq2WufB
5RVisrupIFra2SFAuDaGRvhaRILsoJHLtHLwyE6c58cvOQdDs0Posw28Hob/doi8pMHUpTMBFYv4
MHQQBzOrEWCJMQ0GnCyH6+A9ARoCO+cDcJEX34uGWKjv6nGkB496GNqZivAu+o89KL1ZvfY5CFm6
Hqh3expEPExSNT5lypHu/+lOnQo8eQ6XHoBLH3gwFAu+kSGUMiB2j33OC7YSnGwxk9WF7ytcYFmA
gQlFE8cglY0mRCeU8ExtWE3zo5eAxPUf0wnOqDx1XkFphWx60ORRx9CFuQYdPuZ4MwMvJ68OkOk4
BsnE9FZFd0E6587yMLGJBHzJxOlTM5eFVPYCRaDy7qy7pj7iP3pjBQLxqGaGsSu7ROFivbZSnjH3
X1XdhqAfwZHUConBT/B9lFm9chOES7NDcyvBzS0zop9ghXpFPIMoYIgDXOQX2i4874wIa/eFbjWP
pduZaR3h96xmAbZz4B+XFUMGJV5DtLf3luowouvwQQaR+sZTZtiWtuj8HUg2xLYNV+qW6ugOHgox
VNKMYkfxhM13t0pgqr47+rRqU9piBL+fPlEiudjgfYMkY+silVl/HPZsKlBUO4E0DSGOyVo9x8KL
sDMfb0U2RN4kBPP0BL/GG+x3vjGr15ZhTK9F5B+b2IfAuXe9umapusqDQL4QatKExShBaWE39vCK
51PZm4zyfjh4bYvDxt9lxzx3LwsyNZRevTFd17HwFmJqwQC8f68JzLbfI6L86NAGLRmJeXYMgm6S
0389OGOaLaBD9wS1iEvEPVaGC/IFUW21L202b/Na9H6BI4ALH/3VVdGtNzV0CxLrwU4cbxdap0uP
qepBPX4mfgk3syxmDeDYCXCxgixhKVXf58PjvCa6a3GEvgG/kmj9XpVbVuZUKcr1NZcVOWrYCZx3
NfVvsBfRdjM583Rcfphe3dGg81HL87Cr+Svd+xCYgA4Vz4ds+zEAyxCsKT70z1pnBBn+MRhkwrgs
47J4COWXuQdwmBQtN1JZk2245arCaljGPqc3pkc+QVFJrHNhkYx67LJFWmqhNF3EkjPn6MQNbG2f
PLO3RRAC7eJZSb+dWUG5gy56XYfnksB32SGwPLcU80UjLojXGoGodAjvfI3XKLxDVg6SiFgjVGPJ
DrYUowmeVYyYAwA+vSpCoEYCGuG0d1gLsOlqYBC82wz1hExdKUXQengv6eno7kcUY1thU7vUAHs8
f6hE6HOw42u1yZoGkL6ZAuRNlEmCaqUyyPhJS8PAfK2Z7kK9GmqrFZoIoEb/MWOYTsC4m1HnLZ4a
QtlieDBT0R4U7Q00U5b8NhFSdm7edfv6ra6eJ2YcYJX+i2YrC7tdZocKMhrAIvbSeUuFbW/Qv6lA
n0I3p1hVgrsMwPhd7ptPm/LPhTd0cvf2aKvZ5+fimsdUi6rFnXMXAs/JTTLQhjLh3jW+odrn5m0D
DKpZxyLBnCbBGVcz6f/4Hgr4IIf5ieL3Ak5YVKiEvoPj/LxnLdZkFtyzU4hRdw8T+jkunMPWFF/+
4uBkswWNr6WawwyyzS7YHGbyeHx6I2zxUPyYlbreZhyUc6dmoNVCX7FIm5GnQviT9+prNn8ZRh5s
M173wTL7hD83PYlXAFFBgv1lbfWkzNT8YndQ2jS32PgZBk8p+F8Grl4IsRryUVkkJXwnPDPHntrO
4ZLqhskg3YRz3EcyDEEUda/yAjSvkZOIYaFgJVslQ3p+nBep79mc4AQ7t0NvXuM3f//WAFQGL6gk
+4f9q5M59yM4JByj+XxTRwzWEWWA0Kx1nOxOw3qOxFtAsbkuuqrP7VtzUfoACV2mJiN75XJdUpbO
10+XNJaRmfGZcQzuw6p+DDxCmQtSm6UlnwfKOqT74tCoIZrdFlKtwiaD8qoCnXodOy5QBBDmJ/Q6
euJoSoSPvMkI6LnJqmVm/co8Po5AatDJ1Wstny+yQt5BPI0mNyh1HFQbokNFi3XQ28JcpSFIKiO1
frdROZu3hrnvQWx8CqNlCFgumtGUSpVSn43Vf+CpG7p7tvE/tcXh54GVUeXiyOdhi6Xffct4RV9A
W+5FYuDZzd8wWto/OSvugbWZ3EjfHqZT3yin4rFLrWMFU5NMOq2F+OjEQREzxomYGFbdZzp2hYEO
H8CUChP2RGU2JzcIx0WQGJBWr4DXILra/0BiSlFsU8mT0tuAU4O9tC31C4WEtZV50G3nEBYeCBWn
Jzb/dQzqza48vc2u/KnH+5PVOZT8N0sY59/u2ogPzVB7dBjkgpm+1HkQR4kXSEu1WlfSXAE7wMlD
kjIfLHufMK0QsIwsVqNgR19fOgajPrYjFMcdR5FeVFJ6eLFma+FJav2rPVo76jXzG0Po6x6oVZJy
6GwBWMFgXR6fpuu5f48uJVWLOSJIXsQeNURBfyNXrbXiNl56bLa6HS5URXddyHorWoxOiAKp8hVG
9ZU8qYSy5WT/m+74WJ17AOOEHmt2yPUWVHHzTy4sN1eh/dOrwzoVO+3GW78/px3vJOWVQQijmNSG
omgreWkuvuJw2EdP+vB3UX99yzem9Ke1zN1JvZbnJrGwka28ZkqfZdAqmlxpO6zKumJaQOhHDow9
WHqpjLRkUdzgRAFMQyMPhBLGYRUYimfmR7zoGLclskq4mPvhOccvV9A8KPtSg8+JYE6O1ZcGdz16
fn/rzMpviYyPNXjCjGvLtZo6fc2SBSiirvZlKL21p1Js7qSlx8458HVuUkMT9972t6iGzZI5L+o5
MY2H1+Qbe/w1tNYObhqlck4Olh1m1eb+/bR8CB43O5/DObXzFabsiSh+EypGO6Uq99NNNWy9/iKb
LhXLOpBbm9BiLOf6ZoS5+fydxfJ4No07+j0zCuaYiqDkKMlBchjwRPi8QKGnq48bXGdhTHr+Dvod
drusAD8PFEVOlhgZyKFb+SkWfdWmzcVmfqMEqLfxoZT0GRZdXoXhRcNsC40XVZRenIBDVY4d13L8
ZMdP3cDz1+UOf5CaFoMTiB+ik75DIC7iZrN3Z7cL6HLBVo1nPjkt7m9PVJwbP9HyKfJd8bwLTRi6
BTIOZEMcaYijZ7F3V2jpZPuaaT7nwOhRTZxCNIEzHiSQtf4SBEJBKC5B6K+m25O9/i0ce+9Mwd2K
qejNXsp0RDnJR3bjg/L9X8pL8AVhXW2/AH83vr84F6xqBJ2P8FQkW3xk8gvOMAjZxZiePIqiB5Ye
o2gtqpk+HUgEpLwOjLanqBtM33UWZPIbwZg60x66qSkLjjJ3TkuKxt7V2p123+4f1UaPv93FSY7f
xcetaaGAH7jzSznoBFWLe8Z3VSmJetQgWVUvbELsepnTxV46e+MdgYcarNtAtSfe/0Re0o31JUtm
mkt0/o4xKrCISeDkZGKDKg7katC3PF30y2p0KSsf/QdQq9N+sDb939OW0d/WHy0oaNgSWQZecJT1
ZdpRyNts5Yq1iG6EyluP/6EDMczldl60uuKgIZtA51yWfg3SGA2KncUyCeJXlwA5POo3yF40fz2H
8exPIQwdvkKA+CVL2UM0KdMgdEJz0SoAmZm0x1eVikOqjzR8Fz5crbQ3h88orAPRnZzfJ6HhFrKF
JQVuIrqNnWzvG/7StbsyR1BHNLY7knNaR4snx360zBSW/IF2+Wn61Cp8pLSmAZJ7j6c3VlK1aMMU
eysfQ/GcxD6+6JBchJhlsC4GYElcVa+g31gRNB/pIWByiq/PgAQuHU3DE2Xvhv8bXEmhO1iw2Mgh
sKov8qv0875J0RglRXG6Qt0hV6mURpTAac5v853i1Ed+bZZSMbA0Pj/1Ng6yJqRsX0DK5ETAlNga
fl3adGpGm6qx5Oltqewe4AGfASLyWGAJUUtjboQsZ42VVi8OZ9xFNJYu1ZlW/wRomK1lqH0cs/xl
pPMExJf/QRSP95FW8Vt2e5PaNvXdMZ4h1ssMjAAJ26aNt1zANKiiXoaNo2bucIRUFquEZ9qHcoGg
x4pu0FO0Yammnx45jp5aEJvX6HOYb7D19grCgfD8mDOKZEvBfe0ANXNgTX243mtNjhAacaMyJ3cU
md2hk9zDS8j8jIR8u+WP6e83lYVmGvRBQsQOyT9N0hn83wOsbO+hmHjnAp+YjfqyhbxRdkUJ4Xp7
gjX2POE5F28l3oNdzHxr2npj+PUFXeHGAcR0BnLPlxJ9F4BK+pe1c7uoY9aDS3lmkp4rmk9gPn/S
+6AetbIc31HN7JNUaJCzqto1ZdKYgATLB9Ls8iZmxsPaEwYA/ipjjrvyQBP4lyim8c6oaFKVhYUu
bALp33Xik8aRCyRWu81eEJ7JhXNBAH4Uq+Uha4AhoBdAAzkQoNNkd5CbMNOjPG9bVO2FjavAC5R1
enhAjvYWKcguMhas7eLrTkBu84FbxpAkUzJMMXezW0EmXp5vo1MD8gOsqEXor2iso4uV8CsZBl/N
GKlDWxJAJJu2gWtUKgfchQO3L8aod5SOp/EmxDUwM4tCZ6okqQun+y1fSoWv6sDZcHB+6fs2ychu
tGQpYx5u3PqqAUYQcS7Pw4E0YresBommCjRZGd0jZ4qYQBmUzd/MsOUUQ5RfzcPSqhiTltxro/mo
bQllRIIrHG7ZoEz5d5AX/HFcHTBq7DtUws+E2oTBOKzw+WKGEh9L603MC922jmJxQaxunjkGw8xw
PqAAHtSqm3WwkeNWiL2ratd/fPjFB6Hpi9H+6S10M6JmGeCe3xzhNkStTn4cYE8k8OdjsobKJ6f5
5D1XCJNXWe+ogHk90pnp248Iecf60R1xrDQTmLULPRcJpZdd7+JGonotldwRqXk6bdd80X+UDI9/
Gb+7S+tx3mDkMcm8q7ycBDhtya9m9Xu9QZzXxDVR9D4VyndcTdQWYlZmYuAJwlCXLK2Im1jvcyT0
RQw44m0Gvl0jewSFk0Z1H8szML1fgMCUS1bwI+HScV+uAtoBBb8TpG+8rxonwNkwUrpy8chERMKe
lC0yMZvyTv2B6Dj9C8UBgKZ2wvET+TSjHJ/m6AIREVUp3atyj6A8aXefp2RfdU0zj3g/Hsu9o0Gh
4xAMNuqaNXwT+bnjDp5n4GHVc/el3ydW39+TvhNiMQPM/eB+e8QCF9HAX0S6TRUk6dKT4bZ3yozk
oRLKs9hP9ftQld7V1BcLKePSAxa9xFl/YPT1VruN3GfciXAsdYldkto40mea0/QudEbWlbU//q+e
Xntnu5YCUW0R0wIpKiieXRMk3QtbQnGnO+8fYKwigfN34ptcjRBACYAlocdiatITSZToMlg6qApT
Wm3CEIJP2dPe7x+Tw3SzfNpLaR4xuR7yDastiA60MtfLyqxK350k7NL119mDsdEx+Bw74uW4jwKu
5XnxvFDfQK+itE9kOimvRLc7sa6eA1KnS64jneYogqwcF0pf9fg8MOBMeZYmhlZGpWWuNHVo7Djw
byIXgms1lWmxxVfqqjYqJwYNVxppUTSG+RV/rxYnvZFTsPk69zkVUgBxRrpzUxRWIBbn/mXDrJ/c
KZlIcref249WTqgQLoDtSwjoheQWBuYQMxpwfrGEuVKGhvWnzrGxTePwZ7QXOq2wFTg1zkEt+Z0t
UVU7oGzUW2WswcHvTkZiOFQysp4IUlmihWK/anze7QHYIIaSP1FuDv5EK9DtBpuIiFFn1zp6pdqN
5sAX9WkWvVUevaevRc9XHampdz1s1cjhXJnbPrC4fjnrKvUDq8cz1nDwyQ+tOrr079kxpK/y6mFz
f1E2wqWSRg86HZJY+ywzUwY2cta0WSjF7S8vXCJlm06UrmulPRjp0TacSPqLtpuZMb2XVhqzPtT/
rrjhLuv6MFX2QoJojJrTchH7dgSBZ5Zb8uP/5/CQfUK417QV6kLsq6Eh7KlecLvLNjutC5Ht8SGh
Nb8hlZgWiDdJGON3667uuFSK1nt3zImchCSf1k1MIemn0uRWhYnVCxYYSV6JV//o6KwNGEX4Sv1l
guBotA2SA/J46Px3DKEeHpkTgpkuspE8O44IWOVunzCFNH3gsb6gCj6awyYgeCbvZ8zYWz9rSo+G
8u61ZWJv+vfreElUPD5aTndmyHDVbpEMqnZZFC9oRlwrc5L+9o1yrF5rqeF0RBOlZ0szIC56hA59
NR21QzzknmrxCSFXx/SoP2Q2jW5Xp4uN9ndEek2zZtxc9MurftCk6nl8SiWYrZaLWT1Chx83TaB5
r2SmGm3kClW7vml9gWQ/LOk9isKxGKZJ2p2FTBTOUyN/xXne7LeKm8tQpTYWNsLzp7cwVoafq5E/
Ks92Cn2/u1Hc6qavCWFdykBEhxHP0omnUkE0n2B/Hov9TMJxLj2C08P+2wUWmZdNmhWT4oqaIN50
6G9fnZJ1izbV0mgcqbbGNrWZubMmEi2uGdnp6or42yyRNbGyo89tZC/GCAinDQyfix5ltaXRmDr5
Gb79E33J8O7P4VdMVQHcvVrbeezMvIgKx3+xPUhQxXypLuPVZ3C2R12CJIYQvETDtaJSZ5HcgtPy
HRBNDE8XIDPVpIsMl5pnnWrka3YiQd/vn+hMCdk0FROdCpTOXrhjN3kPV2i9NfgRzMtbkjQTxx3X
gHccHEkkHEkxBS5XRPkTgp9e+4YhCR6/f8GuYUUPoDdc/92VRl4sIJwwR0KkJDBe6U5h+o42FUOE
gSvxiymREJMkCGrcmCeMNSllkn10soVbnzf39nu7Dwq96LCSoTuDRA1JoL63Q60wHnvnweS64tdJ
BNLjappZZG2VuptD6dEWD7W3TNSaqR2LfDZcvIB42hBBsWxwmwzYC4FNbWAKsf7Y2apzXubWuUJq
Y26bhwgDhhoqhMpG7Mw+BhOPl3v6h0YKXbIalTPw3t9deARCPIBSG2ce9v0KzYpk9bZxt5Qsb65Z
pl/DFBLXes/rtEFidQh6qJGF4c4viN7vtIFosS+ISiNsHABLrdy2ct0e/CEZq8IdCxAFm8vqAWVA
WC85x5rgTvfnbG/ZOhQRfDA+z9PFT1gcurM3OJVAFNC4EC8iYSiEkOG9TH/X77tKKDvC9w7Ut7dx
0JdTsIzEeA8cFXV6slRti5BQcsZs0U5vEITL5LtSbUDjRHz1AyxYBaKwJu8nY7ewMIHK2LAAEGIx
0toDzfclT8nXrXD5cFzNJ9uIW3hbL5YcWdBpr+CsHMvdTsvSFzI/TXOrYbDv7zcJadBoV+zSnKUQ
tWHrM0N7rNftllXyKK50IRPgfc2NzHSeEwrjEYhWx+9//W1JgWeLi3bJopssIL3K3K9FszR2W52X
xd0E7dewJY5TxfkD7AIRyrSeVp0QxcYm40ouDxtJalNP3ktbRngePchdV/QFSbxpbZGad9pOP5fH
qXVSkS45qzrRFOIIDGntpSZEVxL/vsUIrtPGp/OPepN4CsZjViz6PKduDF+pgI2PDm8QR5GKSO/c
MHj3WvMHL8QLYb4seNW+dkJKjfcO+1WXr8c2MXo16XA8+jLcGtoU7Xf1kfUGNT48lp7ptaZVeOYP
8aInYQA6Ny6cJSBMKdxWzyizITkapR3T6OfuB15p/BMmI4pMn67NbuT7ipDfq5EgL6lpoFVUffae
o5PUTOpXJ0+KcX6u04AP6UoRD6lNvySQa+ZtSH/DJ8ZMUh6S+Z1W8diqs8xHlYNS7A5tQP7mXoCk
wbEWnbHbtI0A0fSeKc4GnZJVfS44rIfsZI6hIidNvUdb0HhpKe41ya/It3iX0onOejiIJoNJmymO
/qSJyLzaZaM1EQtKhEB2ajBKOsiRx1tZYNKaINSTfF+Z0hTddyc6bfQEcpfBLwCkueUqtS48DVaq
ctW0kxFTSq6mHWPrgHVP7WyuUicQmVs4xe61HgBfjkemr4VGMU0Y5I0FpZIadekiYBFCU2bBf9AU
t/Z96Kz9HCON+rh31yCXSUvHT6dRy0ZR0fa33v0alnGQRkcTKC2TAjRXc/GlW+PC+OBmmzzmQxyr
St2CCLaVnJzgMX0uN2Fl0awrJg4YfZh0riW0MN0KMfWonK6N0DjkD+4awaB/khlYP8Egvgha33/3
aCG6WMswd3XEESP6EomxL8MJFWn0zFS2JsjKJyx0UEWPq/m1cb0SgWxcD7E79jWLKXb3Q2p/1cwg
bmZehmC5M3ZKK5w4fn4sdUkqGztULoe01SRhMtAxiE9H276oHCkcKfQYAf3wT1656gdm9OI2ErtE
ZwUuN6N1uzr7Ozq8/yW7+7d5nFMO2eop3lTTLidZub5jAtbX2o/6d1sTS1lsYYkOCtQLWdpLWPe4
rKiq8yzm2XhiPyeN4Q2ZMW49KqLsV1tj0YfgreYxIF+XogUv2L6Xh+Z/0Xc9cInU6EUaZbQjX6tJ
gHBIqwpvraQv5aMcSKvaNUlqdGZyh7fZRdfIDwQGB2Ph1WyU/eZ7j9tLA/La0A50e4FEd/a68wGd
LBKqLAVnVF/v4uZ6ZmQPic0K7KqGRopefbcuUVmGggLGCt9i4KVQMkEcKnb9dk1HxDJGlEKTDh1i
Y+cE+TZtczL5NkPokbKDl7pRI66wzc7rYKIZo524JNF7Ddd6Rf320EGMRbAUQMSxuJmyKl1By05i
tAfGSD/Iro4kDIpwJCwBk6YaRBhy8FYkuBl+ZTDp/5tyefbH4l61upKrgUDvJ1HReUYGFUTIULS8
IJ6DkwAXzukJjF9l0ecXCC58f8O//khjpi1rrEVsOIVPAwqbL85SSFwChKc/Iwd5bne03KkgrPrx
ACGK6OsY0zvKC+pWyQn7G45+PpKgcWF5oSfZf4VN3tav4BtWKXzEhNkD2byYsm25Uz8tk1rsSqsj
22vXFnvKI2f9rjBLOOx/4tz/Gj4hHsmKrRucZ3ANe+SNJ/PjO0plFI5p0EzB91KjW6q3WuX27j9t
pYsBShM2VLmyLNFNl5e8YRx70LyoL/+qoEcStYPzhVSwrGl61kp87Am4sMWqsxfsJGOK4zEuoi40
lNZHqIuOB5CeGWliqEwH8Esf30DiFvav2DADHUuEbZBO4hEjM3ODRgdyAHjHqRZkQyLVCIdZTEa1
3Dx0VaLvbYM/1hR9x+GGPZp/hTytKwpklyT1A8hGuL1DEkWNnSp2UhZ+0Z5V4hH9kainU5Yi1veZ
l6ZtwWQSiLeAL1Y9/rXsrOte7oX/vzU0ALldqZKDzK+Oo/Yn5Y0SJSFitm9Cq+sGPEocauhUKR60
agqnFAmlKTMvIwjvP05ins6wT5DbnzbZiF+3Nik5plPGs/HgOkiTEnrJeyoAFwGu6CXSy6G1emPx
NxP1FRAtZYMEWFhNLnPPJOtxAH2hTs12Z6AOxcKEWInMOAmdttFv2rIzavEkzDrMAh2iw74vNYJJ
e094y6vL6tazMwD2n61pU5oJzgUQXCL74f4IUFue82VJC1ZU0uj2VrfC3OC+yDouwDgBG80CME/N
E0IZdM27mtPQGcr0bnUd/C7GISQhlAnFoiYIOKv0Y+ebj7zewY8doKrBPVThSUeAWKEoq4NRjE0I
l/9lywFYXWwvVedEcPUkRP/VZZzcCpj/waRqshSd8QoTbJpX8R5BIhmDloyM+p+71B5FQUY1QS1n
aLHiox9N3SKiOlzCmVeroaqUyeTXLhv3nJX5WB0IX5LuHgnivIBjabYn2U1XyUISwJ2WVnJ18UeJ
0Vn5aL53yM9phgyCkTOh+/JvfrVdmOGcMWG0NVPDIXEvJJLzQthkY4qbOz67QpA9oOiJ73NNlzUB
+b+QVXuizUZeb0amji3n4gNBwwvU8HKyFF4mNLMYsJCeFGeOPR39VaeN74/2IpaFY1puTzjO9Wts
hZnodhIvwH5kyVFolX4lj3YabQE//kzH64ZY/D8naLxEtMYJW0gMaRpvVOQboTpPifoAi1YbTg5d
0ycujqEmSlb0vmMpz3cv9gz7i3zqwHtwguSofRLog2r0AirMAHHHxJhmWa1quoVSx2rXR5NdcWiF
bL+1N/Uj3KRXl7ws7H/d9m0Rvt+7mRhepXc2gPBR1AjqNDH2rXGzoOpTCYv7bxhD9ZFv5EEoXsnt
y8jOp4Byag3wRUQfngtivapwHIW5cx8lbTbYyP6oHsUIUgifxo41As65tdlGgxlEVfCOCWZAFEsA
kwWjTn4VP819q++1+rGCtChpAmMFsILGN0GEa8pNxHw3k3BXQkxzVnJQ0afUUM3HDLAOwzcsDbcd
CJAcK4XhQm8EnYkdpe3ZwdjZ2R95cvk7Z+8ZHCL7cXaF4UZcTdR+GzVarUqVpIZioYMKYi04yMeP
WCgJLLk88Q8h7m4XT6hXfcDoh+EbFpG3yoxPhTXMi4REwr9f9QzLyAkBTGv20TqB89qylXHW55S+
2u7XEpP+jxAxyLOoU8tmkq7lafjOV4NRGR5kCUSSC61BGOrPy0vgVmA5QU7vOlycriMxxGa9RDg3
8yl/kL6Bo+1an3Ej/QXIG1GxghgtI+aCjr1wiu8ulIaKQl3XWtieq+7DmBI67BRZk1Cc9jkKArxZ
418S9vk1EZa1lsIikQ/Z+vktKULQcd8j01547xqhIDfz5HFSH+y9TsFXfVrC81KcV6WkBrm4XCVP
mMPXoeQmv+K4V46oxuHeqUGhhFl0rUJf4w8Kr8pqO45jO1vdmtPd53K4KeNUEug7AjacBovfxEbG
ZVktYiPfNG8ITEt56VLTQlc9ReDgWXOz4gN5sDUnS9EY4F9cHBTtW04lrgKneogP5pJKJpPbZ7YP
tpejZHPItTBA48HlaQ9ay8gguEbAfzPzU9cdVe3xOb4AnqN2PgHN0BVeKeRdetcDVCI1v8pwI+pF
RPI/9s3u265Mqhez+6WJ77aJ+u1z0YAq2T/E2eOEBPUxYRw4jyMBXtu28dwcKCAh5kPfKoqfVTIn
4VLCsXhIajHIfLsAbz+l9UkVB7dWCth2kjz4Y2D1vItWtijhXdIiDXbl9zTsxjZab8+gDgAvR6GI
nhYmDIDzdogZ9zDVinKfpW0fbouQpCo5WCAUupUTxsV3+4EJAWlMXluU951VfsJ4Oni7wBO+AR7n
Nj2o0chl7Tw++z1lINMCd0aPBdwyRNzRXIkgGeAWLJK5uadSh42tMpUbFIQA8K5ngItDY9hP4wsI
ouGaKrJsr9ofNrCnqGR3j0i88wkAk7IC1+c9MKXVDPn/i7Lz+gPfw4ziFPs7In08k3vaYr4EQVau
fWonmnEWClj3PiHNDEJTnYkl4OW/0/GuX/Egn6/fce5m4u3hXY8JD6MiDBNXUwjYhD4CCu3xhDYD
132fY1CtpIvoz3m7fXdFXfsbsRe0IPk5nyoN9Ck2C6jpdgtiFqn/Z0TWUJfnbIL6oFBVhk/ukFRn
68aqYNij1GLgGjGMhrWA5T+ShnKfs0o1xr9kwECtucLRbU3Gpk4w+8D4rXoN78VaftQk3DYJ7YRb
PEGG0uc3ulU4RbfQQkoQ+e6Q6N73Gl09Lar+10/Ek9CNMF0jkE7e6EKaGDOvEFyfs9hsNpiFNsO2
HrvCDKQcVhj5G0PuMQfaAwKr0Wiod8VnyZCOrZKBFUhO5IvtShccZpx36GZdWlilHf5EGTOJ5/3E
ZHMbahpk7QOePWC6Url9xS0bnifFddw5qLraHHg2YY4Wli6h3Jg9EpYRdLjhJIeM0GTbdRddWLwx
k/yG1/Rmq2EoA8Nmu8HU5zPmLc7Rg0pED166Ve/wXTDZGWT5vCpekCZdX/5cif2OMrbYsbfIrZOl
+Y3+XnXLDZ+du6s2JevynR4veLqOFtllCImnzP9ApIcDbMs+UXH0l/zAsWBouL+32I02+LV3RR5w
3Z/KjaYWltn1uTYs61YxMCb+8z3isK9nrKjb0sXhw9RXqNMemWrdf3jU7B0y/HPtveaWVCv836Gf
g5zlaoZp2bYy97AVTICqAxUx6yOd2ZbDLG3OqLa96ohM6e/BqKEldnMQxb4PRKFloWW4tZMYO8Vk
AKaiH8Vuy06f7sLTVpnFECjDj8v5y/MjWOFXytISjqBIA8tA0hquBcw0EcE12rSRaPw3flqDNwR9
PyolTg0xDl8YN3jcdKHniv6HCU/BJLC7SD/YZ+4ZD43PzLlZD7bY2vUw2jOZB/c4APObm9FB57j2
ZuVRluP9eVB8aUYS99m7n3ETNUE5a+Ma9MC8Gu9vkgFraM5/BXl4ZIXuIZ3z+kjn9VFNCPs7Awmc
rQ0h6jNZ7rWJ/wfus0aEWlIGI2FVYdiwNARH6/tZW+RkBISHZmjX7HEwngtulHDiXDJNIHzwDDsk
IXxp1PNLOx43orB1hLao0WG9tMl+VXofQXYacZNzBbcGXYamp7W7XUfdmyXfzgzt5eahZqn8+m7f
IiU2ANUwr/+iG4L7/H8sIFE0ZV/s/8wdpsiuP+qezDitfy7MI90tQDM73sH3rIgjPDhddrmn/hPX
mDTAu6ucnERtH/vpr0cJnXigG7NfQT38s4Wti63Kc9k8v5rglQqUov2YtHPXKFqHJYzSLmWexn5l
xzQI771TGfx1Zw79TjGWx3Blb/IgHWB7uOCzPAfuHnNBP5gwj5CpVtr1zDs7FBsww0oRrvlMdPZk
4ErUFbPWv7HXiHvse2YNFelm5uz2/NHPRma2hGy3gOSjGxhctN1Qar54tedNg0UrV9borXLrrId4
2tTGPC0V2P/h8p7Cm5wzGjozHIKAFDO0n4qfFakidlHuXelLwJZJUre6rg9YQiYRd16Offyt6+n8
Gs4s9uSCdzOf0If9P1QtfLB+2tN3ftULwZKA4cZPuF9D9vxy4gvmzKK5OXUlWNGU8SMxWxnAWB5u
QBDybD4k9lldfA+Y5bbhmayfr/p+ETTJUgk5rVrDmyL8cBDMEGAjfvRaEC1nWLelVPrwBrQmXXK+
Lg2MI/CzmTtmqWjpOp2GAl+IMp56+RYPC1EQsRVM9m5FOk0v1Lag0XFsniDtF78bwZAJnOQXjv8y
QuiMJXHyq/civZBBun+rBeRQHPVaJAI/CjRvNA33akBYopyrizJrIt5u8leaeF1YEDq9jfcPrubr
YG8mf4n8CUdYS6W2X8Jo6WXfevoJRlbIAV7gklLL1/XTRAr0Z1HK+BGWPlQS1TqcHuTr9l6yiwXV
HGHug5NBie5wbI9rJxghoGlXD3A98cM+1Ysxi7buqK2NbhonHFI7pshw7suLTSNpAA9MeoknccYq
BIPHAeLD4JVG/PAAnVFP/m3RYb5bMxsn8+JRrDeJaBa9Mh/h/HRiz02OqZ65r8EqyZozPzJSFyhR
0QmOrhfxQJr/mSVNBJK36QXCz37nB0iRqI4oNu0Wgm4x5Sx8XoMbRm0DBo0r08yTLtZP7e+F24tX
nwEXPDZo8EOL9/HJpgpkpGpzZlT7lJ5IXPYW7oYhJpomR5NXTgz4JWyDuZ94gskOj4nNPaCwq22t
ddMjdUeJaYQxki8gxUojiCUFTJHfSmxbqE3Nay0W3jtCQK1cEJHGIjmTAssyzgW4CPFxDpFCA8de
Rq5cf0Vip3+er5+o4XF3wL6CZXrJiBdgoB277tQy72qST8/LbulT7oWdFUJF4o7eccLMEk9zqQzJ
/hS3zPKTP8UPWcgGugSDuHy/YAd7o9+bhxZnH0+uSjZdMGof0AAzCiUzZUNsVYljH2LgQs1q2Ayz
K96pbRLBxJevrtLE/bHQ7mcCLNjBgEBnSpo8rXmKbWOSMm0zbubiujAZmJZUo43Rjs+yXDdfTIyy
Pom9hNqLBX2FXrbnWniVcTXZwMtRCM7zGauzL8gjwmi0YJgzhBx9l+9JXp9zJ+pqQZC7DdWR7cev
ht3vk5ovBbRI7Li15RdGodWP7W3hhaJuHgQIQPI78N0mtD3j5rRN0q0LI1j5t9aM3cXIS157BFHZ
iWkiO1r90Kn9IAiUmD+RlUS6HBgGLwIjYlzuXVsXdTjy/PHcrbfPcB2kXkzDaBfD9JbCiHtfrfGc
gjrs4O+VW9aI+SI/a+oKFoN3meShNzIdPA5z/XHKhkRIIz4swrD71NH4eUNMREkLBNwH4TNFrzB5
lvwVz4uzcQukwRe8jUAJB3jS3eHpBwvGUbbwF/vvSi3bMQGKSVSL5ZCTGaizO0wWVEj67hUwM7Bg
uFa6v1YSQEhcYz7SjmVOXYn2sBHq8f3J0k3i/nETqI95AItdCJ3Wm9PJFrmHaVAr5VgG2u+xjBIb
n93ftmgl6lssQWvKZgzkVin7u1tkJxkKKsGfundCnYS0jJehZOApH3TgfCmJrQyHbTLeORewyCZr
UBxN9Zu4QHyN/tJwpNwhl5PH45RtbPHrAY3HVeet07arFQRQHYmk7/d6MqCCz+Kdvmx7hJZFvUA1
SoGyKSx+0IEjgywIqNkg1mGC5yMTIxFGfJkjiTckU/7/67VARcIap2gx7YaKu+0bO+SX9hQefMDV
YX4nnDdQD0pmlfm/JOhMCPdUlmeQYkRgFGFBZJH5Vue/C7QreUYv+MXmKeWOvAhRbfj6xuRDxHd2
EdtFQyKjnv7V2IqYtf/1uIyvBgRbU7ZQtrT8W9GItGjPHgE08hZ8yy61vpLfJEEyj5gpgWMf+247
23mFFYtWQlpgAMwBpi3qLHpopovFr4Vqgffg6NAQxyRgH39xqRsfiKMeL4ejeDQz9jgmSY/mTGoY
6PnUemjTM4WDOuUzFeAOYLzdxvS2k5g9xPp1qPdEq3XwhU6f9yleWcv9R4i9WVqjT8Xs4LFPUteO
i/BdkpcQJAcQrPBikJAZluzu8FyazpbeyHo0ORBmvQ/0rZDV+47NPq2wUzFvbI8t54ZlT84a2vg3
Uj+SgAKzJ2oEDd66vyOSeYth2nrBbDmhywyWBdkUa4PfG4Zfqt5lXoYYVkL/iWLjohysIUIEpuCr
w4kLTKL+NuUOH0tfq+w7ceyI49/qHDzgumdl8C0NXEMGqzLoTNsd/tB2WZGllkBH2ieMKJP6cJWT
bZ5wDGJ/7qA4vdoUX6n/0Z4+Fvk3pV6gmMGp/S3r+zLtQM1JML9PVM/ltKtRf4UEZG7vCG1Mym6m
6ugUEmlNi0Q1ggmES+i34YQM8iIM7mrRkFw533IDQuRZTWHFbW2hoPZz8Z4pC8iHf78eVqn+sB8F
VX671NMQ+gNcIG2sjgy7XHeB+49+F86/x26WAAJUKhORh9Ay59LjWUa4SlPk0x6NrzoAHcioKXWW
6C1yrMZYa/JnAxs7aP1NQXxs4xFQpmH0IfoH8IFOyJwKVD0gyWjCrZyiFa2Qr+CQgRJbf0NH7jmZ
PgA70xmHsFf/trS6NHPb+a6fGkj76915GQ7ME2lf5jMHcIEQJ6ruSTXO8N2G0yh61/m9sPRfYuHl
eXn5DkcgEZA+nGjXs6NV6PZ8AfjCFWH2xurn6+QwPcR6X2NxO9zpb8slO2BFSxgQgPRJkkJxsO9G
ZpVH1Iot5RVKGf80hgwTJTY6y5IVwSfGYiPDERENN/fwtmvx4pmNhpHlUwenBflTS5VExADSnJeM
kpsrHa3NpVU8T98CvX0N348vn+GUrDEz+nbDKT6rg0J2B4JXhkhL5jKiKrIVQfVCsSzRZ6Se6HDm
IEl2EJmIRvk0z8rSLDvVok6I8qjWXijMRYEhNO497I+diXYkgMzU1ssglc/biPprjPSV2Gv/1Rp2
1sh2L+EgyFXMm+DsPh7lZqbuekxiE+j+JytHChmJnmVNGV6F0UPS4jotn7qSKN5YzIMT19+uKjm0
X9bIqm5HjwWhhVvCD57Q9w8Wt1ZTm+lLy/v3i96ULz8ggGGZ2gUT6GaWg4B2HWMREpY9C+v1AWLL
a6Z+hj1eDaAk2m4+Im51BdcbCt9WXsJqOfDhJ/FuR/DPfYIQ5df3ICl1dl+45zNKc8E3nU67zVS2
mdVid4TW3rJhOfZwRDkgkNFPUGXMX0Ett0aWDxmdFCQx+VqHAdmN/aRQRu8L6eKC6ZA/CdBLqMiq
WLof3dDqD01TbGuvpDgC5bHb4cPtpIurRLfyhdCslgwfGIfMMAiSFV3gu58a0MC1pKUoc6a4DXOa
/JJgjOoa67vH2hAOBlxNVF5ZiCct9BIH57JI3LIUcq7YP9lvOVo6Kco14egcRvg0vcjC18ywUXnI
4fUo0+kvDhCi1tV9MVPSChu/wIFZSA1JzKnkIwVqe8X3oOpfh5Nf1/7FGF5fph6R8MqEbRqaZAFK
TVHMneqvN+zjIKyjtButRk4ynonlWWDv1vM6MZpTUKAHng+h+y3Cdj5jLd8zoatSLd3gtzTDB864
/JDGpY/C+wr91ulX1mJRRVPW2UgVWAoRsgB6gUqeUC1BBc8cuLbml3/Xe6NIL2zT/hqqixMC0Pvz
XrNj7p4np9BhEJv0czZ+bjAfZZZ8mzy5R/FYDYCnZKoJQ/saNEDwRdJm1abQQ1HrjNNzACIsxwq1
6lgf66jhcHDiks1vWeFdSj5jg1vLm+MfmvrajShjvBjmrsZPx9Yuei0SHpFGpDS3nYuMMajq2Nyd
GKuWuAIvdMPaHlvqguGNj4OhrfRB7BJpSetFt2M0Om79iO1/fbXMHN3uVad2OzLdNS76GCrV+54g
mawRIIlr46PItBGgKZwtz+5oN/buZ+JlTEhc5jty5skYRJQUClSUHsHFjckIUn7flgQqXYccpch8
EtNS0inDIAkiiGYKQQ9CHBdAc7H1XjP+PuzQcy1pTO9nzDRy9B3DFqtsJ1JjEu62f3jmJobfiVOR
nLaZsubz3AGkf+vYQrkp7MDgxWxOHpZkejrLbvh3VZ+GFmejke63UDBtnUQDIipIrNpH6c6V0WWB
1ohd7pziNy0A5dv2Nj05wM7UFl9P6Ad5lEPlrzqF5SwCAG3rpeTCBUgDSl/2TAgFy1vAb4JPfBWj
+qIGj05uLQwbqdqWhajmrNCoy2wT378JpmCKxK8CYU5rUHW7wYEVgOvD0KJphJ/wA95MzeuEMush
Wekkdfqu9L35dDn8qeORPgpZe955DYMsbFEQ+wcnit1uJiv2TMgjr6CrDPSs6fc3d+ktzhSY6eyZ
7wVL/L84xdE9c8XUVtApaCGjz1YuUhQxlA9oxCTgMrN6Fje81mFQvQfPil50LB4k5mhQM17wMd7m
l3CoZ3rxv/UEokTAvyx8IZZ2vbB4rU2zfiLy0VTkR2pXBI2pIinciINPwHetkSnYy+Jr5Ef6SRMo
lcL80yZti1y7KoS//8feQzP5vMuxeGOn/9WAYLXZsj2hXdSS/FWxVCczaDNYK31/hl8L92tkAB+s
H4kPFvs41iQQifCmmWv9OrrP1WP4IxQvPetr8hHF5iaBDRiDB1kH06F4yDxCWF2325+9asGzRhLZ
4Tjwy9UYwa9Tpr+d68IOq4AFEVItT+P348iGAZrYzl3vN8dd+CFR1QobxjoVuTc4GSQfz0Ag/P7Y
freFxiHK6EhyOZvIs5l62K1zq1yoRAfXq35+UPDtUfmwEyc7cOe5XzrxE/TaoSwqG1C++9kcVI4W
KTwb2EcbaC3dO+gNnp8/YtDmd5N/fv2WtnSjlMbB2MLd+P3HqnNQB9ASmCXwhv8tE0X0JorMnxho
lcWBLCIcb0Djvu47OiFFoAfjM2jXYNtUiqbN6fbrDnX9+IVIoN58Ox3EZg4Wbnf3WeDLCH3gudJr
P2egBnPIg8MtzALfyzTbYEV4/qKzRvo/bVoPnKoIhciDTyVcMSqHm0GJmMTpp+I1DkfGUpuPbf8L
RIx3gbquDXtF21kKfk4ZXt4bRIahJoU4UEsGbTyNw3Wfx/zVFiva3HQzQ05KAKVxjsk3QwOgzklD
cdutlbmp2SvmDBfyY2bWQq/aMIG0KenXqZZKzdJZ6+Z8t82mKy6MmQS43n4U0CjUIvfMdNGogSH2
XRwPZS/V4MuO/HReZxCXHlGoo3kvaEf80sWilnPm+d35lyZ6EJYhOKSOggEAjrRG5D4LepsrhRSz
VCCDR3So0193FUeOJCNBsdLRvp21oY7iHmKq/h+XUMMmrgFBwI/17VEtjGgOGNKkw8MTD3sRVXud
a92Y1seAIToTzokHlwFmiWclzIMhSvCCmGpRCtHRJ+uyf+VrxJWIlqGYZ26avgdVv4dIS9p31hLZ
+B2yfxZ7hp1jDG5pF75EhmARMT/cI0JoXYtCp1BuICbKSV04Oau5sEBHlpsYjc/odAriQLoaWIC9
0YkJEOve30YNr2uL0wa6WU43MBayKsCw2pQKzBetAzzWR1/M1rnXEetynT8taQu2JSir7/sRHOqv
i0r2P8s3ioH+xLykeX0IT/VxKv59ZXuWhXDrkvzWHxeELFdbXSwk8kcjnuhM94tvHY7XHS5PKSIx
gB1fn0f/Ueuvb7zNp0+KlXqHB5NiHqdu+I/WGXPHR13BXf2I9Wce4c0oQ7LMuhahvWKmUptdaMmZ
aaXhIOsKduY6ZOgwGjAxvXolVTgsQQSVK8nqE4bLL8dxUXQZhmvoL9Xp0TSsICaRwnnGm5DIu22t
kRSLM39zFQdubQsz5FBKrkIbWercK6FMFnNEvabtJfiy9L8D9fAoSnkSUzEOx1NHna0zwF4rywEK
fImK+Uiia92nBeySrAxd34vDwv8Tqg9KLPjbPq/HkhoYVsuIodURZrQQVbtSrr7s3PhjibdFfNfx
NUQAvPBTw2SbjvDOsOHQXJos6kGB/jRnUpuyVZ87NmDc62b2QHTuFEKV4/GedgQlG6pbUgPqJwdn
e6fAXwKoAnJ65dDbA4g1YId/bZbTH4yAgzItqgexTR2ctELpfwkQ1dK6Ln4Pfj9dc9eB5MK8YhBp
YOIQ9DhwKk3q9BRDySc4XbezCuuyKUHB87euFftLuAGhgg0sY/e3/rcWGl9OWZl4U3B1IfcGjJAc
2h6bMsxvMzYHO4MxOs72x7Na7sNhFilItCFvVvYEQP9aNQvEvntqG09kd+qoOlQTISoTuJQkcLIP
mkmiXW+jg3JVIPf7iFgWkuQ/wNPkZr1jw4zPPpMNpIPeJS0Y+W6Tqv7xmqeAZeIo0zj4Wteopr7y
4xUrqAyJ2Ar8Lb3QnT8UoXqdZD6ro2NJyn1aH5cwyg87DxT8enhuykkYUqbMQqCU4olIaXizHKKJ
rdQC7AAVVajbgMm5kpSBiUv4D0e/bRwngMQLgD7FA+S/BmUAWKCUPjY7Iy62YA4PqjlQZmL3SQGV
2+kLXxNzDEAnfBWI0gzFneR4cIGL8lSqMOtyEbmOsB8dwYpH2v0RnUIbQyGHp+bVptkKp3ROls69
giYNnoaoZKg/EkxpDPaS7L6fWq/lxTO1r1Vzjqurt0vFFfGkUHXxmWYTsqQR3I1qhLXxHqw+cSdq
LTOWxuECIqSHNdiCUzTfG6PmhIsm1+cSlrnDBiOZ9A6e74bpZEi8T7PmQ0RgI6TmEFL4xTEpqv7A
OHq8WIuH3fIJV8BSgDNmfLDQ5ZrEEhOEpdh/nkPnuxqz9hAnp+kCqNNdGSgmvqFLb1kHADnha6Yb
bunDFcZjEeFXi2utvdK++gwBNfMr2mPCOqJbkQp86yDb6zQb28LN/fl5Hb2zS++DvsyBvlrJGJKj
qfKs7GsVWyG0+2QV68y71GRoo5tFp2+Gs6HuV4q4zWHHPsq2tVKngcaTpJTwfooYAHMiqrsOgQ6n
wSC8CsEtj8hnLdovm5o+mR1VxFoC8O41M4bDiYXNhONG4gfFgvmkUZchihFHRHDoF7fpP0VxwQrE
NT3DNlMYcqii5Edrmmrcol0oPSztkWLo5uouwtWp+mbZjjprGu5E+Rnx6zKbkmzhoA9CncxAyGDf
DACnQgVZbTqgU4J9NBjCJSMNpYFuOCly2zqG+5LuWXA0d5q0g4x+PjWbZJsdQcifI4M91SZVRd/L
z6eV/onyeVD4zrZm2FN2qHBbHHrEQj8F4cXdUPPGLvxDVFe9Xe7FA2sZVyeaE36U4Juh3YOM2WSX
kDhYifukEFfrLeJ6zqHh5hQ4KsSx2DBn0ub585SThNgF4XH9VX743TJssNnNQDLDoVKh4CrN0F0x
LXROz9eEboN/OUOTMODKTcjxbaX1emSUGfghdAND2EMZe3++2uBKkVujexBNhpUvOVK8ypVaMik7
Rk6JFkSEjCOjmb4BZGVrZAZJLls2vIT1dbgZb2tBAthtsDEIdIvlbKSP5S65EFowZJP1RUVoQB5r
aM084jRY76wjarWBSyit279SOmbLG6qasHikkpXTAMMxaUi25aT8G+XjQSjTFh8GaYvWoriTNrLv
bd7Zxf7SM+wICtxYfr8EtgyMWxITGz3daZgItyzV2Pvb7qTi33MKZnOkQghGO9Q1Alq6gfmcy9u2
DKuq6VRpkp6NMQjYSQOM2T0JRA2sBsFB0lgydWB1KA9BJeY1xwtQlfgIvDmwBQmZ4/IywL82dfxD
zGjtw7uX7kVmvXchdmB9uFkq8QsA450Fy9C1OVPQ94ncvfRRNj/hMMxph6Giaguq+1WMBv+io71Y
JP8riQzuKvNKPXse5OttMNSIgf7YG/g/bb+RcwESd8rUxY0J66hNQZTl3KIftXXkcsLqUGlxmcIx
ka09LEyyYQk0PrWFKC3rIvU+Y89nqYAzIMNcqqB53MEBXZX3aXJAIfg7XVYAKX78nzf1vJm60TnV
mOYKL8wEZuel9MHpUcof0hJebd9LT5L9oyYvaP2qxdW8kgwURAYpd+6cAbL5FhUTgXHEhgOuu+VL
I0HaQPmE10IHjqlrR+ZZd8VToIEdEh66MMZjPhJyRNHZ5K2wvehwnG8KqDRzX6Mc4Gnk7YT27fCW
eNQ8WrlRFXKv2Y8MooTt0Vob/SHOUb1DWfmxpuy0ZKxzyhrN4HTDQzMEaL8loRK79TkMrS0BxPb5
9KG4NHchuwa+Nnn58VS10oTcT147uVlL4+9WIdQCOWe1cEOmwqMfFCm0RO0TATDI2zrK9oK1kp83
hMe4TdxNloTsaPkUp2uwf6kBWiglptNOvRlBX+Cui4QQGLYlSkBQRpnZyKoEBnRLxr8XbjQ4Eedz
5nGYRmxDVYBvWD/oVuVqJn62q29tz4ACN3zvN0mHjfjMMLEEFs39cP/366wmQBPhIz7CPatzTbwz
n/+op8pKiAV6qNERXW4iOiLyWHPhRahmM0StqbYOVze2eLYw4nq6slvvobw9Z63Tf/ccKDC7tE5y
pGWT9G4o8aZqWc5/BSLs4D3XNbCtlTs8nYS02islc7Obj+W/mh8mbzuKITiu/YqLRN4SN4twbJWA
I06JBt3iKhyPOiA+zFnRUIjeko7NKH67HXCldWCzSajxstPkBN04R+5ag0IVBM/CKhSZFMxVD0RH
POq+hcdGwHE+mIOexD1DJee6a1K0UWKSTxnncn83qepPUbGy+ycYsOTfEdGANkdujuQwSE5DzRSm
LD88NjCxGEhJha1rIjFVqd4dP7CfhWJ9jCb5WHuJiYC2xHXVMYQJfaksMnKk0/KivuDPy6eyOGtK
h2aUidBkcehSvsQevbG/DNekPESlQeaeO/gY7FwyLcwsiFST6PXfqKZfsq1Oa8iNPyt6/rhNefZT
9rQ1cQ0VIiVYhs6xh2G0tu9+/6NLvBGkgnqEGJr+QttxZtmZCJy0SxwFaivaMjSlrGFLPas9pXBk
7KQZtXvk2cGQRYinOH+JmKcodsW92mBa6nX0mcU53IpqxVLu4U82Pyt3NvNzzo9kg+hbh7srZElh
8J9VQMyy7Ck5aRf8H16IwDJm7VXd0WBnkK0rURKR2EJKQER3g1wEKrZK/vQOWi2AjK9n322x0cuK
GipF3Jed0PVZzg50Z/XEkCHx4ZDXTqTrzODFn9niWWr2X1kY5m81ybqmKniUucig+VeJWz51BHgR
ulOdzvTwyVa/6tEJmQkTw8/8NdJi6cUABhSvlYtVC9NPoUUW1u1JpvQg1O5RfEGNkGvzrBKcRl1j
ABJQBkNqLbO4iZbAkkjbK+tGH0owr912esfXLBTTY6rUoUqYHvJbCY2J4f95nC1DZ5GZbRZ+woX/
IROiPNnTkrOMayUOuQ4QVYLXdYeYMOsRKi0NMN/XP85Xf97jxxg3euWNFIzrcxaMCbdrqxaxz+95
r+3f/4/NGVqGsczDWZE7jHp5cj5yYZKEapLGClmxCD8roEiDiQa20Ytu3mNoa6mXG7Gu3dd5eLDv
UjE1vNxoFU9xeF7fMjQ4RhkT0L98lzHVHzBJIgoOi3ln79ReHTrNzSU9YfTJ4kpFq9MMRk2fYYHU
CJnxEMv99TQy1J8bZ14Nhi4lrWBI8inN9e7LtNpMGkLR4aHt0QvdD9cLRGIQ5CCEO65erOYBKdvI
r25iO4GLws0OSz5H71Rytw77tLuMhGrgYSqzaCkKpH7d69xr4oVvrtXQl8BwJcVCflqRJxTU0HqO
ZrJdWonmY1X520S+YhlN4D7EEKB3S1uQP19XGiVsuLaNi4KqUpvOXIj1WCuWNx59cx6iHUPUJJyY
Ef9+WekcPSknVcUCGVROCtSC+VmYfraBxUeUnNpYyyPCDuareo9prLxKQdrFB+QfHurmVVH45KTr
of4IRcErdzkse2yp9aAYKU1CKZ+CpV8CWlInvoXLELodW9M4d1kF642BrLxgee2Et9xTKtQgXNQy
2uebJTdlA4mQyvecX+/5P0GYqU0XaQI5jGzyi/+Br2RZCNGwlWBQkast8kiP0Ilev03iseER2dUR
nW+zpPhl9lGy7H5eIN7PJFi/+6q1c5OhwcE7jECSh25UIj1ao6ieb0Feg+onZyjXmRrKflTHEsui
/ZoR0Wl1MLw/gup3SH8G4LIyhcUgVOvW4nNji3SyhVIfeTbaX82T8rx8KO7Kgk4pzXTTGMUZQBeP
qddZ4BZrsEk4D5RBgNfFuPlr+7ehpldiKye8YPHdfzlaKucjGVlxi4ekOCXNVpvfmqvKEq6ITz3d
b0FTfxYb/XLmDV2xLILUDkXSL+Z9IJ8tsNtQZFovFWcMexOJHUONGoJjzaXUH3H/eI1KPfYFMP7K
C7hlmMcWE6RiVLmqKDicbVCo8sDOy2jXRlZApyUvJhE4QY3paGy5psBvJ3O/Mh1ywBEkNhGn/IQy
U0zSc51GjWq8P9E+hzODDYZYW4K6Y5lT29Fttgv1nxe8w3QMJh6wg8i9+Uha4ki/K8ALrja+u+R3
cgDrs2qWzv8MvslUsNk4hV+GMpq8EcNbJSRP1BK4qh/MniOJxyYWINOcU3mWLiYNVy+FSsJ37Yix
AUCJQZ7ZEUwCHQW3LypOQuTSd82S+cECAIm1ru8MpJVORZWCy3ooLQJFURcyGp+6digTJrHvJM3Z
1VT3YjzdUGtUkFgmpMzwLIE5YpgESHXn4XQtl4/b0jBsaVcV/gEKcQEpexJ0QjK7k19KhCYrSz8L
5On/UZmFBHIQciEjrDsjl/8Nd1mSXSu4vBl38xC7RekgcDQ2t8lDbuIXJvC69eNita1v/oPxGCDo
Oh9ttrzPBFKf4fpVqddm4Ao8mu1mysv4uiZ3sxOMgWXC8/uGIUi274FNgdB3GKwGqdUaiB4roT/n
shCkC4sdQDSt3wF9SF98n347dIJ5n37gJ+7TyGmRSWVBPTFFWFnbun8CLZm5yHLQ6KoWl32MvaXi
TI/Cr0sgkXZ93FZjHKMFnEDTIQfopvM3XgyErZtzpTro9cmq4luFFPtfAQldmyAy/g5s5kaPOmaW
iSCbDn0C0PIpDeezRaM++dcPRCOakg0xSvVx12puKKgaRzR0s/ltYeoX/X1eopJF6r7SHrTagpMD
fWS9jLUTsUmEI7rBWAwYRSrPo9IyVHEdxnMRtBKlbhIxQXIqHdsOWjVbEiK0/hCS0FjsMCxUEXIS
utY56EgMGAD83yyq1ibQbaQw9dYRcggUlHiyzve/sEHsgj5jJC/HYHIPVkURERh+rMlQOl3V3YRs
DKPIxzt3xJAxwOjOXsq5gBdvGZdT6Z/vqgSHMpJEpZVIHUflajcE3+F1K00NWDFOxnVjqC2aMgNH
spJbCZqhUogCga/K1VseyrTdhBkd55Bh6KWhFg3mCzxlK0Yqci8/xILoZiHRsf7q5VUi9P43EoOm
jJKsWUg8ZpQsR2aDS3ArQPXywtfwsgA/1nYB5K9ZXTMf4BgzhLmR6e9VuOxYiH10AZdQBnNKege2
0YWzKerPDXIJSTGoPyZAm/N1x80kpyVMqkjJ+7z7Gf53a1S5ui4jDIZQrUv/M5+CStnOr2ZcH64C
lXR/62ZpkS62XFUmEBDoc2Idf0IXBNxCsOcbJQOgSIcHJqU/HnZvVOjksaFbybGVuXsAoY6vyHWz
8eN1b6aYMqObIOHkhnCKBCnboUOD4aHnjpAIUXMobTbR9tCQcrTA23gzb1EZ0bgwaDoFI5rDgCmC
Umko6CaSfHYsDs2zIrRs/4F/7DQY39WDp4HwjmbI2DHgMrPw2JhfpfWb9C2vs4S1u0tRXY10mGCo
D/5N0M2d3hXh6KNDaEo3SEsFeVp45oKEtIisXSWrZAbSHPcf6sCUxTBFaHzRlL5Jwsn13ZmkITa5
4TlIJNXdty5B+0tFh3cQ7fQV89XDxpyywoOaFMYu7QE4GBx6ZbDE1g4JnclF0Ee65BdfNYNNcgy3
M1iImscmcbpCB/W3XqJAqvLR4scFkWMzIWiycyPGgVl0U1iGIbflGA2XPhF9rV9OIufzU015jxox
415wGvrcE+pUCdtWpS5GbQwFhtGN22c9TBES3i2xUgmTDhOhiVc+uqmtMkaV8NA7m50ZoNy65Lz7
d1xs1Rqa5eZlFE8m7Sogh/ZIbdwXUJNekbk8l5C9oLSyymQf/GgpWCXEVWM5cX5pWieDqzX5sUmH
W/B7lgbb5ghkYYSyvneoubTHQZqY26R3fDeOLnTq2MFNue5uoxr89HVajg09sLuuNctthQ07lQnw
PC1fb/LaHienyYG8/Ruf+Kkz5Ou5kyoUk/DMDTkaYl3T/xVayPFre0644NC5o/sgmWcLTIyrqe89
Fla/xbxWUSClrwpwlTByQ/0msRKukTEFjnzvs57+eJ5pwReu2hxpBC/MFTusmX49qpr4r10zZwAW
kXjiXGyU9p1CivAucpr7Sd1q+bzqqgImM+Ycrh2MzSSz6C7ja1gcPSCagSTvVO8Za83ATc/cwvDG
hsciHygp597n0ka4zd0GT0ULfPIaTU5HH9Dmlq+/hRUt5IuddemnKIAxLgnXJLrSnlc2aZJG7AQb
6zsOWtUo++UQAyiU3nhXdmyBn4RV4Ln07WJTZN5TVFvipnYqAzxOkNjLTSheObvv4xK76GiZ50yM
0VJ84Aj/3yqBIjvv8SRapmr+MjkfAbFhHA40FIjCIuPYiOCKg50dKHHVXUgZVngpR4puGRClxcJ0
V+4DYRREbzuduFkapETjpX86aF2D2vzFoZfAOGAEpHrsS3Wax1kLDLHfzlf19em8B7F8N/yaj5Y2
b6v/Oge/l6dXvLdyWK/0302Z2q/Y3oMTFPzyYqEaNBwHVKB3elv0B4wi5netSde/aBBuLFrAl8TP
r2On9IR6e4IzUGYk4zKMb29qLknDfmTGNc+4D3/Vtqejp4alsW8bQwUufLPfGvW9KB8UgSLxVs3x
KLCvhdumli/XWOLiv3u0J3EcawuCSBb9T//891XeO7k7sQLPW281TNBTWUSimHUWLaQ6E2Xw7eNs
4f7HMPBe7D3vf5ShXPM5biioRmXC/jthfqnAh+0mPuK4aNXY0bJ5QejVX9PwgBaQJ1DFcnf+SDza
+Fb4Q6rHbjvfAAm2PAYsSuNZ6JCpJ837Qo11L4GJSo9H0ie24RRKm0vdVdGoek7n0vwA7Ps+zB9B
5mKNsM5C7WcJgK008Hmrq+uXyk7YQ1Ma6tII3vqjCBbqI3TYNl8d4CrF7WPtpNhdquwN2uQ0oOfJ
YReAQTNfYsrioEiMcuvEZaSUTXny6V0Z+wDjeg56R4DWDZ6VZZihiKOqOeG3YikTYirOqLL68Idc
cPvXWnitzsRswnQ6wqyUMQgIWJw7/yj/ebeagFJgrV4pV5fj9fUreXCuQu/yRg8pEdC5mqR3r+ZP
eRRQreDJ1VmI/fYsk1HRgm1MtMA9Akl3Bkd6D+Ln34nbVKNiNBfcdc0zZTt1l5Ji08ObaeHue4Nv
5truM1nFC+9NXM7Foq77/hgsbW+q51lZB+gJ4Y9wvu2vsH+kAnb4eZHsN+nG3qqmg0xbZz/qk9cz
hV3rA/nxhh83MvigZ704JCHHiXYFI5h06TGzYF8F+B0K3eU2CQjKpNSSqcFb0m6h7TZQeXqSE+R6
+9aZvnrZUZZmck1tryQAtMFU1yC4Bv6gioKLhI0HZHXLbgPx5cjKOIwjpV+j2dQDcnVd4HVvugAr
FuiZYwex2XquYAJgcePbcodTAmUISJOUoUCQjfHz3YDrafu/QXRvxd+8S+3KvnSHDDZx3rwyGwEO
I0vOSYFKWxRIJyYn4yNcK9vOPbW7cRGI5CH+Ndv4qdqXlQc4tBL7jrFkoSaDCgMvZN1b8kMat+Vv
4Gdt7xV9G+u/HL6Xu/9RxyO7NRNtFUV4mge7qBzh0pTKprLG0cAIy2x8KI/5c7OwtI61qDuFSUmB
O+/AGhhoui9qhqjeNoEAzM+yGase8yZ6lE7rIXsHpJUdmR1rYN5yK+k1Z1f900M6aYq6B1gog4cD
3Na+oftbH1AZr3amr9CtKDx/CQFaZs1ZbJvHMfPa9Dn59ftGY7h8Za9xJ5hXC4E1enASCo1fGhM5
yZwdbo/37UtY8bQd/MpfWOi0LrUpKkgwqRQ+UOapwBkP4Jewk8Uoipf0MGgoXnSc759LlIiLEhVB
T+DdPRgvajRxdRHWg9HE8835JAPklruwXel+nOSflDDIhBVJakD7OWfKo+kIqeX7DDWHVS14eBtd
QR47pm9T+Nsh+puOS8tpnnsNZtj7XAUufPhd+j2DR9X4khvhqUueN/yuc7h7iVlIlkTEZ2g7T4am
deMxokvAjZUE1FDO8UKRdbjpeiQs2tYa0VCHvki6EdpXj61qO3ryANiU7KNPFl11Q3PVJIRwyC3A
9StSTXbDFaPwK/yEYsjtikfhGfrMzTqMnZfCeJNb8qkNVhF6kePtMycmjSQi0I+SdJVJ15uSXOWd
ml9lYwi5HzSOmCuiQcRse6n0ybH3MX6GiIEcTysyaSAIhNwtw/rvaD/LGrFaQZ4bkEVtL4MxyU70
JxGGHSTjfHxAHDnarC0Tgkcfz15ztqjOzkuH2otbwWKtPCfP7x2U0T3qa0p13ZAQNNVbxQfLCZkO
INCd/lX0aHQrMouz2SRF+yp5up/KpHOxhii4z9hjHTx0hjNvP0TmjbkShkzlPnedh1Ae/HH83H/4
sajQpEj7DBtfdeqECyMMeV/ghkU3p+SF/8GH5ozVZgRhNr2JGiarD+C4nr/iGDABQhM3jLlX1sxI
ydP/Dm4CZIELSu6Or0Fry1D/LJ52dieliGQwhAIL+/XuGzfLSACqoXinHyV1rk9FYIrVAQwScnw/
1tg+SqTLInDSj3tfKacmSIPmcc0sLh4NOyUm4V/lgMGHygAGfmjh0v3YgVoK6Ev7QhG60mEpFUtz
AkJZhcWLrIvUnGpOfsw7OyJcDBUMf46b1D9yttb0ZjgmYKhn41xpHK4COT4Q4UkR/4lGWWHqXOIl
+oU5jpZC5H5wke9F8DJH+AhkY9pi/2OFI2Uq1o0ARRJXxmaYFcqwaANjPW7FigtX+CqJQl5eWfCv
QJu7jecdu+1LSnma7bpMT9dr45VZ6XP335Hrw6Ks9O2J9DX7yuPsnH5ZUqYS0//nsZl8V30H+qJr
MiD+lxCmHR70r/6VwPKQ3Nf6GtEGR7HrWhmbzPLtVeYZMNHssPf7hb7s1g6HqRqiyV2h0ubFi1Z3
oivAMuHB7CTq1SBtZlIgCIWdO7fq3yMbF/P8BX46eMCRFuJUoxOruAv3tyZZoJly6X5QngOjMSKE
EuurWxmO9kWCHaS2wtVAQaU+/88mrOOlp1QnI9R9TD6+Is0fOsVp6Dw/DK3Mm5L1M8Kjyvdyk7Wo
bt8PctSDqkbK0inVix3sOGQKCNYdPZdvCzbR24l2xqzw82Z2Tlm1VLkTZS9iFPENoc4JFZYI/jAI
dOhYXIMQ3tIkErrh0CBTge2kWbvKqMXsQdnUuA8LR86WMcgjvZMn1Aktr9hGXRpa7ExJMrQ2Z7VB
alfY/SANbNIUyZUo+94r04bk21jbJEPzW71XZndsJNMHaz7hHJcIpLi+p4Hf6KQ8oC5seNKOXI4q
n4vxZpHrEHNOKnXB/Zo3qkI2sj7fvCuPIK8AQQ67380Npz0W8o/J5vR7rk2h2a10k5QZPpUT0Ccx
0LOW+/OSbVjMoE79S8Xb2/1L375RH4MnErcnjzVJ7T+rF3FAu0CmElZkA1Efsi2uPQzfY0Z1UHOm
RrEOGyRh/A8o9sMyrhgwtHQDsgBpEO0C7RDsHqvTZOM2S98xbTa6ydFcj6QwBRzPCHC9NWmL2BIZ
ScMqglhftXmIw8qhIc2/hwGMCcWZicZfkmvS1lpxKEcari18cj0gXbM4L/z/PGxSUyngzj9G+o1p
H1SoOyJfxx3R/uF8L+jOtNhvCgfdR6SeEF8ynVm98y1StQFundZu1BsvUkt98HU5qWsVqPKXuHjz
cyHiJQ5+WRFQxAffcJ+uciALx/Ejg7Sro+Ew4XE1Qd1TqVDjbpY8/77aQPY6O8ZBmDJN5Mw0X/zk
B5qzciJt24AkyrR9DRisFoNmzaZfx9Glz7sVKL3JuKQFA8hvIi9DASbXXgI46DErnP+7ya1mjWWx
V8PJuBFsh2EQaa0TLG38/LMg0jwQV8Tnv+bBJ0dhfpI/xddq0qjNrZp7aJosmaGbfR0gGXU2YJl9
/60Rvty3p4aCVN54h+bfZ/Za3lkftuB9unZMYKE1IHjKQNqBmogt9uNp6b0UapCWviue5FMM/oK5
JEs1jsi7EsPWTGSsB1RhTtf7woUDl7UCZ1Hg+o1z8xt87P+6NsWsTgaHLT47g1j8z5SSNDISdJDY
WYcg1G2P3uXoau+BK5RWblk2fcI/xp7RF8YteSodM0Yqs3du+Gk+dnt7sdJxUS6opUoPgWkMUcPi
uWETPpkM58nVuKMiMxJypSbEsLxvFQzrMJEacjbX/VVf2badPmOs2fW8eM0AJC7dkGFyWiZMcxje
orKE4rYV7PlF0BIZErMN4glKDDaPv18fXenw3lTrOS9B0ePfYIX2itL7HTGkT9Q6ncbjLwEzL0sG
GqyDSp8xW/Sf8DAVRw0PZiUJrBZmIkKLNUjew5J/7SHrTZpKmMMktQ8ChAI/BKaS6oCvo6wWNq5+
4Gs8VV27AcgZnNxdZqN++Pms7WVMQ8bThiq5PHTpiVLcRn4ZTqjmRdWoNYRQHFJqWnEfUHJg9HQ8
2O51/IcbufWtLKI4f2y5s1UiFoSvEcrJhBwF7+YdLBUVGxqrdQiZygB/o2xsZpoaYZ9LHXxI867a
jeDMVXP5EL4oMt9aCAvT/JILubY7NwWVGgy5qVm3rZfI5jp9dPNVSyAKzgO0ex/DhfZRa4eHFi1a
Kw8FgldpYMkVIt1V1iM8nzZg5QxV1e7+ZbMHt54OFgHcbrBfw2/I8XYUCFYmhnf3ZH3rHmns1D34
9K0pajrryShn6Hciki31MVEUXHaY6Yb64Y612bO6lOc4RHpTnnP+VmJV9iBdfAy0v7jqzACiSMs7
OYtMCONPkejri2poo7WcOMnnN6JE9M36DAHbPQEsAeOGxF9DTbNVN/62vPZO5dhZjNw4srDs6MhY
azcCZWd8R67YPh+oKO8ioW5cGfX4CG51iwZjnVrvksz09OJRykzL4xMtJwSjJt6gJVhWfXQ8g/ig
vopOP8+0ZdXLhQCpEC1YhTkBq4KkiVJS3jEu1NvhBti3R4xa5FvuC4ieet4emc18p1Y8Zo1Gst07
2+5ZldKdqhl86VbAtFhU68gMdkx2vscm5qBPvTTZiENTknlsOTfpz29WLEgPOG/MNWZaf7wTc9Yl
EH9y2XGm/L81Q/TgFNtvFnAhaVIW5q0lIgyKnxvRyvVcqEUVcZRjwJtSZ3bVR/WwbEaRIIhT3TKV
M9zuq4n72wwZVwV8vonkZo6RlpbywgVnW5qnIHp11LjRuJwEiCe8sGrRWcL3NLUqkgb8DhP2VzcG
JoCT0uLIFV4U/SPIRwbH8qTGh9PLg2B7BRS9EJkuuyW932n540iN6MlcWdNpey7Y8m1avBwRQ9RQ
jJ07iFvtTmJHutzxVZ/JXZvqbKrMgCNFroCJLqtHMAX9V0Sa0dwLxY0xZ0jNbDfwv32asm9QYAdU
xHr2B8rxJlTW3br47vYxsfDwPzSGMb1Rq4fkrmml+niVWQgMjElNxDlYIfJMoT1RjOCZ+lhBaZLZ
dRkNPQffH1GC6x/RkwwduqfHUVyDCPTFhWt/klnjITnrqixTEO3aAO03Otse1HCBZHN76XEALzXq
QKNC4DWLA7icXJW2f0r8yfT3cbyYYnqYxpnC9ftPUHQlDIv/onzq1PACIlU2Z1h0JRvvqDsIqTnz
+RFoeh8gJfpWgoK6CbTIB+VZiczvwzuam2GDTJVB3CDpRIck3lRm7jn4fOd0xsJu/dfuPr+63ZMn
MXzquuwktHIMavxo6OOP77pZqDS3AT788PzpHicELYxIA94q5Pz0wSV4hc9GmX0h84zWriPdhlAd
j7zldbtPm5zCWgLEH3A0+ZnTQJEC5W/Sn/Tx80BkG1XKdoZ55KSU1g5ZXwBEJBwGANvL3v3swTLb
6kRBTA36U7Qrhgq8cN9szElKk59Zvj2sSd7VPPRPYOf379YyOmAorGUj7AMHTxcPDlMjdbV1eT49
IQfXyt8ls5LCNAbwChhOU6PMDTYTklFLzla4FtgzKfx6InKd7DhEpLkMVstB14yWUt3mDaqBscRa
ixO61gL5gOZ6KNvVORyj2sDsF6r9RzY1DTbQgWb06jT7b0YqBxUzR9GAoDy5fviVo3Gbw7yeJjmv
x/jVl2jKeLRFSQKu6V+je0dq0FJCpORFiJR/jSygJcr0/0rhMZ9Bk+9z6IXmNRy2Jp3m7tyKZXX5
VorjPr8zX//HKrOrUrqi4eadCxd3RLV6x53RPx2j1lN/shNeWB5A1hASEZvSFT+qbdYBJS+4S2fj
ub16P+0j18XPOTteaMUwwpjx9IEGGsqifa/njH7fW232qFvbiz8Yk8vJEu0ZMB0Xk/y1uYbY4cJm
0ojCCdOVxMKK4UqJtiBHLyPXtFyuQvOanrXxLc7IKO+fok3ykLd+FhV+xWSEfVcriv9ph1ykOBJU
n+qDrLfH3mtfw0dnxEPV7TZh3FDyHxKOWspRgkOeZWGpKkeyy9MWp8r+s3t6Xsjgr5Eg0/j6Kxt9
eHhoZWM9aRbOnDSJOkAsaF+Ligbd9uu11tWmBlc6z6gnZwxxUSApyZOA3QSU0z1J3z+sS+XreobW
3X81dNByD3yEWhwl5xVV9FxNKts4KHNx4ZS4Ic5v9UzQcN03dyYNdVYqOIounpdd5jsBT3F+8ik5
tg1ZyMEnhOsIglLXr2Gjp/0vSFrgdYHZYmkDch2WIIwq8++4jkj266m0gTH8Nd217wZpLivh96y7
wBUEMDOkIk69tvqROh9nRfXmAnst1/qTxjF+d7sBgJpJ814iLMaa1pTkTt29casGWJBwJGWpa/bu
WAMsMYo/cOT/joABSXGOwN5f0Dxs2kOn+SYCkIM9NRjmudDL42h0wXx46TUqSGwKssdHndOOqTee
UOM+6Nz35/WqqZXkEvnG8us/6FJBmywanf1uFOoB5ighmbXkJn1NlnHZ0C3sZ6DosHy9HXzlwwJz
O/1EXS0BvBWl7w25fmwE3YlwiHbTpkgrXmvgP8DCO38pNEQVgySaFPDRWwAWZ1RdK7blKC0un50a
M/Hy6LgWeB18nZ2JeOl3f8COA87zcTjazTmX3nrbrr0rcVYPbjwtixL9xCbfrhVtrDA+F9s2kofP
LQpVwUEUe1B8A5yd9n3Q2y5QnW/Xmr0iR4BJwoRRkASL7K5O3xnkbyh0boLr3aZIkv2QUz2LiqrM
Y4dI1tym9cMIXcQLkYP0vBGPN3DZFppA5M0B0XZ4iAWXAlNSrlSxiqeuvaj1zXt7B0LW7FPCea5V
tTyApGTReOnUrPj2nk88qEHwFRpJSmmjwSto67CUFqy+l1SkVFfyF3CPJfe8msab2YiSI06SuaAl
E+dZDvxPhfCG7/FYGsXaE8NmrVOyp8WUajfIu30TVQfIOkkALF/f28u2qJQBzfrskHzKxMHgkuvz
Bb30BdaQITk6/Ye706E+P9KUszAYHA14dHu0bzCRq5G9qKoaM01yVRt9xTkmT0RCYUW/istxXUdg
0s+t+74GBkANjm2RQ5qdBvJ0B1IF9TfzjuVWqQ9PcKtt7x81cPRpiECGFYnbOeOXjSiiEPf7Ys2K
eqJW2QznEaJqpgt/7W5b8AJseqDwLBKTJCrhfUiovdkE2h3VyS1gfzqMSU+Vco3mlLb6M89Tg7IQ
8+FOKbts03y8LEksNXmbaEeyKYf3C8UmWeUsMw0CIxzZLXD/YewJiLxJ1WqNpC4IKYQk1vniLcuk
+791CVFFqJZ3TAk8nJd/If09CTShIlQNSrvvTzq9WViZ6JzKN1wP0wTEDKelY0LrYVHcXC6baNEw
BorADkM8/IjylbiJySbG5DkGcNcW4ddxxUxZl6nys5JHowGi+iE64C2ovuwKEqjjtSY09Dkx9UTb
MuoMYdQe2iAtG6TEEHBZZWbD4Kqst1J+Cyq0of5Cg9op59vwv2eTEqW1EEYrCrTxRkiCzUOH4J2y
2zfR/FwxVwHyJ+au60MHxdTjUl9KGWCKGOghRFeyhRG64BmyM/gkjbeSlkRQ2Z7ePyPO15brmOug
paoXZOT0//4iA1Id7u16iJjf6ejz2r21e8tWZToAUV3CSuNSSr2NribBeqsKCroYbaGbKT21QgGr
h0qO6DQAMWF6KZRfNTPxX6Bjjju6ZZMl4qqyCKOsw7ykesnYODqysb2rkfLEPa1zGBtKa/qhOwxX
McjPWi6JKRAQs1IYLK7k2y6PI57OIusSTiZ+9ZM8k/6czc/35eE3pV8FSpIa8t6Sef8F25q0SQcD
dIOPD3lLgjZM2Z8v5Ho+b2didIiW7P68d7d6mWpqJo9skVW68/ZjHF5cCaToj050R26mpyXm6nnH
12hvLB1Dw1JaOerCnFwiM8yP+D3EqmaWfq84gMx2KGc/sG5ZB4GiSUhn/xz0q12l818LNyoJWWgD
9YZ72e5yroX45pEQgGvU6P0pjHIOyWdfBEhGS925QleYZHULb0jYYaJC2KwUibYYPU094uXZmZjD
TPT353GniSJY1fWkAb7P3GfH5COwdc4YqCm/bZ1QQZNynvTUhubggJvK0jcdHiSVVMmdyFLjpoUM
pcDVGZJHpmZioVxn2YIA4vC8LNGIJTScFw2y7sXTk1/EkfQ9/TyueYsKTO9oMPV3ZZ19X6Wsgg9R
1nCzGleHqEYihPCe32BXNK76ItjqamL4/njZ8u3s38g4LKVnHaxA0ogypBuhvU7gr2AWP2FoSGxL
13iGuEZ1XYEkB790+Qp5LDu6mXl1m0b5C9ipIgiu+0rUXK+kcPQoRPLEfvSm6eZA4oGkW77kEmvV
plQJ8boy3HpoT0sFi/PE7Ru++CCqAhJaOpDy5oXLB8bdnsFFkckn52OFTgaWPXkbB4qOL/UqoJzq
sugKLV5MC28Hs4LkMUgmk5PhQt1V9QCtQuYkaPMx3zE5EYRTYdnMyiCuMalbS7jqIxmKUl2yWC3e
u00CrD2w0tZDreNvriwAhwO2JFt6noi4tIpXD+kF1gSJH3z5bYvRxrkXsRfs6BaN0rXTDfld5wgS
3cuIPicf6qnrNTjDzhyKhDpA7gMD4tKUn2BQ0SSvUUFMn51jKE5drsNI79LvJYPEhsEHe61I5txw
omK/DUJaGXgV4yMc9auSk3pL1DaLstBl2ts3OpJadJYO6fdUerT5GkkpWPu/J3Qa30/zENOicFyS
p7MGSYvWf1GzbiCTAeush2pTfFUdGvakGUSXhEBOkTjzPzjHvyuPnD18ResRQYYeuQ2VoKMlvpcD
7zc0+VUeMEl8s0gUA6i1Xd8lJsdxpgScBkq2MA6dISoxsrLUsikU5Rmw263sMBbnVL7SjBOK9/U4
mIzTML68m9JMTnSU780gEehHq9SL8I6vXliNd4eI4YJ7N6w/Y9HSCTGHezmZjGg/zz2tDrtoGlzg
pH0F1N79wOM1Vpsnie8yFiPTgmOoSxdXV1WgiEdaPs9UyJZ5d58aKMUqnpukbb9cvSP6DkAHzJeR
I9OEIGIXUARUeCLgwzkS++cKLafH+z9iX6UyLbJLA638lZeIAHDZzMrudP1O6pSkgDAusu2hDafw
oHWgSR4pOPe0EFf9aJoS40u6GrfPCU65PYSH/waRJBJE5F7AYBOobfcq0v7txPRzXezoM0+6XWeH
ZAIFoRv8DzwCh77c5TXcr9HTLWHO8WjTinwP1fmkLdYqBUupLdVRKoRakmXeso1s0tn4II+DkgG8
uHVxROpanMKCd4lY1rbKQSjIxDNQdoXP4wuwVy4aB0ZDCFBeGCl+w/IuHJhpW+D9zfieM8qOwHAJ
8ir5qBJ0yWlb6meW+xzXaCgsUHP3hZtdoF0McyzJepdrsw+/RtE1VNRBWUSxe/egR+P9UbHnYDC0
k8KfmYG6P8h79Ux/sKIbh3BE66VauUdiYTrDlgC6mwIITMNOyMJA64u6tEJJjptGqOBAMiwmKBVr
BhfNnJacnQ1IVwrfN/m4iII4p4miUcFywdMGbpO8Yja4hrOL8bVRkA7twuQ1wsUUTWXws+omKdZc
0YjTleEwGUp2Gl5B0wAMqepFxZLyJ+nizWdHkDRwF/XZMSFalLwJ7HKSlh/hYSKPpjQEyJB2ZBeC
HTFMIAJZtQdwkMl6DbGY2X7ecegnPG9tnhiTvkzy2GMbdfvZYCWLwM0/ccEZX85pjoJVfpWDdy4a
zfdKausNU7yhFW1BcGOEGXMASrL01HtCD+PeeTCjRvW7p05Xv+bJ7Bl9jU5knk0z7b4VE3o89qwK
ctCptzIkqRjkqjISbCcXc5ZvgdkUyWteVJDrdRIU7uXORMmzlNXkRJ/XzP4NTdRwlO7dgHi1ysTr
YYSum1arr2j+TSvJSsBBbkt7ELlMaY3pd5R5G1de4wxJawGDi1KFY2VPoi2ogdd7RguIR1hRIBWJ
g2JiRFuGcNjLQAtmwWMp1E8Qsw/qXYvDJAMz1QMqu/qTn1ET1OxWFhIcWwxwIin55TGKNoLEooTA
Li2vIvgzRIfEHo3lknRRvCp3ISd5CAejaCfQSB4MfuQ+9o+LcS7lQHhMVKDt73daJzrXfBta+kTA
dxVxt0lOK3MZHY7DWK60dWp0t4F1jk583/p0MSca5sLCII/Wh2OQdk3g8eNw6LsuMSaRBsrKs3UH
Qprz80JArxMZbB77NtsU3/kA6L9WPqz7m0VCmgK2W2fi1Y/nkxvt+bqhFwbKyw/GV2t/aoTphVTV
ykFsstQ9drZIRNL7sHphWna9lwwr3ys8NVDPceAXgvujl83nGGFq8tU+Ecw8WN+WbWoCCpCWiBZz
sPGTUFN+f1ipKZHP/Bzbus2vdDMgYyr2GLbA7FUvPHaOGRRS/Xj6Zv+Lm//Aj17Lv97ymvecf6ug
3ums3xbJRbvde5YW8pK50f/W7emHCMnKbSWPpenu77TQu+cf9375CkrpTMrJirXHKdASQISm7pP+
oEkbp3AHdzEadHS5p40G1vHxWztxT1pAO4zRLXqzLRxp1waEiK6WOvhE/165kE9cE1UpXonoUY5V
tdYF2lSCm0O1O0EPmd6Qt8spQpluLu9bgbsyItnn7GFjHBqo2a2esqKtWoPxgJdTxAQPUbaHU0MN
fpYKutvOuj21bHpuTGuPDhG8BI/R766HUyYl7gZhKD+JYTI0r3uyCEKsEe+uiOplfEEA2ST/j/UD
b0Uff7RX+GlWTxfeiSsmyP8gZ1BoUwR04Ewb4tg94KOtCDbmCZM/2VgRoz8OLhceyQaFNEcC7ATr
jYdlBuflNlZ95rPd58PXL5/hjgD2g78movv50XRgLxJIisnwcCflWhe8s3wRGSEI/vivVivyhA88
XRCmBeE9JKxdpIRjxX3TtEJwM/nIYUgWpBLHNP2VyLngAV1IdmR+Js7PGjssusuustWbBQHnNATC
yCMLbDIw2CNRlARo1JJVzeTNgJESNJgC34GkqfqVvRWiogT94bEDbx3z0wYjeh9REBF4KMoAn9EE
H7IVZLI1sebNdU2BoA8mSaBTgnLx53W3ltbsXLrsKvbB0dYkg5PppEe1QWxdR9s8jz29AegYEjVb
QNF9cYaIXDLYeYIFHChckX7KpQKcwLLu7cQOwQDVMEAtAVGAbV+52sznC5JRmAb/tZLYh4yxrENp
XrEZIAXlQT4cQrKQ+/FdqUf59YBEWYopHqwUrpDve38+FmBA+ZUtwbGoHHaqxfehukJGQfEJOs/k
ZCcdCfP94ryrtkWS7tFFfecd8KAkATYU8IJLFrqJmPh0rWcoguq8KvMYgDOSB8u3iTsfkykMXQkD
YaK5/gVundgkbRBz5w4Jn+gAicPrL9o9KAVZo0DYoV11/RM+lrl9kwaeHUTgB2FHozl7Mu/dKErK
pEI7nw4oDSQGeYV5mHUkiyEbYv2xzcXW6JI4+WCAFG/STdio7cgQrPUzsEj4OISdheKHGbB09C5g
Q8JriOv3Kvlrmf5zdSuv6dvhg27kRqP7mWevvvpPiN3y0S1AQdd9gWNQKINF7oLJOv/hXxXjDxsl
h2HgtbQn2VcKnIfzcjf1Ebw8DJAL2iabjJWreaGbxg1cgCk+nex3Kb0ke3V3K/L0bxEH+PCj5JNe
bnxkN9BFY3kHWPdZRhp0uaIFQRCmXQGKzRzkrlQI2AjbstMINi7U0SKVV/BKFnc0o/YVqEHyq9in
QytBwXV9KGkiQc5MnwK9CArrRvzZrNUrybJT1gvi18aOYk1uMRaZT4s5dsfav0SF4EQ7LT2ssGFG
fh3jBPp505i61bnSyk4gaD+H9hDfxxib7m2oWrZQ8/IvezB/t4nLG5TN4u8vvcq63eFjuyUWrBrf
yJ8EdhD1SWUgPD3vNdQ7cpjkZ902lY3HC98aJSWt1ok0LdhMdALbUI+7GRlPlcP9rWMpyDzO9W7n
EqOpVK9mE/buyWaowne65dwTzNHoav4e4BQlDfdHU3KdPgOQgdzXE0idc6PTk+RgkBFFwBQB2Wzw
C/5wn0lokOWdVGO01zOiWu7k6PshPicZBtX/GpIXKi0fD5AY1kZht7xn2/TNW3LxwezcFAjp195a
fJE3A3fW7KvX2igmdnqVoRd58lOwZ55ca+ZChT3HR6UZJhjSqxCmAOw0oro4Mat05AjgxwUy0qER
cOJmfeXmH/AWS6VZ60QgmZzUPpetSbK+0OQYaM9+U4TccHqTlA5u2Y6aJN+b6uBLDj10RQ5oMyui
cY8ltRvYP9tDTDWirBaxTSOTHquk1nvQETDg5R0hyMWr0/WVN/JaolAsEwo3COMlJUp1qHHfKLRK
OEpQOKzY28tGM0yiaaz6Tl1NxziVDIDBzGQXE3RIa42Ohzijl1SpHrzjkr6qON2CZL5H7CVudC1Q
GG33egEDxik+N4qX7MN4f0TXDIXcZJcb9tFq0I9kfu9FldmK/VY9sjzPNM0ELV1JGNF1hsGnTcYc
TUouOgTx2i/oxmu9VpnxCDQlUkCyic/7F0Tz2DvbO9StViDoC3Nv4QWrqaBeQVFh99obESA0Uu93
95sn1XoIxpwMZNhPoOe3WUkVgt6op6+Pd+twsqIdG/eG6To6CS56WLA60wnGuHCZsQfTd8XSJCbQ
JtmBgWHc4GKwoaQfgePNDejT3aGDpIzxN3+hG0mg1mM9Cwmdw5SZB2d55ZPrWIJhfYsvbMrvHBGP
QhxVgtMsiW1Ghddtn3AYeqpLNVsk56tx53FXwFHGkI0NG7w1kaCyCniCOXI7LLyIXuuhfkzIQ5ax
zF0BOMy6oEfANt3Kp8qETIQtXQRB5QqzRbG6B7jXxoVRs0dB2GbpL4H9SqJD3RmFkbNMr7Uzt2r0
hJDsUXbdtP4QHQEc1RQUngdB3QWePVFnMHtQiH9EqSo5V/Vkpf0D/7TJKY1hgGtECfNo/bWUQ9+N
Tg/0Z7JBaAP4O4g7ICmAI70UE8zEmzit8lrFCncJybZDFuifwH4nmDyMj0BUKLykyBwd3g1E+G/h
Ia6uLQyvdHeP7pdQ449YY80oSLVxWgsJ7GadVD9pqrUOkAGRwFkWIhHnqVnIjdBTppJkYjtUqMOG
SuJA7SBIyo0MDguTZbQa7yE+0JCecg6FXbImquLcyb3aY3+dlBoz0FKkIGBF9dA/mtanYNzWuBAD
BBvg0Qh/rKbsEV+BW/5QncQi43Dt+OsLM+m28UsSyBMB9vTgTRXD9HAGoza7kvpnb4F19+jnVIrN
cIuEuyN+raOXwvAosX8PtU+KIKrenkJXU0MQ4oVpV6svSraeCI/TCyX4/dCNbZVvCf6nxScTVrdl
Bglhx31/h58v+AJ3gtD/8I2sSOotIaQux7wmXY/rksg+nu1Q11DRllCXgKr+wus7QQd6g+/BYpnc
Gf4neY+LVHyE8zX0mF9uzA/sDoLqwck3ZQoGK7ALMMAPZLiOMOUeYTrlbuqdUglt4kgfslUw6229
/n9JY+SEniKX0+VMdncxRJGUGDRLXGpDvid3iEQoauwe966uc53Plpf4gVtrWTjcnV3q8YMUl4bp
1bli2r9sXJIeMTqM9Z8C9JY/tXVreKyqxInA3nz7g9nQJEt8MD/95OkMM1kQKjqj/4JZPm16Fniw
z8zDjNICxozZvYYa5u2ckKonmSxcMV2x1C2psvWhQlz61eYN+FMcYVcMAVCs5PxYVXPRU7wJXiNl
Lq5hq5ByMC+hZ/fwVn0/hn9PRiWPIF+5lakL3NQBgPq/50NO0y9DXvUqTKkEAnqyOIgMln7316Dp
CWkZwZrEhxYDU8C5TtWVPEhFl277BqojyLob28ZHCemeeSlLq9OoHdF4vSOvqxuVWDxk7wjIwL/D
wa7naFVK3vqzb/f6x1CXxLBJYDt3P/mPGhSZMP9Q2dpTXP6TqqALN11y4Ho0VAZar6gblQVzKEF3
wsX04QrbRZzhTqXUa9VMUYNH3gtor0C6YR1crlX4iyRbKN+NXLUxrJawvdg+okLQ4hL56dcs08Rg
0l+RsvcwNSwyI/1QX+WDEdK+pxvW92drubnpb31LqYcYwK4TFCNzDYR48PfxpKjIjUCO84L1YctR
L0/E8yim/x2KhmFL8uOUjc01JgBypSpH6Quhq3wLNbQWUjZ7YgIEU4qHysXAAmce/uMZ5qRX03fx
/LIV2lhpEOkkToY115Q/Rbb3wSZFeyR1aWSyDTWqLGALfBLHkUWrV4vjYAV07TG+Wc89vXY1TpcW
vh40GYJgoB7CY4GVn+2HwQNUoaeFBBIjyEO2oO7yQatpf0Ae+nbGZtSea5PXO9RO+6z75LiUcUQR
302eP7w94WuaphRKR5ByPTxo+tipBBDhrOtEETLNWon2cD65XhDH01uoJ3wcA1WguLb3CgIPH/C7
zNrIWLQklwurAMoL2Stv98sEtPKw3ZYVFBqdoetd37FsPsj0YjeTBR2pidjuH1Ky3aSuryZ7VH/9
mwUVOQ7mLVb9DSd+m4Rh4I5iqU5VXDmHvTUn6yK+PPGVUqAOYm65gCY0SWRTiwV66Fad0WUtPLN4
GlqnSic5lMHhB3/k1ZCvAF3t4r6kMzVbiOz50CjHfDqDEAQgGOlMhd/vR0YVX/dMJNQd3RgtWf+R
9rckfPi1LZfrW/8b1aHUWauiaDrxuUQUeqvQDR1Af3J/wAN6eBFXWjyMluYnoPaY7RrD8YJaI3/c
j4ZI+tTUvXdF9mCiq3tsVO5Svg8mzxt+wEsGKf9pYSbnhnciPa4lmW0k+qjXq8nf6UZ1dMx4+a5k
4/wJ54pmWIsDzKUSzQjbZOdtJ+/8UANVU72JHRH54z5lctYOH3NHSGo9PvQ4R20fuq1BjnyPOqgP
JG/BiCoOAhK650CyJFrqOx/znSSV9dUP/z5bJ91BjTup0Xz0k6g6/I03vqw1HROC64DTqJs1R74y
4CE+SLBe/SzZK6/Z2cL5oOWuD9Xhb/aaSBqHb/zcQ7jc6TqYQ3a/R8f0x3SbBsWxQvNrtD7sh8Km
Q9KXlUyNQwldFspCLODmVoQh86wKTY84MHohUqt5RpCQXDEayH5FIXUryaOrTMUIZM/kVLftnCyu
MDpweZh55w9XYAAFuqGh0WIjZwOIG4A60RZIt4emfCx/ijgemIGGX8g0MJTYX1oWWk4sbt7Oh2TN
fBBP1KQzZc8+0vWekLj2BaDMPDucvnPsNQY3xuN2nKc6h53P0kiNlJg4Lb9V7KES+a2fWwa1JSj8
aemXaJgWJldejRh1QMqkZyLg5OQ9H0WvQQgMSk/NaWeKMX+SLOfMXdrEX92ogzJrZQx5xpE5R3xZ
yrAf8xe17S2TuwsdL24jRl9Ykj2p4MOgvrix6dz235Z/tS22rIqFT0ZqCr6PvMQ9BBskTxHI1K33
N1O9AJhtSujxV8X44+UF7maFckcSBem4/MWBsH3aXTPSqIrmk0SA/HFoi9mYQLEiKEZopk0e/Fkw
07oe/kIf3JnImJBFydkUaZMDXZiORGeLjMKVTi0gSgRWKRXb4eOQH4bkiDjGuvvldussje+RjXKp
56cfyi2xuCbR4Z7Ye4pFwAZr7cokXNB+msOaepIIg9WHz2V4K8Z5IhOVqybirpRtgjgoHDy/9Pcd
6u9wzzlhQjBBwBgEhU3aJ317mkyUrtikTnjr5apYVYwGUONS/ATMoF6RffWMFyZIuQ9rMxAQSUb1
BNElxPZh3jE0tVGzF/9NDuwCoK3ZkCDkYqcBjuBbYhGXmwYdx0bVAJIHuBYPhvz5X343vxlLwmRH
ClJ0H9aMp1j2A2Yfi1ussMQ5ND65kr4GXAkBGgZU8YupJ3jvec6J2YnM1KkvhYeC17TzihXEkaSe
TaqEQ1yQO9UI3exDqUBwPJ9I8KHB+ZikQVBkzeY4re2tz/vLRhceq8XqvZudaWJMj7uNkuIQO56r
0iMuEJM6WXZsQhvF01+5oKhe81RVIfONmtowhI40YFihTsSzbGKivBb8hDUhFP4dmDBRuByWiwAp
kmoSYUQaRSKeBpy56lWs1AmhQVS9zluxkgh9rQEVHUtZ7C9i5NPjpJpq9wHm6W2QQQb4Z8wcxlzC
WL1oSrdBGJWc+yeX7udfmkIocOtXcA7zAiU3qQr8J8bnfkIW+Hi+yu/UEuOl/F75v+zuJ7mY/Pfr
h06SX6WPAySGQ6oDeFB99FPGDRKtEktoD7oncqBj+/iT0ZnuunTAMa+cqNAxnBivWhU9SR6/WE5s
ihH5qGVGMelMV86YRdFSeinb45d3XtrGzw9X/qdX7O0iZbkSMDNNbnXh4zximOCyMKn62VuUhzF9
GGjczpLXyK/QUjXIdH7ATSdvkmB1ON98bKSmL9xTTMxc498Yj9b1riS/52qLiLaoJ1Eea+yyiyYB
PxhT8C+N6Hh5sN9H/wukMqwLjYm5QcJHZV+RA6+zKiSEmKPlnSXTPDjT0LVDhgjmSPWLoIhFmW+T
aIZEjSI0OpHM3unxtZ1b8aQDY1pDvCBEHQu66OyfGKfpTL8ZDCS8UbWcVHH3FKkGxeIHa8X1NDQ5
znmK/AMhBn1/L5X18CNOmChpiFe7w963nNSeiacu0T+4pziaawrOTLyeZEDpsMi/ZSmiyp/sxSqd
FsSVfrKJLmPmPAvSPAi4ip/HHi4KIVtWXlQqlfg+BU3Rj0JPc/WH2HUPNTaAFEp1BbzFu5TPMHyk
4WEx5cY7bPXiMme80K30Y6WDCgH8Lw/zUxX2bvZdiTQqJcaCSiW26gkJdXavU1VavVWpFYmgyU87
NOt+byXnLGvqFLaBLIQVXIEhwFta//rH7gQzaQyNDeb3GLCBVbq5f8/oD9f8yv5zRpJHhMWJ2jB1
UX6LnDk31NAWZbKBeYxWh6ACFXoEqLSbCeB9JbseZ4pCXjw1Kd1s2GKgBqVtlI7flNoUqLrefTM1
e/oispyLxbWFPQAhF1OlYK37EqJbIfwHMZGNUZ+eqDQ8LMjNWZHpw+J8sER6hB6l18UTbVQTuFGV
nkAbeW0x9+TgYM9y/wYpA/JwK5105ktLZZA8s0y4Iba/9YlINZZnT+BfApROBHHqX6+u4rT5vOeB
EjaP+DvsDslyuQeUo6fgAMMvlnZLLWCHf35UKiShKxQMlSSnO0zNSVLT7IA1KqYa2S4//tR6+6Uj
BU6M37+w16NdS8DLvpG6WcqrDu0iA4yLof1eGhPFFwk1TGWcZeMLiGKcQZgTiAuqaeHDm+6fSe7g
1khI2c886X/106FV1cr93K+7Em5+fHWvT16xPq7SfkEJ7hmanAOV00JaWg6RZzykxGdhbW0XMgkJ
jR1UGfSqESlghfsIZeXTHkJg0RdZdeeOaNBWI1IBjyhI8luil2QmZgavsPA1yORbKp5WJgX7c7x6
++0QEyhrBas3uBDPovs3NYDEVlpdMdq1g/kk4VAs1/k7MhaTbIE/PThLHqBgIV09nlf+W56V8dGL
3NsPYPez/65H70dG1ttDbYt2uzyH83n7wuCVfuPZw9jxPZze3grLhOWCsjrrAjK+ApNZnQeEc/nn
kpbVM2ZffdRwcVD9Qbs9LQY6Dy1juCDIkl1b5DIJxIfTLvg/CmPGHHi4UoJ2RfFTcwF/mJM2cyx9
UJVA49BXQwK9pcs2YAl+V4EHf2o6Ls+Dz8u6xjwbNYhEHy+6KF2KBhP9WYuDHn8f5ESB43EYzEtd
eeXbIBvZf2UPUbimVG7F1a/rUoxhFBXRdHfJ1QByQAvkv4akK9N8dvwIMj8s6jO7uJBgqKGEgaPO
ydyd/2jMYeTQMc3jWW2Bj+iAd/UFKTv1AJd59UUkRKI5snppG0VxQvsaZYy8eyD6kC/2PRP7BorV
W6nd86Ii2QJ5w4fL8X9fvBC5B3ZcEah26Ayzz2eFrHLBVsmi0yNzokLGTWW1q9vbUVPBv/23gWKK
9WcwfRTw6LOUsdMZNgzZwS/d77g3YK3RbIOK9fKls9S7uqgdEzUp4aCRfZQM2MuzyNVfgnCi/UzY
sRCckuz5GklQQ52v0YeXGzh9gqL5dy+nb8F29Y5sgKhQ0PuNzYcf4gkv1HEwwEH8gq8zWahxgD54
fOppQL5F0IpTcZ/cUFI2tbOEPvpXQsIpAsuR+tnHpcXIgFznk6i2bvWB9GJN5q+kWTmIRSdQfzDe
ViJYLPYfxGXDb0pCPI47J3ZXrg6qQhyHqvDUA6HvLwxFooT5lhEPX1/0FB5jXo57Ea7kx8Fab922
DAmQjfxSNmU0tRBqOJASwdSyFwk9oroptkr8wUPX7ymIQlgeFmYL6cdTZ9gwiSsN53YSkKt3AHb3
7KtcLQKQACmBvj5JuUnWKF2uRLE9k0aU57g7KN18oU+gl4B8LAMHdHkm2wcaQnDCrQCpXmTVTrZh
XXNm3W6rSApNXx2dps7PEuoib58sYbVbMSYOMPWxXWN7/uTLnOo8p4ql+2XUHZhaOfU1ebDkKmrp
7rfoV4SWz+zld8Ej//UR7R3V/+dVjVXtR6oPEWzWWdLj8kJOsn+lH5ZgHjvxCkjkonhE3dBfDumE
9akCFFGkf6qVUuLVo9lSHdRaDu7ZlfWYuMHI5Df0/F9FGbb+p3Fo32wS9iASxXZGlkR4C0HjE7NA
IFRqu5/k54Gr4KHE/Kc8efoT9ljXuyjYiwnrhUtHCeSo6iGy2li5Kjd2qrrdIPFQMbulKdgeAMNG
KKMj9ogpvjVEHKWWwfnqCTxRgypI97mEwpWgmvAHzCS5yMRnh1JD7jf2E+ojbCYPIzXwspKNNdiR
MZihBqygNel/UefbXWXNbafLBEox8n4S6jQATrB9WdmF7cspjF+duI2zN1f7bt5Wc47LYBnOOwgu
2qveuuNX9Iw/0TP+D/b/FbnNWVrohzD1V3PTzLv2sCbo0GJWVl0i0fCMmrujcuH4jZWNUI7ndffB
FFX7qvx56gk28MPwQ7PEa46R8A7i6BDhrFFy3tx+TJtlxqK83OmTiT4vayORAmgGypjYFitsxdiy
SiKBzmAVVvX2+KdXmDR7Hfp93u4v33iht5ZmIyEgs01iYxLnn4NQT1ovK49+wcRrkbzgv/aiF4tN
DraKXHeLPLkLoWdgf60OTaRmUMCqxlIXuU3XTKsLPgx4DEKAzGMEoN+4mZZjm9xt9S3k79hsHRQA
YSgDlhEe8C5n3V2QMNvk00dBrRRGmb0kkkDarK7mfsi5pmyjGT8kftsOQaHkqJN/lOvmGy0o3nQZ
Ix1RIoA5PVP2VFaiLRWjBGgPH92ir8KZvr1FLZlZPcyu7QmjIOmWYfEcQ2ECnIBAQP6d7QSObTe+
D571uzIHIw5nsyhoj/sisZVmGdTVSTxqU2FuiIcM/PhFybRqWA7E10GxuBVhQbicOJr1RpZco+Xt
HzDmccH2CzuDvjT7Fn9wteNKRNFRzAx4/cZY4EubZDknoaEizlx82hJioKczUjjUpTzGUiA8vQrN
fDgfusrhBQ/lMR3KV9saFOuqUJd5ONsgEdnriyUqJDo9MDseRyY+qRTZ4B8zVXVc5JITmN5K4RUi
TIppKHI5vjPzUBqY0QtNH8KNgN9ihpcFB7k1so9Bm/Ln6brpppaId1QJEVc6tIToTIhWNpKHxUQN
2DFtfNxPaJMLnYV576LyNaDbt8R+vAfNjRaMzuHDFmiFQlZz9wIH++14VRHXKUCtxTrjuRoy8xXW
rB6thVFJPBcnf85xWl8Gu3W+jXjAftqNCIWzSHFc0qSpUocyc2pPReLJ7X+XJZz9aQqeajl5zimB
IJzdyBDFBogyuBV3Zrz9mPmp6z2ctD4CTZemWDzdiREYtgEX1d6VHemAvfxG+Kz6Z2GKBo8IK0Cj
2kXg6UVLYKede70XLX8zXxv7zxVaQyb4BNtlK/yGfO7TPelPmysT3BG1aDWXNw5eJaBk3V7dbNFE
6m9O2cxS0F9EJPNBH66d/8vtyOEmKxAYL6lT0qztfgJaV9tSoFtXLkk1zcKxljVFqL5g1Vyw7C1d
aJcYf3W2iwlslbnOBWRGyn2xiEh6KcMEcJKqkH945Qp1CEDYro5aTZoZwcjMc02Hlzcg8oo6YDms
weKkiSOQq4KAJzEGGyS0NQmSLed9MJ+KOQinAwtF82OYQbMO1Gco4TVwMGIGQu+oJ6sGi4laDeUQ
dBPT8bPuHU2qE+HDlVU/IlqMMfZc7eWOubxe53ZNoYYh0JYViAYshmt7XrMBthUEpJHqy8qUb0iX
sR5WRi9NV5V14476vopGR10CJVRr1FRI5Q8vXyiN8UMK8/Q/9IpauSn0kgifRfs5yxhkc4YEVdXM
PDD4j1OJY3J5vyJmjDCRoJTZ4wrG4t0X9ALJRMQw/datks1kADJwKHqv0Sk//XFPsLF1cfLgrF9v
nNQtwqthoNEx+b6ySSIsp1UCskZuUc0Nifu1KZuTkBo481cNrPDvtZGkOvohDAwWhPhio1qaM/Lf
DP8rmJ5nL6BdEsrLXM//Igh4RJB9JGRk6JbFwigjQ6oz58WKBj56bi9PO8zYxrcLxJPkefXClQVx
Sun/ZRe68cMwE7XhhyG2EYEWG/sjrRGNz954aT/lK3ocoXuqZFXYqvP515r7MjJ3HIKwDzunr4BE
CyfkYmFR4YFJidlCYT05TxxmwJ5SynP2J5CnpY1TWqER8vll3Nv/4SKBHKJNUWk6Zg1xJ7HjDsrP
g0PNY1pTQqFbk2Hjg+KMDe2HVAMH1T75BlrH9+PM5WQHa18Yr/I9/dRGDt8HIYhp6iXMuO7KTAJB
Pc85Uox5lwAmdWMwZQn/se/UPtuHJUjQcHTSCtJ3fnNWHK6dWBX90/iJB26H/s/x1hqMjhU/4Ycm
oUduuCR8k/IE4uLsi7ap6tpsnp1DtxM06RognazSk/OnS67hILniyANi7q6micf7NyGf+7Lvspgq
It0lIOBJrK4SY21frEAeyAYO3zgA0nqiiuwcIXBYeop1CWy7D/mel11+dhxg0KN2ivNkE5q6IHBi
SyAC9tvsltCy+he5iBABiJTXdPmeasw+9qoQEZXZK4UseRSQXAnPrbtikT//22FJ1wKx819FTvAx
jvgo52uuTwv876deTCXafTofdz3/HmUmk+NxmW3CJWcOth4Im9hC6F7MY7i3LH6LCbIiVecjhc8A
+zh0fzSJdtAx+5Xpz9/OSAUH/fmJ7m8QbqVjMzzQYJvlUFvltu/BZxGZ0xmYewxUpyO/pVr2uelq
+VxUtauwyF6ygUavd5cmpFcHewzygdFgU1sSg4RkNZSGGWP4KhMJl58d6MdJIve2cNU0rRk8Qv5b
oP8Uphyu4M0kia3rwvgqPO+RH1cO+MMhi64xS9i/6K8+W84xrRwGF4EEUpndYHeImuwrnVkgXsw3
xeX53uoSyehCKLMPF4iWa09MuXGZpqpL/x0EB211Uv5Dd8TOzysZoVoh6HNCQwSmtKUUAC+vQ/Ig
gEoRjGwQYwLOpnzZe45f3GXzUPfq6OmmYnxiq+hOO8tS+RblN8UZXbtP+HpzItVlh7QMK6GQyjq5
pjNBApIw1Nz+ENrSkZ+rHSvnjJH24ekSMmfqP3iqdDUWkCJZeCuF7hCXB6JDmyaZqsCy6LlVhujb
ADHR8yuY9C1KQwv2IpfU4WbS9IStwt9UQSFI0dAg+uBPJHcGSNbD3QTrxRuoz134CoNwZHW/osiy
4d9YV+lAEZqjDYONEyA8j8Z5LL4pCvZBrCATd++U8x7kso0Ff+a7zTYTDRmYtmihpStlrxPkCXMZ
fJGQsMvvW+EouFZ5ox7aRFP/a1KhWfHY9ZmW6Bjj9LPWzmcFzLgNmQ4rDN2pSPtqPzz8M1WBzIWn
NM6cjIR464fGTPqrv4cqIM7fxUibYgTOKHtMs+A2UTTy90Al9GQXehODdspiDk4yo+QBFr5d0+pp
ofwNX7M/m6uDVgqQqbXA4RGy4EgspY1rMNESNMVtU93DPGae5uWSqVfjLIp7QAiIPH9RnaHx7ogn
Bbig+nm8vTNX89StWthZ6rPRIYEyENNW2xKHDRVYHd+5FuPzqOrV8dDEID2UOoXoTqCSy21horeR
nuLkzpDybr1lgCRERT+dIfFof5SVnp1eikipk/baFdHl9UNILomaGlfHZXve38oPyAbhFKDTptno
5r9lORfvZA5PoC555zSlrvEF/seirVoBHIJ8PQVx0mKoKP0uomGOlec1OasBm8DPkHYBlDvQOQxd
jXtsZ6+kRbOmNYI5A34y9I6X/rQ3vs+FUMtPKzHBrUr6+qnibJ0Deg3scMIr32WO3AjYzYD9JWfE
wO4U3hETOz7fVRQXUxRakfAkDM//SnTdJbAeKPqfd4JmPfyidvDAT3BWfGr7mtMwje6s+SmJ+Nj2
tv2wLl4INoP45IfFYr+Rnri45uAE2xH3D6/HHo2UeZ3hkN5CFvwmWcSUu5ih4rRJNXGpk/fJWUQq
9lYVh6Z79m7Xx7r4IcKbK1xRgnLFo9/GvkymYnTr4EoytQY9DPdFFuBPXI+vAUShnHZ815owlTx8
MjDR8G/VGIkpGZGQTltv4qSw6pPKtAE5Z7RTr676CksryYWLiGyF61Qty1G3Am/fCyJTyb4EdwJj
QVC9SgR6D7A23vrBgRRKdpBbR4GTKKcuN+jDe3V7FjyS3EY76MiFAf0zoF9hMnTUmxoN/axPSCcm
JnP6PO9drhi/y2tMXkm9NuxgaE1c2jwxN30EGTRq09HX2L9/qXIKfLOTXYt6wthqfpVmOAgyrr1Z
PE99RCD3L/56OAYmsFKj8U0Ip+NcXUQGMRjLHuxEHGBObNV+7xqDU26g/5/HrHNJL9ahs9g5lRs/
4fzZaCzesFy1DqVC6w4jN4uCwIFmcV6OInqoGfivt2pPonU0A16dO6wrd8MQx1RTsJvlqqPMzNjL
ffbushTEGTbyzVChsEoazHq0LoSRj99ajuZPn0L6s/XwdMKCflwRzzO4cFUHmFJUKyiPMPwG3rea
p/0qFkdF2nrKygZ9GXkBarnwCvAXR3HM3B8/NHiKppgYD+X5XxltESCWH6dXOc3/tF81cAYrQwTi
MBFLz42CrkOJNwoF6n7nlt7q/muXcBizW7H/KuKYRvaNwawwRaMYtn84BA0kFlTLsxRXMmrzdCN3
RbkrRXwugg4O+KfvLTrhqP7P2ZxsKDuzlCgS+FKjDsq4Euuot7f7AAywerAC/njHnK64U2CMCL1j
eNFJxzPq1NVS+pWlLFOaVlNTDXYS/hFK8KZvfxeOAsOXSv0kMxaDxgNWQSMPY6f9n2gNYUQsKNu+
dEyE2/Lz2SzAYziiXRXb+V8Xl6ltljx6Ju3FONYN2LR/ksFg3OsULteCpR9ZQLpGpuG4sErBVbyh
39NORc9XB/uRyziE7aykWenIM3+dbX1G329bCv3dkMdwfb0i0QMBzVwJ5r/xeSFPiehLEqmyZQuF
5F7IZ1L70DkV66jpdaM0YePoWBemWpgPg3GUr84H7gFsFVduiY0zyZA76hrn1sx+btD5r8p6/W6d
MLQb7AcBO51J+cBH7IeJFAsecnRchNqlB8TWg3aPnHhq5/7em39+cichLVJFEgKiP30wscZ5IbnZ
CgAmXqve+RXlXYWP3/zwX1hYwtLmkBV0WYY1ETfYrRrQx4wZgkx4lhtuH6yRB1trHFHukRAc2/2a
9EYzLjiM73b/9TE9JxVbk/J7Qd+MJ1tsghi+fnKrBy1+47Pewk/aTjgD222QT2klaB7T2WzcPKNj
y6YwJV8h8mhZwUzWwZWRwSztytsFRvWFUjbiFQdSxGb8HRNC6Oh0qWBU19E6A5rudtz/JM/JmAaz
CjPcuw3meJEPs7sXg8rGfxOg2G4XkPo3mFv2YO4L9KzrGVsTJ5aY4N0W43TutdSmmFaHMjIk3/Sz
bDGyiVqtNXPbOV1fnXZAfJ8v2HUptbWZoKvySwzbYamGRbs72AuIFZKwqybl9KzSVH4zzMYawFeb
0blgQGtToCaGLxn9nxYDIkrDIMxzxYJtajatwEXFiWZjGjs/btEPv0gNWrBwbGtjYI5mDKk4erGf
rTuZFNuF5FkWySNvBIhxh+Vn0GyNDP/tCPpXl7Z3lq1wEyyNMvh9PQeQvvrDRYCdqrm03qX8yc46
wI1xZCw93aQL81biMxMClRXf+jUeTenVyoWIw1Qj52lp4f1Zb/pC2EM0dmu4a3WqQTcCz5MMJ0wm
bDlykBSbz6MzSMdo0k3BeEk8hrzXRXKVa/hYuVzBzl6bIMpE1Cmnt0iGTRIy4+ixLfpt/tr3wPiO
mIfF9Fd0/Qopqi/ngXHzPcyaO4PRctjeUZ8x9DNXmnNrxpp7MYL8QK9XRtHZSSwGU2Aka+K1K0WC
C6ZsiPV2vSXUhhSyQc6T4ul/m0qo14nkYleLFIsr7y0koOSVeGERSAKphfmuoarKLonwziaUWC8K
LX9HblqnPgycBI8GlxDGnF8wt/ZRjgDCXfTNRMUWasPulC71QZWONhLLaUe6m1b341OX21AX+Mxb
w8Y0LAwam7pLYsKy2fC/tG8oAsk6vuPh4yDOHLQXB2qWJZSozANew/6jKqUam8cx6ke1M6ck3Ofe
cv0XjqOG55/C36xeautNkXeOqQTTvrtH5/r3dIuHYwRmh+d/NDWe8P2p4iHqwEue9T53JV2Lxk7g
tIDX/czh15UoYQcZhdzqlZakMwXVBV5nKnMq7841tgAMlElNfUF1GQJ1MN9Q7iMrmz2Vt9TJQgCz
oE+MSujzRGAeW8sozasloky/WaWvsIlWYVspByFDc/79czs1u+mOnoFG97TV+iHWfLw2Ox6jsTee
gj2PUlIC+4p3c3ULHr9O5x4P9vFRVP6Z36Db6zGBVPh1affHMa3s8e/v7OxH35b9uAkgADp1yQn8
fS74HAcqLr2BEtMaCVGr6PQ/8TS+cYPzkMl44mmBH6OnfyBUa/t1MOJo2C1Fzk5q4s8TUAHuOgs4
GoAVXVT645SKmMEMubY4NC2kkvQTOU7XLjci5HYih5kTFlP4Dc8IetcXPrH0BhrCDMUkR9yvP+39
ggUdOycQeAlwqxVrWf88dMH1bxzEtw6HV/Bufms8Q68PUZ6s62GvVnzsjWT27xDEygFaPy5zP2V2
3HuJlr16Ubu0U9B+y9Iu9hcKsXMFzuX1MikSTu9XUO9m7APLgzkjVD59lKVJNZpjcLvUVQ3sUxX5
eDusscD6UG43Wp7Zfxpe8TdFINdVrdonD4rQzWz9AScp7u7wZu/FT+BcWis6boRDNCg77dNpKR3K
LAE2n/aK8XWQ6HLYbYQmSlibfYg6MRzPQmNNI7ra3lPEb7H8XsCkr0lg7Z1t1t5Rw2t7nsXBd29E
QVBBASVKSMhXZ3ZC+1ThvHlFlqBjtq9aiXeOS4UIRKCNPEU+kkP+p2oVSypE7maHzAg3bGY731Na
FpRiQ4WY9gTorRjkNjVmFSiiT5lKIg7f4Q6wUIEkLoU9Cd4LqyvQH7LPnXvrDZbSeY48yao18gkk
Nn6lLcxsRspojPfWhlVnrOWuk/c5Sk/ncfgDnoLchGI0YKfI1/0No3n58/wXQUvl6sTXhICjEPzv
R5yASVyjCwbPfDYTwa+8naUf823DGet/NEoXA5ocKWuW/LZhvixBL1vmnY4TFJD2kbC0vpJ+sUV2
i5dc/1BRMevvCo1Ivpk1TJT5CM6K7m1pbJeiELI/btkBMtnm7HCkXGA9sYm0UOdo1Ln7W2Wm98h7
kGbNzNQoVOl2PG4hKTC2O/LGPCM6r/+90QAiXflBPlCeWQvVcu79AvlkYhqnivSyOnot9B43kl2g
tb8yqCIBdMEc0Xo+6NWgzkArSBr804JLy26rvysx+TglTA84c2fFI0aJ12mPL0DYv85RPBjyYgpU
MjqOzVYTa32Y8kdrgJixopN1eE3WwpJOkErZ47Eh++39wyk13cGkD/fZ1bHI7TExy8jiDXoDGJFi
6I+annN6gFV8MEtg8KcQIzTu64EXk5iWJ208eXW5I6IdMx7uVjLJe8f+g36qCd5bR383EOLuLvSr
bPdLWsbH9GfHdI+pAvs168BJGLTRRjq/LvJ/2tWgJQTR5SNb0o2i4Hm2/CKMqCv3scYxuGrYCYPe
EkQ+MYILtTbInHC1K9DR/3T9gseAhxXLLxcKfs1V6Y/Hpn7NzQiAd4sF5eKOEMOnlvkK54jX4Emy
mUGyEOM5s9AXec554fhEoEaulrcIzYrsLgQTuDidAHtKdO14p5EhhvBtecRsBUdSuLT+sjDoGUq6
uCRVp+uYIPlKwaZbTpbYfa+u5xc+X3XZQT3SEV7AgqMRpmQkfWqPmiL3CN/XrkQCP+JnVpHcdYS5
SJHJ6xcEmI4knG068kHCS84Q8qV9PwVXkD+7dXB7SgXMZO82lCdwN2ahA2dZCphhwmCww4IVfV17
dpBtfbqzU7EaPyXtXXgYjQoASVE53dTLOr2j0fYAVOY9eWVzqzRIpgY8oqpoAKLu/BzFEW6agINf
nWCr3XBuqUSoB+L8Mst/dY/mNY37Bl/Vmk/TkeEP6n7ErI5DJpSpuRUAltZYf8NDUdc8uVHq1wTp
4TmunamLli3aiRete1ySvqZ0jVmcJuuG80y/ounvx/1hPBD1hnQWVyiVr3RG2Xob50rIU/715nZ2
iAwBpe5/3A3obp04jrc60TtBM2NGjrSlCzfSstOF+rla5AMSbjiCH9eR5s7c9TC5w0m41EFFyDwp
eA6acy2ZlG9T/6GKPffIREkX25cSDpAg+z0vZIBescniAy5Si1iI9BU1bYPKIgpkbzVsPF/BzDZ0
n7Ay7BHdw0urrr5ggIZtptB3tIeohg0ignNCEn1M2FpCnoLktyKKPQGSagDaWjZP0bHGPgdfQqIZ
VypXLAE4CTcHQiJ+cMyDq0EBM3FL2t8eRi9lUMXTJWsh9FEKDH5mlNy2juumjoTjvB1ha/inmwHC
/otf70ONdScE8OqSsYUSogpc3mWwca72Jm9CuO727ciRMtoJiif0jtGqjO036ooah954YsrmWuPA
YtEshGcwmWUkuB6XSY4fkepOzns1hDe9UZ+dzVsGdzSDHbUcNqJZgNHZMVFe4qQ2luxrhFmBBTgE
4rm6UWmGHgx9tNlKXzo6nEl8o5l9rXE00lqXQkbtzYK73+uC9UHyRZr6tn2X6onFeAWv6hZnX8XL
B84kIhWWPfCTCwC3GbWebt8BxZpC9kFJLzB8ktjyg2ccgV93yaerm7tEF+iVC+3hL9v5dvhrPAEe
4aHmf/cLIdF8abgGXRsPdBDpysNG1INjYQ21DrrwDkFd6TtfdMwQSwTLoli9P5ot+eZpvAMmyf4w
kCgLHhrc5Z6LgX4r/vgoFH7/SwL4cq7GXkrmyheeG46UN8v6pgyF3HzFUkMOSz9ZDMO2ggdyICtf
cNLQ0HCM1KHVpDWxpvLQT/bFiztT/GbQ/pF/6i3aba03rNJPVz//cvrYM0Fju8fEWmILYmbAkfWN
u0hdoUKNwQ9PHhbDjWYc7cE5sb4EAaXPKwydOlm4PvFMfp+/lg0cqsquas99OQ27aYZPd9iKxPCc
TAaVjHhFzSnPQedomSOo+5CGqjfAKvWOK1zYm2V6irNdjqTwOzhTELE5ekoQaUCixhkikd49y2tg
QAjJZaF19jILP6sF903+oe+BrDnEm0Ll7SgmO1skDtHk7Cb0qoYw2ue7UFiricSq5N1rTV61aPu2
9HO2aOZIHCl4rhKuejokobTobEwTJtolp5Dk2I30xU6fdlDOj+WYbOg+/RU2ypVR9URRglNmhXfx
htGvWNnQJV+lh3QyJO0jFY/Kno/wZi+/3t9zaxU4UsmwhFIXae8ecckkU95W4w8oMA9mUkGhcN1n
kvjcfy2TCAhHBjmuqF2mM6vl3Y6qXFKSlxs4ZMZaZyGG8Y3cZSKrvzYSx6yiYHnwKPdPBfoWu8m4
4Y42y+Y/q0exMPpKbrQ2IT4859hfmO75sMjpUjNjwOQx6UTb9/5KFsFencBA/TLiUuFl8DyqMBmP
UCKQ67iE8YeX2GWnex8X0WJkXy0OKoBiPhWLnoGfO6tkTCZ5OtW5tChcPJ40yyBlg1o+yr5NOvwi
d8zIEwwV639EPxw/72P0vpvyeC8n80oEhfG4nyjpHP+wIInKeRMRkbp+/ZVG61Li6wVvd3XUbrc+
ap+MpTeNFXF4GaNBo2I9gUUNR8cQOlb2Ki64ZxzLWQx8yxT4GBuOeAv0y8hL/ATfeJuftlxjmRyS
IRQx2Vzoe1FY4mxlDFCiZUMK++ZxmbDvSqwtxGr7jdPNJmaRum8d50cjwnSOQ6PJbxRaWPiDWFoh
GPTlCGBtgEq1BAFp7jOSlnufiFk1IjPZUiE6xC3bgz4w7w+dqxVMIrBi5ErQuAX8aYi9B8bh5dCq
9CPbJs+a/e8+uK/qTCxdfJyWj3WrdyvaTojWIBHX4rXA1HcgvbVLS4T+uf+Wc5n6XeqQTjBNDf6U
BbjCza4iNvu2RwPX1NGaH90zoOTuRSkkYZdCq0k+iiXTohcNx2gKlLqKnFnDXIm2+zqxlzdDdCVw
dfQSOr6aT4hsIQooxVb1uO/04B/REWvNbj3uHnubyYtIMaOtczZpRmHkOKtfGqNwbZbZo/gv+l6r
InBKYI8Nz4CV012bs8QaMCjD4lebguBAcpkW2y1PRK4nO3uXtJoKSP3kXnGNUbIk+Vd4if0sisYR
8YLSW3fpbut1HdWKvAOZYPTit0PU8x5pG0BbfBO335Xv5km/1J58XuPbymW8+s1qGLyNpPikecBG
bQT5WVExc+nsbBEc7eryg6L/2JTTOa6I06KTyCU02pqm2+HMTiLvYayOPlh3SOh+IlASoNd0MQq4
Kx9gsn6OElkIcFqDrcunhTJlxPRvZ3ZJ2W17bKdgcHMfBRmL5oXJEwbSwA1rsTnkLE7m/cfMfeE5
mBcQHTIqEpRzIc2Rz0aeY0kfdo/Xh4/nPD97h3G6PtklClLaSlRwBjMStKG86gWC82SvakGwsWp4
XOpO3agyPJ8L/5t24iNWUg1AEs23evLNGT9+6famOvJXo6O/pr/dZ46iYlwgr+V6BH5W/AEo50pm
x3Rq4vIsdYJwXVP0UZSWzU0CgipYN2bQPia4ODRmHItOhRrkshsrQo9vtajCFozATBe278XykfjG
yFEQVB6eZ82KikP9bMGrqVZ6xhhV4FN1QfBo2x+AspBFsKvkrce43vHuPMqfyFrgjkECKi0CMjHx
WBqnM8TojXASbTAONjLdGSYEYcesE8kA8tA0hm5h8VT45jB99BAKavNFCtU4r2E+qXmulJfcHbQS
wi1VrJHV2eYk/mNXf6nhSYCh8bqqMy8BkoT481TycmiZhSzz+HZz8eJfU3jXINMLIzpOeq5fgh1X
z44BVxd7ud6As3TGzJKtwkWoqQYtvN9bQmqXTJI6yIW8Psy6a5aFspa0oqXmF1B98D1Ww/1xLeL0
sYJYGNbDsT4UKzt7TWSbiXae+3KuxFg9G4J9WVfHRT96pe31Y8JR8PSV78tACYn6ogcOR1S361sC
JOCj749HdD17lxCtk9fs0k2+0vi05xpmr3cB94Hh/mrbYaerPkhdHliilLLuPax44C2zv66jPsIC
YuNpHAI8abyXrDoT3Hnpr+WaVKpUQqV88JEz6NO1lqD3ILhRmQ0rJ73U2DaYL/CzyrtYNlpSBBYH
ecDXxf5WLKExhwHE7kN7efKRRMCo1qGx0EuQEU5dHHafCSemjeWlRtOed8sNeO5C4v6CIYAP1QHI
7VGLwQma2Qh63XTOxPEzelu/uM6uIfiC6oxIiUF0ozAu+mcL4kpZw/XsiQcfAkvQwHo8HEioBZox
yhmsCLFBaofS9hc1+GJD3DLtFE+BrqyxI7sEMQ83beq6V/w5mnQgVtnQtXkDUthWc/394vkBPjG/
q2Ju3izd3XEty00cRsS5B8ATEePjnOCElH+t/+BjaDUnPd5+NE0qwhk1gIXwxi/CD1VgqvPXPslE
zO6ILmKll57aq8LiTyIgZ8pv0fPV96nU0jP83G83+X7E/VxPLp3Jsuqtq4OBsrSBk8mQA+8K678M
OeYZGl0Kv0wpXHGZOTCfVq9h6gG5l3kviyRN8aFzzafck2CwbjFA7bTe4tTtjT31G/5EObJD7y7x
P+A8eEGvbyMDNUTxWMegCfQ7HAfg38j6cMGFx+A0ztxDyvSjOmhMKkY5H1PPPWg7AplZzaITO1xV
Xe1vCtYZ41MvFkId+GOSXkdkZfEiCTGIsZXPK/umNk69PJy+7bksu4QgffwDPcIRMk+poAu6uMS+
7/sWB+nrlHmBzN7UkN4aGYhsHVzpYXLWr/k6/wtdnaDVvTWu+q0y6B7rAJx5vHirDZ7rB4iuQwnP
SMSb6EFiBLLZ8dlHgv9unou9bOgDREvkTL99fHN8iGG00g0nqETlJA+9o2EYU33Jsqzb47yxlDKc
DbI4kAgDO7PeY1RNtyXth/S87X+Q3Qxqb3a3Ukh1GHVKWknp6k9M8lDdB71hm2yFsFOZqzJL78FK
QqOGnerPv0EaMp3+ub54z0jS40wCk0n5BZq2o5omA1S8ZLT9ZiIGoglnwDDnkrGzS/yOvenzqKiU
V6fxaaaCxGeDUPKlfbi0EcI9sQEC6p7a7TE1kGrLgpAKo1qYEZgm76m/ujfxdo5gc2ayE2zv4nNO
m/sAE449ctC99PIAo0S2Ydg8+9tRYexfZMG65bCoWVvd5i2lQFTKnegGgaA4Kem7jj7huGcvksIV
8y0Qx+2dV26TUMEdOiDBIkhGRvwjmJPqcq/KZaXYyMlKL3sIM022pcjIG3YOJ0C1X0SODl6qUTS6
TiiUsQo0FvdMy+aY23fDdh20OI0JRpd9dU5MR+mKq96AMokzjD4iSyi+R1UjxWJDNvMA4YkmRZNN
5HiqP9E3grdlbdV7XhbhOqiuMlYmiBByTjCbqpQvuOCoAIRak4WZvIipRZudNdn4ER6IugSb+Dr9
oeLfULuGSUZGEX7f7/gd7jwMLsc1V7yK0IOZm/LMv6Ohbiq/GZtlgAmTSxjKJva54/OdUoLJ8SwQ
Z57XeEL860/24I7nQPqZt54DQY3sX+4PCqL2n+xhsnZqgIAB+5WWhsk9TGGTFoptBdFyJ2DNmeuT
QUB3M6ZKkMzHuDFeoU1cp7Y9YRg0VGpbHwcBC6aP9BLqtVFV+1BQfy72AgMm988cIPrsMv6zzPZt
FiwK9aukuwsby8GBQJSBYb4pFGdmQi2ZlWTcxHlVka3z5GlCj4aQocMqzFihVPPRnTqPnE4YJO1X
NrWLkpCBm6pTlMIaKIjYPjNZr4ihX1NGcdsJrmSzDuGOXAXVDFtF8jT6eas3FES1q//awcOPEVBm
VYrDrl0Zqi6MAyovENAzrB0a0hkvpFF/qfOti2vruPNJGp2+4DOvIUj/BQrdwZqebEnYfBX4Z07s
rj3vNP6blX9t1a9+oI2991oh2JrcvGpXNHM8e/DfAQW3CgodrzDAgPOETMLkXlC5lSPNohSX7aWG
ntKpPhuSApHWU0PlzpRFRLXFB/iZoE2+LjHzxCvvvz67iF62k+0Wx4cnQs2FoQrBvkgFJSkVVMQN
YnSNSkPTV+NA0bph1/8+7U0HxK1OMt6e4ds3HR1pYNZzhGqhXKsAki4+D+zoMq2uIlsnzeiIbO12
SoTLVcFr8GmXf8t8LuztOINFmQvEKHm9DrNveH0fEB9YCRxkGBhnIUV/VR5L5NVP2m5IvZALxM0h
eJFtuGIGa5YyPehTaipR7JWhp8jvFISfIBXXLBjXhJI0JhM0/KhnI6kA4q6LXd7Kt5oKZIWb2+mX
tGhZIlsHBbUdhbpwY4lLUSzjJGivcpNDff+fDWp4ESUJtA7Aow/74LgM+5rjF3WRc0jjrH2dGyTb
xv7RHKVlJZw9baBPMYtc+Fvw8ItgMgtt1YFZbYGv00W+8qo2pAt871EAV/XFaPfjL01cmXAzuU34
fvemrCnwSrxFbYRxAtZBT+alCN9N8r3TZrPkwAlM+GYzw1kxxgvnZ5R4g00ZT825N3zgBxXtJ9EC
rQ4m1pTwsmfkNfXd+oC74Zek8vFB8cPRs2/uWlyGZdkCqjrNR90jlRjgTjEXS3c8/ZVWVqSk1bBG
eGTMnnJOGTV0vGjx8ILv02nQtAZRSXvCUuqYY/ZlUng/rDTnI4ApIdF9qZFFfePwuTTRPLItNCWs
qfKY1lJfvxKxgqJKJ7ko8Z8BVSyy6nLzSLvYZTNHH9F4F/jsN2X7hY8KSMeoRpbEUkowJ0fbgDpM
/IqRsx96VobJSo7sT5lssxwdyfLT0pSiOFZ68920dcFZjfhb5sIvKw2z2RNuyFy1GBn6oBxHNa8U
zXTxVzcqsOU52kli5gE6xXAYExqNYNZYjVNxO4+Xh2L1bK4WoK9ISduyH649lToVH1kDgIuEjXSq
YR0DY1ktC68pQk/yfMNuQ5UObo11/kz3wp7/Mn3jlDE52OAcnAA143aW4cCe5qQzyUpynqqorKR4
WDAh5YWQuxe+hDPi4PZPOgC5f7vT7x5hsb0hSORgCgtmQ59FExOvT54GaTi/+wE5EG5Py0fuAm8J
x67Z47vKWF0uXG+AL6cjihfqrK3NZERsUP4eIo6U4GNGxzLVoPzHT2/xBGck6GX0mkfCan9WytpG
FaYFBJMgkYlVXLtDygmpqCALJhMnQ464l4XjKcs2tZ9K+sDw4P8mdCzjigr3Uy/HXCcP9EO7XP/M
C09IQsyFMPhjv8OjJ3xD8WaFI7YWR42vip3WqxKyfjd2/mPcFD2mRX6XundnxP4J3Du7fDJcFxhH
oA7RK77M6Iq3lGFZemRw/nEHbx72tn+EUYEocm/4EddHc9AHRc2x6Uy/dOQzhDNidRCfFMe1jn6d
m93y0UfL6UoMXFJB/IqU7RBOxT/PJdXilkSuYnt5rbu0LJR89pkfytn96KC+c+53zfNuI3k8n9G2
bmAkKj3y8LVFmrohi8q4KDK6bIP3IiAjdfGIaLR+wP72dlBOFwlwW/8bwypBrNi8nNSsYu3KMsRi
f+nn/DunfBLqKNXBzM5EeJolIOcx2CRrtKHtrGwE2luZDyWxP8BcMaRI+Ru2r1BDfgPO0cF3V8Jo
8mErcoNJeFRbiSceWohprge/0mB8+z2CBMXGcjaQIE4eKb1lY5/Lv0Gxu/yVq2cBk+eKwMkm7pJE
rbeAYT9E5ij5KdVzP63vD0Zn6cXVrVu3RIvezpFMkH6do5MkI76MApFZ60uBdOHACVEMVUbKiVQ+
rK45Orp+JBiM401hg8iK3rQCy/u8Be2tl1jWlzoKFJrOOtliKjztS3otit0AQcDsN7O7RT70lKgL
S9tUwkjc16bjTFlDg4nZxcR4HF0QV5iV5FGj73hxRsh6YHByBB9m6neojnVkANUCxhnYJWrjccaV
e2glYWJaFq5Zxq9x53mpfWGjdKD9V8hUMnPYweN0OeP6+6oxT0xnLyGflLrr88AVqTpetBAUhLmu
ZzELJDOTx4XHxrFh3qzjTZzACREbnG91muUSsRi1bWq6adHJiRGamXgi23xjBaOp2hM4PGMw1HBh
HLa5lDiTxiDPkT2C+xA04XQuNbT87v/Kc8yNR7md6p3dMHnRrndU/XPaf8LseixUgF5+dML1VfP3
6a4O8T5l2E/5T+zSMlIUlCCcGLknS3hDSNJ9ATVnQQ781B0VP8as9Q2pl9F6NQ4CNrmWLYplQCjA
AAfchNrtkBRDp0jgofGDrDena8WCRh7J7gvuBTfa4Ix/sK0OTuKOHHnMoCE+d59eQfdbtdhxRYbH
YLhwWMhrZXnAOi0KCvCMVYoXj+pQ1Aa5gy57LeZlIM3cf6fx2bSCthBLxJ0XQafyZlrk5aF4jfQB
oL/98CgcPngVsmn8ypY46bOZZr0mWK4VslskqzlqdWoak1w+E8Wifix4YgPH1okkVMNJUhg44bqz
q8x3Hpl25DS9cpHVn/5XXA3t31nnDCR8qAhnLbtr997jm3HldQhzdJW4dd2neLb3WTSR8VzOrpgp
ESdGK+zYVqHB48pbIgEwDZW2kdEeA4PtO3PCV8Cup8JPBeiBEhyUsYL+BJU5mm+cQUXagH+/P8ZT
gmX9Ncedp6mjJgVstMFjn7oeBOOcKfUEAsFUywau+LIyRuUtMtt1mtLDXSzlzvY1ha9G8dzD5ACR
wzSWSsEoHTfrjkyasrMsDtog2ZhyIVy/EOeqMH8NVMIMRMHlT8RkCf4O00vzXta+i1IROHheyV7E
mC/qfICLCZEbQ5wDNeszTciwMH3h2WsHkHAzAs23lBHW/1yFY1wBySsTLKfr5AOs8b9QAYsGs39/
0AZ4hoM/pxnGNwuniiTazFDbMQo/avyObQcsfEJ3wYDDt0bfoCca+G0ORY45bDRV0yL9Ubiv0gS5
x3P0oh3bA/OzCzoI3kstVlIvkNOsJI0JKW/QeBrv4fcJ5BPO62/FAlMjKJhFp/+TQtmvPRIA0h8c
QozlBOpGbEaaY871Zqaf0phU/zYbn4MxnNVhmnaDqD5RTq16JwVlJm9IzZPCv6dQ3iqlpvqmkZy6
8GagwQ+FZkUYQEOUVV9oE4xyKnD7vc1uMftOQB+dGRxcjhC/rTnY2QEmIVLAU3FS37G8d/01W1MF
Gdux7aRSDJUJZsJLKBsclM/kxls0SVeEE5R4BI3swkKT1/scfQ4A57vV8mrHsIeC7eOZZLRDwSao
s/0VHQR6EueLzfWed+02B+VzoyXMI50AZkGiPJOrMKm4RCm0KszUiRcRoXzAGE68TVe0pCnGWHN1
GW3VhI6L2vehJ5CS92Z1ulA9z5+87/SsYVow6NVNPe0Y2XO9lq91hKPpmLvBlQv87WhU+QsstMzD
FeStDOgbI91R1NPzPXxRrq0aNgodY85G/qPKaPZNCU7F3UpxnedAAoiE4N/ch+Kv9PQyO/EBiUD3
O9ZMgSPVnG4/jsVv/9RbFf8GW405JVLASGjPnu01LSzUc0oedu8T43zJmzby6PmerVGpVuzS3xK8
iveieTxG+lUH8e2bDj5f3Ly/+P10sWLA7NfjpS+NhrMmOjYlqP+JpYW/aIIGgHMCi8JJXwHR0Yv0
inIT4yF8I1mTfEhjibRVizmixIjyCn0OYsFYaoyb6ds4oHrgRIeAMFcZCb3lRvisGsTSrofv3uLX
80lHW0AfRcmRImjpWM1K9oACGcu7clO7x/QsrB13+2w37/LHK49NHruvUY5Mc65/3EvsP+63vduS
k3tBBly8OiaO6KFIDhgSrrdzOEeaB9IOlkzSdJqOyLksrARsnuQOKSzO0VMbkfgEe8On3QkPJDSY
JghSDDuPnksSdGbY8peseqOR/eVejdX1ReVGHA0cjUWTSIMYf/SghpR8LEywWBBJxtiQg7ukTGfh
lROJbDpm7Y0xcmZrEah/rzaop/Wrv9qsOjtxn1r2ytgRtyGUt79E4+nmo0hpIJsbrtssJVJATPKj
NMwff76jxTEOKRXRv9LZzRK4hDex3nA+Y/1V1LKV0C3aPcvf5IezBdfg9CRvr7l5pMn+hN4rSNh+
OXk2y4f1axgxrZnzNtQmHAg4IcMaKNCX1RImClZFT+AfgRYSN3MkCNx/I8aaVm/bYK1kJz6/NmZ7
RnZwYga7DI5naa2stODajveGrWpxCeWOk6nL9eeGf/xGs3MyuGuQE6KISxpAklmmbFV8/sPsJO7G
bkNsRiiLSbjhdap+DGJqbqrr6CMRcz7/AgW4D/WXVau8WkEfymBwYn7gTHeaDQpoJqMS5BoQHbSn
3lLWmxB8PuBmecbuBrNUIx0Zs2q5YX9J7RSlu3J+fNCaSJ308isKGO1YZwNDregcyRTx6Vmd9ZF2
o8sN6prIa/qQMjdq1PLyWteW5jH0ykSlxRxq1u53ZCJ3987j5ZZ5M2MnZk4dlxG2GRT3DGfIqPS2
RnTIxDWV8mBsUxMd70+kFdbZK1a6C8I/rBvFXMDfGOvUuzyfIRz7FSJemdZG+b1PURJfrsg7ynY7
VYWh2ENqKRDMCsrzmwSuMC8dPaT8To+Biw+OMpv0ze5esO68sfw4PxkuxxRr0BcT4//KjNv8hFE6
Ejz/QwwBYDj2yWQF8lXquH/NhkH5vfQrHC9Xp29MbVGTeFONzXjPL4Voq5jQ/ysjfFpNjmIcCV6b
u+T6y+fuKj6fi9ocNJWkF4KK9Bmn63sRK140GOSUP3mb+R96eScn8DZow+HonyrTc//YcRFf70Ns
bBgiwr8UrvhDYasE+9PhlRxvfgsOWMckiqTMKzlbRsoUNB8BSlS/UAhe5b/BiCVbHenluTuhkEON
fzaqNst+kb3oXzB2EfvQEush3A6HRQDKTyBY4X/KRzeTJidMt9NtG9+3LHhIaxAWtKoJRQNjSHO7
I9gkqah5/OQrA1UfAnTGqGxA+EiA3nWBi6onqHba4uh6KVNgNuAHO0U19u+zN6AmUvhS4E6+EdxS
CgM3sRdByp9VjqSjTwppCNPLvbb8V7E+coBQex8cQOzoCpQOCVyeo4N20nhAkMd2TNDXqaD5+F3q
usSxpRJXGhDjAHugsndzqOwOW/iMonOS2z94lS1HHEr9QumqEsYK6rnDWvDkHbsCV+LQc9jLOWOB
Q2RdzXt9p2sq828J50ToGZFRn5/4yWJtn6gzxbHx6bLO0LhWeuN3+Fn6hL1oNB5mouZnpssYYJNh
H1rOwl2SmJo8NgNqyKaFY2GwHVFd1GwcQTsSRlYNUF+BChJOW0f19olJSbJqZDXa7tc9Fz8rFtYy
9jCBMGMA2yYPAKltBr4cf+Rz7DeEui80Q7OoIA7OG7x+9u4nTJDMm+JNlDP2BXzlSVs0LpaFDFWp
ZXGA53/FIdEEJH+T1nspJj7d5bnGwKyxqE/f8odPAuAc9EkFlklmiMOZlOt/j79E55gDdrtLQuC4
GSuaeR5qRiSTi+khb6UExOegGJZaY4O/0qwbTBU5stAHzZ3Zcxws282996BDfZ5Cbsl6FIaIsniP
k9FRB25iSXZwp1q+h3f5igBtlimvDc04jKnrDU0mht/d15cYZQmZHx4NB5yl8885daHvn4fy90Xm
eTlqB3QaI8+Vjw4SNwipUHvKYRm+Ta4gY5LUl5u8uVWdi2I/9SbUzB9DOEvJoH5CXuDfX3ypjbFa
HWl9smpaGrztI9SXLx/ABtN0H6M2QEYYprPSruiBUTeH/tcxii/XjJreh5+N8DeLSMISm8k+Bx4X
QJfIjQlrNytkn3zDEV1Za5w7POKuDadsRB+fsLLc5g3q9wySex5zUvmTrJiebD+34AsvpZ2WVWkm
wIKkCTMHpMMR4ey/rdf4WnNlOMrQSOPLTtFbN8BGHD/Irv7AfCP134yLiLg0CYzxssC1FebQhGOt
UEMod2DHoKC1w22X0ytl1vZHTnkFnP2BEqTT/OdIrUwz1phx+iQ1RKRdgoAmnG4omXeR+2Mbwwqh
kWJVouEUnXa0RYsqvRpHd39Om+uT2Rvl5Uu5ztq2CIpjKRPJg9KE02N5WoBk81ltPQNFYPYdKCJt
RPYm4AR9/JJc73ay3zO4KBJcUpSvYQIVBZSlY7c5y5e/k1DIlHxLlK1mVRJMbugsCvLvr7u7uia8
2x8jh+hbfl72h/yXFSS7kg7L9vDuhj/hz2mxL8NPI/LKGLMZ2etrc0v2V+FSBkORgM0eEWTeUv2P
RC6aYLDdcNnXDmlVlF0zc+J4vH0ODHPX2e1j/Tg67K3tgBN9VyWXhaUpJmNHNiv/bZDaD4EzdIwq
k7nCEUVlUx8JaoadH4EYSSnygyxc/GYudiRF/fNCFPuHrRO/IaGkD8nyTMbN7MLb3uI+pvYmAnvq
43/sS8QDw7KKCbVvPbI08kNb15hm3LSsH0Df4AJKbfirvUgLg6BpHSnCqCGqgJaou0tbehj0UzR+
MBkxggefZSKjXSr3toKPoiA8/eQWgDytSPy5WlXjo7LdQZT3QIWvNNtRUe4a4xpLsXjuGD/KBup4
r4xqu5UvYvLCfFej1Aw22hhgEAgIjguUHhiPUR1NIV2daREBIDm2QnxbHGMW5lO3gEtXPoyrWcUV
TWUDflmsL5hoWg4TL+yfyi9oA9xbrPXjeVs5lKPLlHMeF6lfEahRNk933TtWaiHQ+1Nk51Y0MkMY
HiSXn7PxnCRxf70mYMvvEWcfICSrCyC0AfseltMv5qv69h5GQ135UdYYBFkDivgGV5ENlZ9bI4Ly
J5F3SdtCZ5RSdoN4uMyi0HR5TsvAm9OgpVRZwn9ifNPhlhnQjkKZvLqysFpA5qEbfU/SRE4kpFyw
9TdQNAEDv4R9slNSPk7j0X+95WEHZeb9fb6iHD5PRiClpNHfAMAnBZOq6XAmAvvDEqpil+ccihoV
HlV4JMcuUilY4p0d4Ec+ZfsWAP0mzsMalmadg6wxQHahUR4PG2qaYsepPv8eLuc+9LUFM3UVj9DB
+fRmSfng1VNVIBGjc+CSNpeaBjf4NNMAS1KkWzAo7ruAM+cxk2AUcVVG/XGSccd3jaQj503HBosM
MUouUFgTw+98U7MqjkEq2ims8NfFA+TmG/bKVzapN8H7Umj/Mz9HwTWDVtCQ9YPwnl4aIxsy7SNq
ZpU1Z/kNtVs9YYUgPDf3S8mWzKnX9xVVGBGJNUsAm/Vr1g5wFIGS1M6ECXtM49yEgsZwY07ahD0Z
DjUnmkY5YPZXKaXVEm6vOWG683rtLnSH4T8wD7QHi8B+lv1P0eg8PWe3cpenSu8HdJuyHboGhf/z
PpBrBq6SlcKnQDw76Bnz03Kx1ANLBXaPPvKG7jLOrkp21dODstuqMJAbWVI/emA+JcTHZOWbjSqI
ONyQC2PMgzsN58BVfmvrfu+k+cdJEF8JKiG5gYOf4tyUAT0DokVbLJhwUDmQmbyIzlKRAp1igMKM
kDE4SKbPw+jCzLamEHxiwodgLGX/EY/7AJyK76/PZu1cUfd+fMDODwsKCgvhhx3YWhonmhh+Hzky
G+WO6g25sRskxjzfNZIHq5XJHICFgxqHI1C/gaD3oj+dAQLx5HPxnJYbcrlzhUc1iUfcql4AL/V+
VFEi3g9AUlvoU+MrOU29SydWDMG5dYtdxfbG58ELvx+cU6rPB1NyQNDW2yzn/7Mu+7jjahRCckWe
ejGrhJt8usIxrmPuE68/rqFKwzZss+DkRie3hVqa9b/JE/F0RqovBZd8VYl/H6s6HvSD6wUtb6wg
g7GebhIK7067VCDQdDcYk7AlrbSPRSY09CPE6Vd10ezA4/1MbMEYg87pm8OjmsBZbD+As+5maHye
DqDcn+OFXM0w6q09sExlRGUwSaKazPrTWXZQEvJBQ+i5ZPsmcpoAgyb1XId4oqqFiKTrMuiq1fas
jaN/CDbPmz2l62PgPWs1ydlCw5OBRaHrGfnFu/gN95sFd1d0/zt3yDcMOqXxF7sTt6EDjXymHr82
Hizqm7JgppVEKkJdqI+WXjp+n4vZp0Mn6KlGNjTm+wS45MsR61ZOQHSe1Gon7BAzJXAoujFXu3W4
iDu/uNKExwltZYlO74e8U/xx6UJm7WTRL8jsC07lG97GS0HagTN0SWaA0DP9OzDMZpIFkJepDJQ8
NHAC4thr1F3CY+lmPypxlqQ4IiPtC4XFwleow2Z1FLuUJn9mIW5iNJkVUqJFArS7591Lq+jcLD94
//1riCtJh8tqFYiaykDggQzyB4UYnpVURePBP/8BQ3g9YFi/ZAJTLV9d54ChaJW3/UD9n9xpEdQ6
jKx8zytD8sEZI3GgMqQoj7oHfOeIHtKccac5dAdXnorsnX+LrbK0oRH2+rNWjqIKu562qn/JwBeW
0aBphNhN43H8tysj/XegoqZU43FHbO1g9e9fwRDVUqzT1RR4BDTbDByu5mWT59o+kXB4W5JZ1wRN
9L7NM7VyqK3g9gI4A60Un4UJJ80jl16RJeVWCHLjPs3U9SvnqGnMn/8dBVl0nCyrIcCAhpbdRVUg
KqoD8qzIV2I+0mFkZ8jBJ7vID1fM1VGBeQrgueXXIEKeItpR38ysMZsJtI5lGJ428bTSH4Y4XENq
sHHzm8oSTVB0X0MFXRms7v85TdPglEI9mGu1QFffGOwREzoXNyIEpbweAlF0Bq0vRbz69uI+ljf5
cJht9vSKFjAkSiD+gWvXMslI1jXwqDpBJ10LQc2U5XjY5yFgKn1hmgVrUTHZd4ZtXVauaEPGgsUK
Vw+hCmBWleEej3SWXnFMVOf3IyUAkc7N0/sBUSm8FU7dRzlrcrr8CkyhF5GDQ7Nxm1zO+1ynHXBq
LZfI7OZY4YsSQrpzW9X1doHuLZ1dxCEhW3p+PoplYnEA9JwkWfH9YEtAErch4qGdWUao/GumoUhq
U4w9tmh8j1E6prQagdSHwjRCjBmB1dxNpdMAZCjdDydkqx5/gbaGdBZtaQ8dn3Z9hjsAnsuVjcVa
UdOTNM358mN8AAk2aqfqG/dQml0gilWNgUgivl6mK+9J/P1V2MbQgwYgCqXmLYiWMgN6oIJkurbK
lcTXChogPIQNyQ5+sbRyUvuUxbHFoDKgPC2+vNWeC/ynLoTqZZPwSEHgleO7KsKnDRNsk3BPXD2C
9DaLD/C8KphsHDYgbeo++hepNmsNCjay12zC1W8MrGt3xVSvbhuAgrsqj+TUzaddx1BP5N4ZJ9Qr
xdUP0C348g6CUb1fnYY+9eo4S4rfSmJg8vAc1fwrrbqbUohoS7WQdFTJ3qX5+WYkU3MiwOu65Vlb
A0woStdzChKZ5fgjHQ6SQ4cpPJT++MOv6Oa+mC4R+LCsX3Ohc7m4pQtRDsTAApP5toRr5xtsZy+7
Y1QViMixnEfi1cpLCQ6LR+Xs3/xesr2swtgLRqMIH0G7TUaE3jug9NBk9kfcplgTV2TGPCeHOr0K
lnHkRTAMeRJy+oKUjt9Qmk7KxctrIOkKY/C/V3/lHxc6tQpWTh0fKiKGdGmL8BhNJ0jsgdEJrZ+A
VI6Xn13CgbtWGUXjuzdk233YS4/uxUWkier1AjFk1E+/v7oHbJkye+NGnxgeTA4+JV57BsUdGeL1
CZKGwKx/4yT/mENxZHQ7D0d9Lbi5n1tjfMuQ/Kao8CgUvqwSUYmhKhckmyjzFZ0dmb7dM0b+jmS7
vjcG2zRuke4ehQrwRh4B8HrRs+7o0zFNWri0FlZvNna9bPQ/Yg/5TsD9FU7Pl1Z+II4+rGYG8EP8
ACsu++gJbcLbmaOcyFLMSvnlidhwfvIRs46fk2eBpouF/SXjt0mALMGtTZvthKUCcH3Ic0DjLCL2
zXl+Nb3rjTy9TEECEjLKoLE5K8XH8hs+plO7UaODaiwydEXP+wnLMlElUp2FZZE7VkpCaTZXlDBk
uYHW72tuFx1vyaD2kxbqWaRgCILeyeuxd5nWwEHz8xtXIfk8I3p0cV+pozf0VzdE0456tkgt2AAc
Q6VSjaHGwXpH+Z8sZUyWTuDpF2xoq78qT+bMD7M7r4aBqw+HdH1zd6vMAE0l4q17ksvWLDhvKHMo
C1p1XHX62746TQt0qyMH579BIzO9+PLxZN94GMCM87F+bgpApl6f2THBBisAhSZNhWHXkRahBpw6
QGL+LN+vh6KFM2UliDex0QxEIjXU8A9XBU+2liNwx/U4zz/VloZMeO4AzCiurKAxaRww9DyoCE6f
fDh40SiugQw1PieuvxFTU0LyMTEURhuNoihMEMpoZcJyP4L7f2pzsXgpYjKcd+I/EbKZ+eMenBDX
/dprVxB9vRHT0JeYe6Xjngz5232U2VZK0d3GHOgXxc0scankZtfd8Q/jvryV/hV+uODqnCKXOZEZ
BmQxf4XT6aOu/fr9v90ZsbpvyMHtFVSmLuspW53EykYPsn9wp9IDtfPuObxSnz6OPCKkcyl3+Job
rXKMw7utNZsdOEMezjpkH+dd6VIYr4UkPvTCy/QCAd4mAQ4fdYcbR4R0oALVYTMaaBjZJC8sNaYb
ug/VCfS8iWuIIPGemi6tuSGYnbzGsim0w7QWwtfn6kaA7vscXLSqASZw4nLILLYie8Qxg05w5UeT
d3vVLpXfRp7MMS07gRxjPQxKGN+BrkHKlWCYsQDdBRu/1uuH4mxOjANcdeDgiFF/7CEXoKr+Xbrk
8SbyK2t/LoCEz24rZ/0/VlnZnzHR9RkY/8qdZPt6sHUtb2RSTakG0cBWdpFMbVCoqmXYZHxJUY5N
/4akDgJAGU4oYyZxC9Et1hIwaej/hS47w8JrO55rad9DlHar+6VeJb3+/sSyXencwAuBMsC0k5O0
+DxEKwfEq3SQk5FAxjfiVjqog/flgxabCdjlR1bT4/QNHUQzMHQRc3G9WWRx3k3FJFtfMHcB3Kg2
AaI4Oymw0bDurRl7eg3CZbueIplnRw++S2UQGx8hWT8nIEkCJUAoSpUetRaa1YxasIor3113bjiC
eynkLzOqASjQxDNHaUSds0p17q9QXu6v2ncFVce2Z4u06qU5078d7F4fQmV6FJ6xJ00imI2wvaMZ
qtUaq0S5uUFwETMGaG2tkNIIBI6U/1kBYw/nid/+rvjRrTrv37tj4rP7b36sus9iG47dgKwcSpiS
1LAymkq4LqwVzEAbMk5DX/aF0dVPwDag816N/7+kKEo9z88MPW4U8qslp395Rv12/GUTKKnspj6V
VKvBg41AsUW+9CcNyvS74n85019803+r8gK4arLSXF01IdWXXMQ4ISzkDCyMItB6xOOnuIZrLlbg
j4VbYU72sOToB/BQeBHLSBlawEU7BNI4p6LNhzB0spsCmhbcOlp1Ddnkk1gFAdDuIXgFqQzTXd3k
T3ajKis7dFahlBOELgLuevY2gOv1Kfw5gDGucLStU0yWW20ABO0fLRPhAu/c/uiHro2yPwZXaRYu
506U6ocjfggUi+zzDTBzDTpcLammYGiW9KCSqEdS8EorHFytkfonOvwxx7yxKaNME44uSc/Lfm6D
/ktV4r3JCwrocJ1tYshB/M3XqK5gIlfaeArLw03gnBWB3k6smQQuQvIk/QjMxb+PwZu5xO+TJnS7
FAWA2FoA7Pf5UsdjGY1hgaYyHMERQLJoWb5DWDTiYWyuADRhFltl9vHwXkVMWje9BSejSSQxPHXH
5M0u4DMjYP7N91e57YNzFTjeqJlhlww83tUBWKmasO271Wk2pNRTQlnKiuCCfC1JsLaNAPwKbNH7
kjUMnOqzvG2YBgOMO5aw6Hm7YFmGD+tD7XNv2SwjaSUu9X8tk3reX6+VJT/GaI5UBx6L9j09ojS2
SbOHYI4MO/g10qiyYg7ZgUZd02ZmsOziwquu2H5VX3/wZv1AH62UEHrcjZbQO4slIh1MJgFkW8c+
93ompJPKRMy9wEsMbcK6Idy+0lIbx44eNQ4j+O+3eIzDq3n3EZVb6rx8vkOpKm/wgRi+a+nGSN8q
hWnb2VW+2srrY9DtwsQngGrZDRmoNcW8KTDeMV7VF4o/1WU3niSWfMq/Uz8NAVJWyw2V6Beq0VD7
W2ZwuL1e5biz1TS1lCCLZGlvP/Kx0+Rq6J8D1twCXD4TahX5WBdnFH0ZmZA39plSTpzwVF4kZIkm
t6eLUhcBI+j6OyoCMj4MgQkXxK3krWW+YF9fPjZMm6SHLKxwYZjB+uFaFDRLyNoV6x0YENWv97e1
ocNXuLOZBbMzm7IkSdMwexWIVHOGsKo0/OtKTKamyJbOxNhPbCk812/y8eL/+kwiDQQdcY8rLCfK
t3/d1AAkBkl/cu5YMB1vGfQ/bCUqkXPJBS6TZF0N/bHpUdVxQxHVz6xSGg0IUQlmrmtTK2HpKvDD
tZptxL/XXPxk+hm+0Mc1DJvPZO2bFTzMFyKNkd1uDf1lOvQb/b0cIBzFXT0dnbrbmAz2qQ0qc2rS
KXdauO8zL1NY+VGx16tR6k+JThf5qRQOuMzBwVMqYgfPNDSHn+IndQM9hWCqvEuuQQ33Cc3DVhi6
s0/W/TYIIbssZePHUmshCBWY71WfSou6FKQ9HY1dWBgQcratpTaZDqqhnBzb2FE/Y6kZ5FfdlR77
CZjk73urdhD+TiyaI7A+f2yS+1ukI2d8/PD+0m3ctDzmoYCOU35VaE6ruuF0Y6RoXKrCVnjyQ1W0
3pGlbvzUvVG31is/mwju7DzX/AqLtR3YRO6eAFPvRT4PyAugWOhdOpMH95An1YLnAqrHxXbmZn0p
q/eiacLWiAFixHPN4BSdA6By5nY7HZnbs5C9EHF2ivjmOLsAaFH+Yg80o2aNUVaxjHqm4c9O8V2g
K/2wL8lTgDuiBs4Kn7/TGfG+eEZ4/HVCaVq6SSflx/NQfHx2+dhAuSyik68Ne51pH7ZVJlobSzrZ
5uuIbaIdihNuOMjN9XbweW4EKvTu9Pl/tVpGPeRJ40P0AjDmfOXkXoN6hhbv34f3LBUtkGF0h1pG
Z5hXgi2gWngKWnueFRVKLMTBKgpKaKbrJfqbxHg4CJ0pEoRqQs8U/xAZLf74KOtG4fBClFjgctJ6
66MHlcW5tvYjPpV71Nnr7TXrDOYAcQbffNl4ZYOCHOxf554/gvF3zzBlQBO875PTyKKe+CxFM3Xo
uyIVun0gtBYqcz5HnZobQk9QnCn75wFmvm4pApo243BcbCqsOS7udJ2EwrpKEBpg4Vcj30jxlvCc
Op0aT2eikujM71DNw4P3xyTkO+H6DWPZoDMPrqR2UC2dotbUkTpOjtw2uRryFDIlLLXV9PQNsgnA
7cjM057NRg1e7M0T0CSdAY6ODM/AFZWFp/1Wg7YgslEgcZ7NPtyGfMb+pAt43HJD2omA7pylkoIK
jox1SuXJx2FrwZgPf21HSulWI88XfBxMvFeztRtI5GhWHRH5YAHOjRMTJCaZ63HVe90egOs8WKbK
SwN5paDudUIOTlX5b2DcnhnEz5fkdJsw6KB4WqUXfUy3vtiHxUT0XAaJ2FdpkaP9Qh7YzgyTIbWy
k85X30HwvjDIe6Q1Qa6k0d+P6F+riiU4WFAMZHbo3RTNzvT2QiCR3yJP4VTMkDz65uIx0F1fRCac
zrglI5Rq8HcxrQNs0/3jRuAErwEGxq5VdiSu1cZt6Wni0PIABfm2RIctgPUhRxuST0RZivUclqqJ
suJxQuIVLy0EPRGaPu1thYiiVRVoLJoUtEAx6ezaxPjEs7tvGZztQBPn/DGzLDP+Zc6yFg9k0p9R
/qI/eRodjl88KnHtvQ6Ps4Au4Y9Hmypy+8UMzjtAngry7wzS/rU59tpANVpOQDB+/JwJnl8NeIge
ioW6eQSlbWTkXa5JD9DxTOunsd5+CrhonUny0B4LwaDx9wq5LJLMlgwGkFyQcQjdDCVmXGCg/KVX
X4HufylCJAhUpzevPj1wDgFfFQXWw5EZPFkQOnfDsArePi3Xy53aScBjn3P7jItPz4VAN55pUEIK
ZuNRWMGHzOdam6FJmZDjFgU0Gzr1/4Jzw6McMgmb7l+P1durpfzVrcVajKBMhALIIZzmsTluTSn0
2lYZN0YugeY4S+nsnMwRXKoemGiAe/rDnZES/fi1RnXh3l/1EBTOCqXhY0rBl2NGwZGreT/a212P
sQ5Lx2sB+17beBoRtOMc0bgoUvLmFw4yWV3AnDRtqmsyP283e6RzJAScnH+u6SkgYNYuCqBexHg4
Rk88VC6lfTnnTNQNT+ZwJZC3pbGpOLb38axjAXVBf2+iCJhoK53j74UNjIRgq+Ko68NduFWkmUic
fjkktfAK3EVSUnSAd3PWt0P2oDDh00d8r8WfdWXa/Pbzyv7AWyrobNzeUiWgjxPOEEgRSQewVOlS
l2udMLSne6jyEpqsEbOqO7WN8QPhbwfm2tkDwHD/bpMdDFB7/13lcQ9+R/qfGsV7ngyqmGCuHx5Q
WUt87ebFkDhs2abNi4ZbQsKTurPlKcpgb8OQIoYKj4CRaJbvl1EZLHtbPGdDeErb7PnBiKtH/OeF
KEoEDGWwrOee9V/po2N+ocbifyu74nyRSwn+eolt80mjOFZbjC8wA/Y0O64RMmq1GouMcNBAjHRx
nKzn7do5bqHTrjPNdgtQc4noSL56n7D6M2h2s3OYglZOxT9zWNGzxvq0DSEUGh3F23X/+GTQm659
zdzt2I7/skcoI+AbSqLPBhDB7DxTdUBNT79JlYY1CODm5iF/Ab7y2dPCS7i2W25jhGoxfPfXEK3J
81XwFAmsyKcJFPCid8iewVHh7tep778sFqjpWS0MTf7TJSwD07PnVYMUY/AKgHMouQdJ7986uDVt
t9/tr/p+ZcHK0f7vP67o/g6yQQ6kiKPOfbCj3FU/qzFpUnXcAdkMR4LHKl3IRAO3Cu/emm1AEt4c
1u3Dv1siSh0NeamKOaNmbNwt2GFQEd4MtrNWDIa2JF/mloP2ZdZXijk+oAl9+CanXqPa0kTsKhrC
8SVWUgMmJFFuJu2D9du06MU9puij0txOcXL1JQ5T6UWQcY7OPbenLbo95YO6AC/ofm8onzwoQ36d
RQLsw+Hs4Ryg4UmUX0NT4pFIqthK8aaP1ikTBz+KOaYsgQcfgZdBIdEhnISzbH3Qt1Iafpg1ClVh
4tWRLEnP4inIVVmqu1yZ6T7uKJKFTaQ7YkOqIz6HjKsKJQkgve8qiCRTBq70ruJJQuj7TSDm5k0M
vCRcRtbGKvHSNxJzvQdlHrcFcnpDimhIIZ+0YiLqItNbSvEQAGjlTjE6wf/gOyapnEF76Ps/I5uy
aJH2OOVoenPHxlMSUt6HjNViKuUy5LOvgnTEJJR/FlEJm1SzebgC7PuAMwtrT2kSgiod1o5SPdBy
wAzffhPVwflBFN5qHCGnbCLxHdPWc1JnPIFsijvFMASYXZfzNyxfOQO7Yenujq1VXL50haSblwp7
koSWRyLqB16ZUpIfbgUSbWjNhAR7WrcOMOkjIl1dZIlF3r8Klg4LXIQ6h2PcjXt1cVyNGg7fb28T
yfnLJ635rsmdUVQk0dvurmVsmk6DIFdik8F5j8HXVHBaVhTCqIP+1jaMEEVIlVZNkd5T9NKiEwzx
JYD/t78RjMrVNNP4FfU5GoZ2KjlEnjNrU0Jwmy0OFPrQ42EkFOZTZegXxqcs+TU7dqtR6f+270zP
bCga52+CxwB9B9DaYnTwab0v85h+z6hmD+9b9v9YbDXUuxNazThY/GfgXYokvIBPBj7CpDCqN6Gp
wFi8fuxDVnTzHwB2g70258GjQPzuX2rKfKOs/90elVHQU1dR+yeHGpZ6v1eTrwiIRNCvW/z6z6ce
j+bejQ/x7Nv/yeSwta0u1iaMaI+iVK8AgodWf+70jaRCQAXfyKSFB3S6BZjmmTnfHhZIBudh6Zu2
lHpaNdQyh77dbWZTIRJq9sABystXm0rUXT5lG1QNMARu3nZrqbTaxu7otyY6rHSei9lEPDDDoMSD
hHCIJtT118BaHmSZKscxuNujNXZFXkawsI7DQ8dXM3DEyy4CabQY02B2XTGxg3AOAn1KZxrc2Tgj
YnxdlXNIRLPtScn6XfMlrYXkTAstV+PyTbMB1swpYigx4nPhoi1LawUVFoiqgJr+iBk2aM/puzhy
YvHu+osF5htmbVROIBAL/62pMZp9BPeCNUosz6B2BmseAII1QFvOl2BCPK1kuPr2XG9EX87evEAS
nWN4z48UtmThEgYzMjKVdEdUPCTCb6BD3idOggE+9sQJRmwgPre/n7MxmU7uGStn1C7ENwA225mc
0WtNf6EXyYsz6sPYVT2ZtJeHrE01ODXkqiYbd3JD7Z8O04KN5Mq2g1iaJOizTw2UZGTP1jcaRjHN
gNDPBZPUWeinDYrpZ+1DVWO9Go8kfnpKhEcItieQx8Y+pQRaG5kp7vaVg8ruYbtsO+mLavPZCrGE
sksZw1I771nJWBpWC1GVwBu9KuPcvbjoHHWOewRG6F7ClmctMUIsBpQ0mj6W5pXsSLxK9S69RgUO
bxXETCFZ0icLBqXUTqX2q0ytwqc7L3Ao+rkwbYo1qQhZfPIQiutUHpBmBfDv4dM+06D5K+fw8y5H
P2yZpXVYH0Nu2HYour1clFluTIF6k5RcsXDiqzEZFwQt3AYL5Hi96iDYLz4RTrVQe7LsH0iQvMFd
rTgF6+TxhvTRJjH5w6ZBhj84XLkxyONW+B0wBdzeqPZ9ndSXXJp+h9Z86RXSQOW8VIgRYbDCxkRC
Xj/bDnixybp8V4e2q/MXUo8hF/GJMk9cX82uvPGpVw5uz4kVNSZ7Nlsq7FR2AzcG+q/2Zeg8zD0g
DeI1jNFRCnG03y7uC8AHBp7yDsWZvOj07uLPkjarTxidLzMejImr7SW1VZfLrFVFaJjo8QiQW7vR
6hN/25OtQeBKMYV5WWolitk9/7S20Ix6vdOf6i1+DCKq/nSfmWvTwXM8Gdq5j+OvHwaIU6EYWnxv
dR/oHhqFpgjf9eM6evE+h2QrikAMj4LgnVRrtf7LGWABBwQ/hQbQRrgrvT9WP4f4zZaZjs1kl5K8
3fOY2IHgV+eFuWPRH+GDGrgsyJQOSZ+3qzlHYrM2GDrePi7nD9Ho5RZ6yyOenWa+dGkN1D20G2xg
FsNaSorrn8TqDZsvHBZnwvyZpyuQHMIvziMAIOmCDKMzMWkstgbyaroor9CMBpMxi25Dzs7QtAl4
6ckzuEElAfsW3rMj+FJgk2CN2fB8EZPN6WBqP6vOeFg3QrsPasl1nbqChG6JGS4xnQV4pFgz+k9r
vM4teZ2EQXeUZxVMDBv082TKwRrzjIRUcviNJzW8Kj2Z67HabeFGaLJVHC8cMp2WmzUK1pv1Yu3s
seIxjky/8nPCl2qwQnqu3zcJvod3QgMbeJlbDD2uLsgg0GWGuZxO4lhMrBp28tS58I9zmI1leTiJ
vEWWmnJ/GhGTbOXSxEAcjPZy9OLhwF7P5RyHM2MGcStBdfmz4OiU40usvvvuqCQERlaxb9Qj6CKE
spTn04AyCvZzV0XPkox5B7+/SnAszqJVgoli9WG5pEmzAyqpSWvII4gzphPGRGej8VHHohvQHR1+
SxZCshFyl77vC41lho+UYah+D5odqTafDO9lQoCJbfeUvX87saZzo8ubukr7dJReygMeIGNFVPQA
BEZAtW9EECgeNMsmKX22VUnMqnuusIz8TSgZZcc8Rp1g3HezP4+CIAZvkO1Co1LX/4i0S9o/TAjR
tKyPKkh95k3nqw00VjeI2aTednGK9b0SPgWoFNgKsDn2G7/EPuUutDs3DTkUR1LdS5vLiNy9S/Qm
f697FutWD8qzUROJu1xUo81QF0nZ50nL8imIIzeqxed0S8JzFMLXCXobMjvnNVMd416WYbxgDAsI
pQZVT8lymH0i5wAbm4StePMSeQuXWNDY1e7yiMuXczkI7TpUt7QlZWyecFg8HLULzSSzDSW1n3s3
Yd/EqbimHf8uqXzCrdmXSKYTLtKLSWlYb9wP3v92nLNIWOr+iW4AKXMWBW4oJjEJBZ3Du06NNdk2
kvW2Pij36xdDyNW0nMC1m/bc0LOnBcQzqUXZbz9+LpRYWDQvfseyN3HIucjteO1Biq2aogtYNPd0
aSR7XMXQOREEcIUuaP1556xa+ZNbVA7U+buF+SVRjesfW8jRHXXrBITO8O6gWUpY2g110MmTobjb
EES3V5Icia4/XJWsm9a0+/0k7nNVJR3cJ1Bil8yN3yw8zF5skdCNSHjjnww1wctXty/bLZQIgB2d
0bX6tro2l/YfYJBZdVHmwLXc7MJZ6m+NDacylg1yr3n4xWTQPb/zwRryMPH6/fBF9Kwpudo7n8F0
pqeH0tj08UGk978iaBH37Bf73nVEmt6tU0i04NokXQatzSC9aS643LxYFfRzLTZAcQDEkfv+TbB2
Asarakj/KGtnxHvATwmghMM6KtMH553PtvxvzmZl8DAMasIQjdZvBJn5PXUCK91zWrdv6C1RHyPQ
wmQIrNjxGEy+5ouVNDRI0YhL7NSsOJ3U7ULgLB4gmK4pRAH/SPkuA7/rbc84MEnV5AlHY0LZOoW1
KQPsvP1zY2m8xc5CKD4dvX02yy86mNfQZNwf2wN6O6S/F2sFMUsFdAbVO57JL1THIxiPXE0EnXuf
mWzD7jJiFbSBLFVxCCC+GSjzJoPMueXLkSMCLBpecEQfnv9UAGGa1mvW8aKulXkLtrExShkhLsOU
RiXdjCJ7CF1eBluLU646x3v5tkOWsBq8AX9DJT5zk9uARFcSLfOI5LSBkTwnezCCsD1Yy+orDLjd
O/CAdUd9GIsq8I7vO1ZfxX8aQ5znMBJai+HOR/Y4DZzBSC9ykU8+4sIIGeWssxzUkBJcxU52hz8y
pybm73XHBHq27UwSyCKOhNuD6ajyjQNIiqPSoK+E1Q8as/t4R0Fw76ikfATVQL5FgBk0glpNJry/
Y5G4nUEM0raygC1Jm11Qw27gLZGIo5XE7UXOVDNKpvLs8C6q9yckjXXjeKNPJ+Qkcb4r+lMff8wT
jB2Jx+KXBcUuF7nUC4TDJ3LyWxh2KsiNB3aw8BMdYE9d0iyyn3iahy8+SKvO+fv9g7urnNYVe02O
CH2GPWe8Co2o2uZELE+nv6ww+SGxMoqSU0s86pgl74qA417PvEOQgRBaQ8eBxMmqp0DJMxq2gT+i
W/v1jDoceePvhMATR/0Al7UkXSlejI/yULjqTJXgTokGIKo2sZxQNPtq5sv6ud6NezGK9rVgkmti
iYg7q8Cml0J0LEeu3ADmPpWKX3Hp4Y32FusHKH7h3ZeURFXn39t7VFqvdvmrEmSVxPXGHwA2Pw4S
nMhuMe4EDDGJC5t8Hx47zIgQuxdTBqchbTyA2HtMgPu5fBHlyQ5GuXeRB6jRhRfdwUQiME0dajUk
xWEN2mZKUYt1nztKDtd9l2iM0K73rnNUnqBnF0G9k0E/SvK8D6gXTrXdJbZ2fTXTSe+02I5I5a2k
U4sVmi61O132NRR/ZaQlBkTSg5OAwssJt65uHMlvUBQ/BuMXAVpKgOXGX4lh7y9dHgFMcwGC2MCk
29KNOGUbIlEctRMdBZYeI4teqUc7dzDWnZ/w0dWQPB1+eefObRoShzDP/YSRi1gTAI5WnGFB8nx/
rVdJGi+60vOq9Se3hAD3ssbMgAN2fQrWzso7KojnpaqwdzjO5znbvCrl+/PTmggWNNwOxEb+rOha
Slnsa0VBNGg2PC7W0GqUzWA71eMeiWItaRiN6K1/g+copCqu/9vV+WPfUHqA/8LBRAY27RNRqxrX
uME6poWfM3UJPJM4F8uMF6S79MA1WsC2oty6qj7peNO+I8kftGY/ulZVxihfy4N4vmc7B/hocILf
HTaOBYRznYcngA/XFsZRX9cJJTYTnBeblx5c1maN/gPBClsJp0wlUWMrpx+wCM5wPK++Ga3B0aBG
a6HNe/8bUtucAwcDyOAWp/OryB5DCWh3qTJOJjJZ+t/eDFD3+zbR/eUVLAllCEmtgdadUF2mmzeR
4rrtT8LlsZfpGT6vHYZtMcm6xJz8dCxoRDMglDFlGmEqleTx04c6rLr1xU8PyR4hKsJeetYJy4Cl
6SgXvi/dAdUnWglqEmOrDMG4WJmRZBzK57u7S0hI85y3wsNRdlGh7iXvLwskuB0Xrmz3ca/gAj5U
JaAp00jDqDvBQBuvzvLLuTXV3Vb2RUusfk4AEVho/xE+dTiZBHJKCxMDjCKUrhifG28tOc3EPcR3
GLXB68B9DUQKPUU5jYcYVztKVMpnl45gx+AHBeQ2hvyM9Ec2ouoCY5g4fEX0RQk+ZjKPSkUNe6mq
Z4XtKQ+QP5rYF2Mo1sgj1r+D7by2P1ONTIGuvgf3hgmdGeLcmg9BQrfOTnqpgEtmtD2/2YI64Knt
GsAbnRUsJHzU0RXW8AVytk8IEdHd6eOPGerBy/QbKNByl2/bYyNa7OvqDQP8xi6DFtqFbxqU13mV
2ISS5MSEA3i/78WDrbGBf+DKfYR+rksAkP/nyi6PIDnaKmzcXIlTYYVZDOp96E2q1G4kPMnVJGSf
wpCxipV57Mmn4g2dSEPhqqPM9T2ZsAg2PldtAy+D4/rKfeVcehJYkNPesfxWdtFFK56lyhHI4Kox
GX5iSWIuL92d2xFXjVIWlznaA/xjB9TldFrlBPcIV149RdkQ8Sx6u4OwZuhZdQ9N46ROxVUjE8lT
IP28fhYVV0QVjA48LZys1BXnWmU/VW3BRtCHmFEJHrPTi2ix6mRufalxbLx40cDQuTxrk2fFTwNX
w2JPaHrOXSl24e63Iorfuhs1m/KI0dKKLKkipJz1k5U6Kawge2EVdZ5JTpR6oEYu0dwo4h5P+7aR
Yh6A7kmeftOx0vmz3z6XnAXUWTeffnQM6zeGMQZOUSov+cCrn+Al6n8OsSy0d+Ir16xnOOTvkx6G
vdulftsdG4TuAwVKjmUs9ez7E3NqqxIflWWS4TNtUJXwZqASuN5HaJ/lH3f9H2BoREdc/CjsSloM
n95Kw39NBNBwYajeNDn01eX3hVF1mjClUe/nZcX/fwYHk3pz3VSsw5yOouR3VB7LP/T1ifdaQ1F5
j9/mkRYCca7VEmwF4Bv20hYFh/5egPK8o5i2yXqm7Y4RvPLBsXm1zadDCDMnhcJ3yWAToK94z9ys
Ju2qpvYsAi4QNMsbOd2B1tJEgqnVrCRU50wL+Rupl3u9/yDCz/DVoqce1chtEEeAr+YAb9gVLddH
67TU5bmkLOUmmC/yC3NCzh7BlTJgiMVlPXCpmTGyfUs4QMR559RFdlP/XLvGnBPkstmJnDjMyIys
4GC2Bf4VFM4xsHQA0Bg3t/LCYSM5fcsVXxOsciLGm+C2piYolWjU4R1sfqDOkCb/PBUPduXFQzoH
VIELU9865560HyfxBS1OpJc16VQrFPHY24r2PJ0nJC4gh3YUDp9xz1mv0Y+VF8dgDniO7t7RGqEn
K+vQQ1VwEVnzzftEnPrjb8/plsBTGv+CI5/KwcUnZ8xrcC+gC0IwWvtLfY47kZUw3Bi5Tzbv8PkQ
y0dUd8ujLYHNylMcFuwy9YT5O+N8ybZfZZ8IzUBLGd+PEH3Do/H4mWRStk3TZpoSy23sVGY5FCgP
vgxe+enM6ly/Ugd3CcUAk8KAuTr3DxCssoI+xbHqdjF2iOvkRLTdHxhmyouF++JgVnL0rLzjdX8s
QHTo9hkfr5RCETs6bh+EtEWmaduEd2s+E4uK1qtsX6vFIHG8mxcU8KX598M/ecoch37L3FblZ8yT
iu8oza/Kdn5Ym4FToXsiOOU3BjKU0KUbCdKRNAXVyd5pVQp+ZYCd14F5LC5acMwDS2iGN7z2uHDf
54vOgdveCXxp8Qr1cmBNTZzgYK5//uI2CsbCDW6zhQ3Kfta5OkCILoVT0uHJeDdO+ZvT9nfsGAXy
L1qwbaOpMgZr8ZmRLNN90/VGMjBvucYhfbCNMqizvd4z2dk655J0fJSBr9EB3DgZ1x4oc6La6lDL
zEejbeikNSur4ls0tCIuYNUKzVkmCwdMgQOfs/p6M6rJIKcJy2MeDLbLVa3g28nREZ21QR88KwA5
3iK0TWzzQKNTH3ylhHoy0s/Xpb6BU7xZcFVjQScUvzWZROpJpBiT/5qOZF39QFPBsPRfMki7nMqj
gvlhdpzOhDcf7uL087X5v6uhaKFh6c73Yj2XFEhNBlQvZe2iGMYUdzERdPIuiBCf6uisAJwKGyrE
vyNkTyrDA030mKWk05s6wynOk4iSBXXTdenR9Q9REOCHMftDHBhAmvp6RjtVS9AZrJf8RR8HcQ3c
cmnbGKlLeD5Jf1WjJIaUy4b6u2Hz/hx4ahiPIfgRAuQPJxY2QFAUGlOOBpMtOzBL6LeZWaUgwKel
1HXJMeLVflkT5Hd3FULpl3aSc9yoEzIXq8RxBJDlCflFoMHi3PFIzYhS3TRGetYnMR40tK8E8x9n
7d5HCkG+u+ckwr6AygytWFCsD6OTW++AyI/cKDdNKKYs2UewY4lSZF3hG+kyDiZuVvDuFzX6M+Os
hTQHCjVDip2gFIEQnzuB04cNPU8sKOJKnbC+itEXbaL5pHKrgilJwWSc3MYt3Rn46dMh9jslZNke
soiqFUrKzXhIA4xYRDeAALGRRlPNbNvJOsS2z4+AD5MLzg7v0HZTPfL3af1nvYGHUZkLmJ1IO3QS
HoK4+1MrWhO/4+9fTTWzZfXdF4UEXpBrRTOU5RjSJoDyR01jG6tH5svB3HqEVcJgqY5tgMoV8L8y
UDF+qd4XRYhXOSvLWhsWQZF9o/ZO1Ika70VVGAyWL0jykOJuJCVGossDAqMR59mqrRSEvpk2VU/6
ausB6ZD/9FSpklIaVwqgG5NhTkKMPG+YJpHxgrTNB/3CRGaTK4jkoKUX31HTY6GlwAPtSry4LjFN
mUI5qGrAOeIEnr2qSPnsrFaj2RtWYwQK3+aoUj1QFj8yGvvtJ68l/1LaQCCHfx/NFPBgWo6q7vs3
xYOxwvIArGEYzN8QZcoqQDgfkxjCz4x0RwdhgwIfN2abbDlUUBxnnOq4UrldL5lEPzOX+EhkSMfB
aO6m5ilBEX/xDrdbVy1ry62zGtwLnHrnV9J0kKEb2fBmzuSHZ1konYlmeP11/4bJXrli4AtNZbkK
L03nBbv8KDCjCZQ+/iLhChjTv6UHaW3WTdtottWPj801y6yLb/4VX3J8MMUXAxQYiNfV5swnhhDX
+j6PfyvVqMFqDlZG3sLUpx+KxL9IIHyqvfkB3GXn1gyo2KWn9HnK5r3aiYSaynfu6CCpUpbqquD4
HO7zwxPP2fOzUy68g6LKiLNHRcPEWXg77v5nwjsNZvLcQqiOxk0jduZIAgLZWnvVVC+mgg7IlYHF
gXkkbiSXwlf7p/txrNMWvz8uBXTdbjVuNmldTl2gFNxjsXNOSWVNtRBPFNEsHMM+upVOkIdsZuaN
mas2FkDefgYpVnHDtaj3lwXJ13hbBoWmy4JW6DQ2rPOkhu3J73tVAAzq7A8zoxXmdzOmH+Fxs+Ux
YYylewwnuYqD4Ljd6C/nS46zWE8hvALXK6ePwugs/JwapizlNOiEM9d37/QtJ//JgdcXxXt8Iuym
5B+7qgvUtfBZ5/f2Nq/U0F0prh8eSjsAl2Vpm3/6s+DQoMOnRlpaeelhguFQRQA/fBhOG7rsoM8y
1V2p7goE2MlzULQbPVBGZhBfkiVkb5aRLg46vEBueKe52teZn80AhNCSEaOEpeTNBIeKXYWjLaGz
jBkZObodLcjhBtGZ0Mcq60jn6O1SVPW2x3QK1RJOpMgeIvYx/DDiD7pXdbZqaCixznuxO9hxqBBh
KgPRuajHz2igSjGTzpnncxoviZRa7Egqt3EqMZjVHPr9DUBXBIvBBvCqknodHxiKaM4NYVF3UgMD
r2xOrWY4OanOdDJzM3p1APr9VBjxEfsxsDpmW5kwzI6Lxd26rWO8506hZ45HzQoQ8FAyJjuzY7tn
GhPv0h/7pme57yZT4hEQcjUaS2jb3Objbf30JsaquYrbK6+vy/yGnYz4UWT3sLoo2QI1LbAPiT7u
gy7PDdSW1Qu+8WMrUZBebx6dDtJwouZ2bWmCx2Aq6HDWsAjzsJ2VNai21eIqs5z1txdnSP++wwDo
sGlrFdwRR533o8E5gE6/FTIRe44EInZ7kWUIGRjoienkMCKWQgxH3oDIm6a0APe/wa1bxXhLpE4k
/OkWmwZDqn1JJuSn0jwEADSSQMV6rndhgxO4f8POAQnmHbS/v9GbowMS6cRqnrbNfIXtLbTl+2VB
Y1OhFZEMwGYBImAmnFjhnhuwUdMhiFp2bVX29n/iF6KKWMStxYXNVqkDOxqhtfMThMuUjutI85vV
hKxtXtFU9DjsOq01hiev+ELqe4J48KrMEmR8kwVKVeuOP7lINrwCyMDevMlRJC+0slqim13iY77X
Ib4OXAadGMCIUhtmGlTJPmdOxXm7HGB4qjIyjQmg4E1Z3nW96J2dr2STJgtfAbmtJChcWY1S8eGm
EEgFqNaaANvwB/jo9WoxnkeIp9MifQIgFBukAK8sJm78r6bVC/FwjTtsalrT1o63Cnb4hKtZrcGn
JruOIqimWH+O0TyhXgk7pc0mNllHxQ7HMpA48EJr0B7C4+Hxqk5ycIV9o6qVbJj7KB6Hh1ouyTaO
UI0VO7t+wjMtGOuf3gC5e8w2AuSP0q1PJF3KojkTLhesTc5GlSmJmiQ5juqNzoBxZdasM2ApxuBm
wnbzRxU5o5u9j776u3qxT6W+HyBqH4G/cRtd8duMaTb+EAPHUyJ2XfBaS/K13Dauuswj+eS0tXCy
uIscvQdsYHFxhI9SpuyWmq+O9hFN+sOilZldgzwo200RFRBNsb9+zPfKWHLTFkB8uttE59AlKUXV
zRqbbeqn1pIMQF4tRLPfLQz2NSLrz/CrcnCQ+hK4eMWxKSas5kW/zDFDVVLBd/3KG2VElf/92c7a
rwC56Fj3fcbfsgG1yPhJZ5Ry6QKwRFhHMIJhmaCy7fqF+pUs0nzFngw4xQUcIbLwV/zLkaGouOt6
WoZCwCdqKdCjh9t10qAU7Y5tlzsbtvTXuklabcCp2xpMNA3YWEVQmUITvLVOtTvdebcRKLsIFiQs
MnZBt9/J/cbaRI1xX2+kiMIyHD/eawAYOPwpsTDGbeWu0BZUi4puCZVk/9RCE6xuBWRwo8+k8uzX
SubdI/pzTY42A3CJKEKnDupDl3nF/d8yvP7P6EzgMYYKDbaT4p7rJ3K8h6OxOtN0tDdvWcoHP2ar
we8MGhh0EekuQaya3dxOZsms4T6gE7DE4+w6mi1qdZqVYBmxsKM+W9im/mnG7uI7cDxHaHvITOCV
cbAtfZL2NnvoJdafys707oCUNUbid4rk0/7k1xJK4Y5N5BCMKg3bywDBJU8XrWysA/fxTVVuh5sV
cUeZCM5JGl/IeKeS6MPodGyIxAAGjE6zgSpUM1sFQZILwlvIXKRUBXdI/Xi0n5TTYy8Un/6beXT7
0vLocXB4GafOur6+ckGOeBN7MlKaT8eqjfD2pfhXgT8F/F/veFg4BOBR0Fwwl9HUQDnxd2vAiUQu
1nFracgzrh0mtQUY78idWMn3HJbD5b/CS/28wWrlMGpdT3o1fxwnffXcQXs/lLEXEsUMBy9juUYm
c8xTtCV9tfvrCzpWgQEedMRozJ/O5pD4ApqjrF6ZJnqs9dMNExssdd5++RWp/TLO40tW18JdwTgY
6LuX/0HC698+KFKKXnJducgKnhdg87lQB7OMet6WiiM6RVKJmh7xrLmsyU6Tb1cZIx9QTG8iDSpQ
x0aIQADjYrPDWpnPB2NB/rQJ6XiTYrw9kDMGf0fPs4oIth986PsrFBNXtEVL4/f/3IvGTJ3WYjvW
IHppV0az7iMxxfQnMBwjCUM4tAezpfdjMYW7ju8ZyE4BLiuV9qku7F84KaiZXc/DW6bnErQMy1dn
twF3qlhSbyuBDHQ+Hmut/uYkW1fFlPg+hTJfFXdF9HJt4BwficQto3D8vdG6CJH0Gk1jdpnDobO9
3M4lqlhZEtNqy0cmmaVGgPnyJPXgouMAH2EifHZhCljZx4HHJVzxhd88ZrSaw5xIWiWIeoM60/Ex
9YVVzyik+CayHAxSYOUByHgUFfJh5kQBpoUwpHrgSX6gquX+muNmXkuITdHfOAdQbVXWYz6KKMmZ
iNyDOWCXwqXxMCOZzHaPRl3eDkhY24/JZSLRFU2vxw3OtWmrck8D4BKRX83VnWXieVJVm28k1m4W
Es9WrilroiUMo4M7g67san5NqwSQ+hjGjnn+HYSR87Cw/taWcpfhLSfXzDB1nyfVBPOnLdM3uD36
XbSSDtr/KdfPQXp/5fMX4JQ9Y3TKz5Fbca8Jgb7F/F6mGjVMpmiPYhqTp2gxY8xxjSe7TxvtbUxs
U/2k4tUBMrXAPoowzAi2aYakR7kARqS8/2HmPQrN7bZ5OrE+2+cMIXTNzDhldkH6G3cWGw/jpHYx
rm2vfbCmBotaRflHe78LTs7KCBOQWalNGtrXyz86etgJ26FeiRBQ+VRENWIXYfKtTNPR2cTZ/VdQ
dN74eR2ILTtduDgRK1pF4NFKplPBRPlXA+JoI/6ByAm66RoVYwXi4o0VH13LJcjH5wawC2JmUf/6
HkwvmK9wrIMQmBCczSMdE6PMXsZAuYeNXImUUSQE7WbBlLOFC8CWs8ZQ/iWycGAYXJwVLM3Ff7gf
CSMYA7PfJsMDFM+eKFsUT0I/hym5N9puf/q6r3sCYDyi1+9hRXuhumCHo/FSfLp4fVUaOrod6rNh
Amk+k4tXvewegMCtZuHrm5ILzHHPkNIOpoLz2MRc3KmitaVBHFvL2WADIfZXs2vGqYuvzSE3uIMM
CsUe5dhGjUEVNRJ+8EHqF0iZZjiDjoTHzuh0r4KewIrNZqEpMRurBioevOPHaGkKY5f7cdqnU8nH
9YNCbmoOL31Fc2VcRl4G6le5OhCjcSaqbaN9yyPhUMDFdkdH7jjn6o7CgcBuVTmKowVTRaZBOK0g
UgoFhmSn/tpeeyvLrXCSqoLf6oyD5/z/3bfx48+Qn1LAc+GAyun58yq7njvK7mUmpMqt99c1IgZj
vDB5xlV5an2K+OyZl8cS2n7gyrn81FMHbYyipHGX6v1qjlEY9Eq3iqjzoN+9PKOeAjJkv6q29QQZ
x6LLGzUBkjFd4CWcrIcSlKmcg/6dyLld2hKEJ0BYGZ3ujlTxm0hPwVPYRKcW0SotKuRBuKg4Vp1O
xL2Mdn4Gb1sxlt7QDROGT5VC85vMDl3e8U6nCCOQoYP4lKjZkE1yn97/lCK17J0QoKRc+nQJGsE7
ot+r1QW/Lrh/j8hVYldcwf1l8Q/yNoTjuey+wZvYNIyxCbJr8kjg+Auc3dYj6KFzrPm5Xfln3xot
dQ19yNXVQR+oTu2sRgnYrzaM3/huzGq8IqGk0X7VpC0uMOaf5ag7RnYW3aHQZMaAH3KOIf1Ggzaa
iXywZtQFnigpuQSdd9f9bmYwCxR/sN14R3oITCTT07cUe4LKESFTTnFggnjiWeOC8yFo6ypmwvBV
mfrS3pArxlqLvbg4MIsfmK4/DDrHiuwSmxu2IcF2jWZ54/QdWQgP9jLSQbynP0XvE8lsA0N+l6ew
3Afy2wgFN/4eFECgofHkypTkp96blapTqoZEVZT+T7wLv7H+bhGeobHeR/1zQP66Q63ejLV8Pqcz
oStUWDQ3ZXVWmDaHS4ZoAw3jVbjDytA0rnYI2Ai8ZFVoc64eNpoSC6qKPSzbeC4x9/vQdZS7I/CJ
CI8iYUEiuJ9jx6uQR5om1z71CQ0ocs78GdDR1va5S1pzP/VBF4aqwLcR2Zk9QM6RcxIC0lWUgx94
UcWpXK+1QHh5qg/XSPub1XnFs48JEpyQdqZCXfdi2GZLmtjUu17SvSihfvbg3LR6p6kcT7k+XukJ
x0z0BVXbh1Nah4+XeFEDssCD/RaeUzwhq6GcEUQ+zZ2tBtMozjadmvuwU8LMoh/LTPuXBSMihWXd
vMhr4yH8nUnB7azE1jrYYb5QX90yCchiuQHq8R+9Mn0JyS/Yymu72yoNYij8/wonv4W3kq8+Ul8u
gRWfQGv8oI2KMrOAV4gbb0ly3eYcF0FxbM+aBn6+Erxg2GJZPRszjcURrMha+ZF0zZpcShBQg3+b
PIWdZjIzJgqsuabTCnJd1ZhhqakWS+ehfSqILA5xJh0ffHfZOUPeTB9U/LbWbkNKb6blTEo231Wj
z7OfCewsihE7JXo7izPW8JVTapYDGdAgTG/TTYYT0KT/Jtwt9NU/XcF7Ykm4JuR6VbLo8LM4qw9R
pBh1jTpLH+bAHAlhhLkak5TtoqMy76RSEKJ52YRzQSVlVJ/I1AAhBZnW9f2mTrScqGvl4dBO8RIJ
g9EQy6WHboqA/KtN9k/vakV4aTfeRirZ7zd32NTfu5/opAcW+rAw9eoQVFXvrUuD/YuZLd6XNQAP
5SjkIENiFiZ8VVQeUMVQQFhfTHKv9QE/Mie8JGJBjsJiJNEZcFYsfY30tC8l4MbRVrZHdUqTZj7d
8eUMy9oWFT9WjVTovvUPFJn/7Kn4BXI4z6LbkvZG1cD2R2mog4RBQfCOoAn80SrX9G7KMtRfAC5s
R/e4X3BFhRB0OmLtEMD3Eke3nWGdZUhtDlDfhpgyuj2yHuw2Gqgdz+npwg+hXLwDrEeFEtYcQw2J
/cEqxFh7k2eOerDmyxW7l2JVn7KdhqGc8lHLcLqJyaQgwTZfjW3w8JgHFgQ0ojXZuMZrqRnYHUH1
5CtN4HVUi7jLT60k/WMhS7s+89OzBE64rkHcIrqBZAdt/VvgaJ5jIMQDeMQ5m5YEYoXnz6XgjJ3l
W82YVGskS8pbtcUTWDm7jSNdwbunZEomQ8lkQcF8gMs978w5v4GOqrvkDC4TZFd3CmgkKD8SADZI
jU6OThSxAaB6toDzrha05N0g34GMPzUSBWxqmGmtNJIV3TarM3S3al34/TRklxSMUkMA/4Di14zb
1BHbbQANUgtNJE9ZpgBpT7jaB0+ewQ4lS0GySa9vgVD7PBnV8b4P5Y6hqJhnlAIei4J2sYLQZQHs
SujFCelD9NyCDGlnMSQU/41H3z7SRPEagEekQuBu0P+CaIRKbn/Mq1eqA94e9dzAtNM63rjKXMIv
++Mja9yYowy4ZAkTXE69VLcC4P/sXDkHkItnUY32DlH2Um1mPA/eVtK3X+Iiec+bYN+XDzfSfTJN
5d755DowoaadqMQtYzZVWE01EOBuM5jEA31xzGfj1ZHfbZl9mtOxsPK8QZjyZsADOdBz8f5fAH3u
9jqQXzUatTsWi9NYNvEf9DzcsEveWbc6LfarqJucX4Zjf6NAzBP9xd36eItfRWmopg7d0yWJnbte
7F0AMB1eUYbVa2RtlLIgT00ZZFOQFSjM/90eG+fGHKvV1SLNkPj0N9nyxTYy6bxe1H2iz6VyqrpN
VhE7TMKbNyQ15EDJLoGvSZBcTmxPmAtPCYYYI5SfSuLve9cyef+3D9qYkLTJJDDUtABBfDDLacEC
R0Czs00w4oPNfsRtzsMKWpP2E4UH1b+YxHd+rVfoa6LDMqli09d8+j2EhfNQ1rQTTGx9Bh5uqV5L
DTAIS5hH7ado0aXmVuNF4OFaHHk00XyIaiBApy7RkrNT6rtSL8NFrvP9WFu02elQGpDsM1/Gblxa
D7HE7RE7W0qtdKyV3vMyH+DAmgOHPDISfZWvbT0o4m3rYyjcO5bKSab8wX3MgwLBYVvmgbYtsyGu
/wsnE17VFVQux4RBayHMbc7Z5JyE+sipvTTGb6H47BuSTC22CtATILUx7RjSQ+pjm385aeeZhWuj
xklSU/6umjicU8krn0cMGTry71+9xdZ377H5RjktAkKn8xE/lEhTj9npcS/TJWNzQzv1pofH492B
2ItFDF8xqk/whTy1EE1MRbGbDM1H4ZuvxJS/tB8dDjIr0w8mgpjndXo3pNwOSiIDSKvfoHXBn3Zd
4qCPMrcB2uqSiSOlLVxHq8JQ7G1ZMl7Q3icHsub5jhspDxRk61kyTjUFJlXqVGvNC6tawzoAd498
N2MMBOSg5eP2FhRE9HEkq3iDlLM7zqAdwISoSmrNIfVekZCisbMyuqmKjeHc0wzg5d/mTcPKEVQN
TlZ1qrGWKlRkCIXki0LXRERL7cpCvF5opbzRvshly64CF+EVN7R03E8wHsqZDM4zenIudFNJyfDp
fJdb2DXzcCDHEkCYy5L4UqLdhb7T2WRsIwIlAMnpWBF6MOXxTHvW3JurcGsCfb6WkiXFuBl1KRK8
2WWeTWYEILDt3RrL9TFD6tZ9RDvfRst9KLFXXFmCURkfOeyJbEk65EVe5vF6om+h960wHq2YaPWw
v5vVYpSnVLD7f+8kGEz5O/+zrXrSXyUis0Bn47VBSQuIOYtKLMzNLgFKi5H7ueFWj9e8a9TkF+iM
Lvr1Pl0kBgphJ2T5Zuoh+iFWsPlRU5FCLg60VrheQ5YD1jjfoqwpiK7cCe+5VdKCxobf/efSf4lq
f1QPRzMuR+/mNKc5/uXweWddeb4BCidocX9885l2g4z17z19jik603e7MyLohJzfjQF5sLyIyBx+
dpDZ9T1LtDre8aQr7uOhPTqRzoV36iWO0pKsoQ3uYrFaUBmU9lMW3CTg4oekDvQ3NWOWguQbhPNf
PTbiCx/60YbfUGABjlz5AfHW+P1enBJzvB89LZYoPw/B1X84ce4/RYnzynF2Xtox+hs/FCKDpPmT
hy7rwKXIHXlGFJBPxAVNIA2jxbtyvNhv2/uZXH1mqvAq5NJ7zvuPWPemisAg4LCNRy1BulLYzrMi
x4i+++ntDRjy486hhQVYQRijN3dPDiboqMo8Mzt7PCDi7K2Y2rpdy+HCJohFDY5NFqBUC1YyL80M
Ev/UcgA2PK4yh0S0IgMp/6kZ98eZeilpg847X01I9Y+/thehPNE8rMcTN91t/jtQiDcuruIoU4UB
5zepCMuGbpGZIDNHyL7u3v9WmlCM7n2p9S0DsYlbWS5x/6LqBfktRQSS7Z+RBg9KCfVfzbUy8Lcj
7yeujZOwJjeKAztFHl6h/q+jTmrZi8ZMX3RCT66GSFNTynCVSPNRiwPKbBY7WU8WTrLk1l+g5s0V
F1fz0qE4aEkJpGkd34wNA0QT/frqGKFlVkEH1GD9pOOH3U4UzDtWfQtR9fl1ogrmgSu5A61FSUHc
Z3HD0vNXhAp10iraLnZz+W/AWDOFxI63t+7ye8KXDe/h2Svo5XW3i3mSQYbL7KWrOIzW6SDWehlS
y5lsWzxc6ZMhlIBeY6FJQRH6UGzqHS+d6eQFXH8d05wttWu6e7rEyDnqe9KbIZktT98BuPXJ8X1p
aReDIgdEOqtZ23lqePkaoVuXBlLMegIkk/Sp9dyD+7t+q04mN2Fm2v3GA93/pyvlckdjBZRNyvvm
i+dK/HFEov5ruEtZmcQE3bwgb1z5y01CwIPOdGsOAuFfXlrrY08iJ/W97zeiQZuzXowvhwC1hTX+
8wq7DUNh5XK0h+lipzoMiDT6oQxSwolrMIDffD3UESqhoU8YYVxEXAd87WCKEbaEJ6MimdJvo1td
y/9Zl9oCXgBagq9NvzB5d7nXBuCj+78BYEh+yQCd/gQJONA4iLyui5gizGmo/r68aOchUsWmsnrn
J00uOWABRqf9fDdNAvMUvdY4SDlfkX6Gor1xqZtEHyYiD1AvKLmxjg0D+tYVQdsgtHF86O9FMA1S
sp0LrftX/p0IeY2flQP1ALkLP2AZZBVLcPMb2JXLvl7hZC733owFEo8aKOV+Xt9qmkWti5IqllOG
H/K+wIHBQVMk9w8cKxqMeTNwmCdhj8B8ffcSex6SVZLTFuKfUbozx5/hLUlYM/sJvMZ9QWH2NDk9
fhn0EY+dk3oZHj76Iv0fz0js8iXENbVFnZ7x55vLIjLyC3vRDaHhjHgtPdYFDsJtSo74Uvt7Q22M
+Mi5I0H/afMhoFwp694A0kHy4Ibq2ivLkQRcINJyNrFgOTcoBYRKArovQgjtNAzgIRDPpfW6RbJJ
wO4jaMeChduM2Nnp3LVT8tfQNzTrxRjJU5gMJbomGzzskdUkIjxvfMdMhJeElr8hh/F3PGDe/uuR
Uc5QZvf7TJY58RUnldeABZV/N3VouXWmkPf15PNDkeF6Vfqs7+hqgwQUcm7TK98jJDV5KEKuapJk
npBopbHlhqY6V1oaP+OTF88wGmESOBJ/jTieGPoXRqjETrmD1jR1IuzkfDckCVKnbmIbljDVFlKs
AFxwAKy/9WYN+qSWSWgjuPGiq8aNQgSUIxTUVYdN7Z4Gt0XPR4CwX9U7mfRODU9+/25YCrUV0a7b
5PnpbUOpdoL039VB/OB+R2E2Y/JUlppNQjmo+27fj5+Q8xaZKPQgMcDhQH9qATwuh9PMysstpUWq
oOIXQiO+5Ba2inKAMEXXiFIKAp0qu7eULgi2t2529b8dZCO3Y72EvBcNcSsatHZGLWTPjYoSs47L
o+NWczxpG55ERb+Ax9IVdKkBVsqNaR4YlaBM24pjEsOLJRjt5uCqOy5F+CpyfUfQyE7ZZaOzKL+m
0lzhXZmr6t8cb6Y5j6FSltDVd32JTyT1yzx6pZ1oceohhmM2jP7T4amaege5xqR/r+GV0UrL6CbJ
BETjg6WZ01t+TC7KjU8mRZnehQNwbJvxsOJ6EgXDwPrmrfRB46hoUhyw9jT6bh5m0mS7z5P5kFnS
C/fCHZdL5M8Y6yMbl5DveCfFs7qoc0AX4ys5gVAMyeN0o+2xNsMw9SG+jUHQFFQsLhOzPEzHkZt/
yCFA7pyfTzWEKaM8X4V/8GGix8oE6Ta4IwGPUpk+DHhH8D8ROLle45HbS33c7OJGu64LlEeynfhY
PgMe4QsczHgAdLToVJBTz43QZe0AbXf1jzCSMZBT6+uIQq1xGxQenjHvQyokClXSMIHoQG57ICcT
RlkgO2l6pBS/38k4DiWmthtBO2AOLBH9lKGX4OjN97H8PWjcXEFTCpbapv9fF7Jl/uWI4ofC/qEf
cwrkJK10n4NDG1UrSVQ86owynaaW25n14gatle8RinT1agPslUTU/eWscL5STEw17Kt6OrTmOQQs
bwc+PGxusG3Ln2i4HQ1DM3GozNOJktxR9vRBwiO6jjS9ZRFnEfdpjTg1x5eRaOj665QKNlQgJ010
47dFZIsm4xJFNjJJCa75oCQRz4hJwGbyex6NlVwmsNMm2BCwsBTwG9U022D/YMgtb8EEAPUkQKtp
1xRPb6AX5/PMbxwA8LNMVCGsW+wqLhZ5MJGw6uJ/OwTGYm5v4hL3Jihox/Lt3MIZAW/5dtwd2icQ
OuVXqYDQ2WcDKhiJMYkVQ9RtzeWeNbxqD2CBI2wZE09ZB5JgBMRUReKjb+2SWKdZu3UN80uX6MWs
bvUJJg0M2M7TRBt9YKfbzMZb9NR4+4keIKVdl+pDqGcS+GkFmVYgjrBfLTATmqWQnWfD1kKzznz+
IxjKeclBnNvwDyqp6lXMiyFdaI7rU4lR/vNyXLh7g+fWAem3VPF7lsy6oG0sZxRhoMW/ZxalJ0HB
fw4rad2wYtaWxn69vVW4SBAHuhJBLKu0g2zgw/vxHBRMv5b6I+UbIjLYzwzOIi8yKwgyPPXdwtcx
aFUDultp2SmVfA9mQri9+KPsS/PUgJi3/bovQfFM9Rv6s+uVM5oqYRNW2RZwAy+EzJhsyuh1BJ0i
dBtTDljoMhwa3VJOs/BGJ5QCaCDAwMtJVEacM6NQu4g2WxuZ3UolQ8wVjnnuWSJBbvD3FVkv4Tvb
XCj0AagVG18qjcxkzkEZktv1erOztS0PHv1VvCcViUqgtvTVIbTRyCkq0ZrVnQi/1qsiipQGJDhg
COq/7lhq7xeS1WfTkOMlLnNs0iQG2ScnS7pA6LvcZkEh0DYquxGY11jZBD91nWh8cQ6GXzHYOPwn
Mh7/VX9vNeBJi5JwabrSLQowVseMmiO6yF5kbTPkEiOonj6acZnf/VzM2ZiFqa0MG1Qj268ZIVdc
Hi8FrUaDsOFnDw9grgmy2Atuw6drvFfGbU9eL4nyqG84D5Q6ReLUmpLQsW3FEtHfe/RbnldcOyok
mi/Q6YYTpAglch1IzyTGYO7DDQE/D/BPSyIqiIbYwRmkpTdLVZLkvOdfbNJ9ou17G4t0b/RfB6L9
FDhA2g/73v1YocZjuy2esxrVt1XFFV1JOsnt0IxGDgjFcwQrmCVEEoRbtXExNMWHIK7dVtFrfDrZ
bpWu/rLtnFW+PfTjkZZrUtQWzMoCBvNvbK/cM+qKrAc8C7tPlvUzBcxg4AvqCvgggS4tYN+bFD/Q
lEDCk0HAwvKMONnOJFlS5g1Oe+lL1oyz/hUHfNhGehwizKrc5qE2nr551v9XjP82vP2w0MXLZoWS
VHCYg9ylnc0Qn+rSEJMz8RssZf6syuz6y1MhkzWTLWphUExDUYxiOsaVIXmpuZIAyOg5WPwpdHk8
ndIitASGO2pJCwP2BP4A2UysYNv8nyVhj96r2PvfX4vVQ/CQobScTC2jweKQKmAWzoj8k3e5QPxx
AwNO4uz60QmlSgzDUXrzd7KP9WuWm2jbctQsOvQDyOA1e8gQfULmLgFAptlgqAjDRE3t1mN6bKW6
GDzGfRQXsvIKKNzbOMiXBkmiRf97RxkTg4vuuRKQJiPK7Wl+yKSLQCFrER0PleSoloNSdlnl2sGp
kqzDBtKViHqO/s4jIkC8U5LSr0rmHOeaqrWFKBrbALz6/pQNU6POgOwekRu6+xMAHGEHSFdrfUVT
hezMKtdfn10GHhqQWvenAsCldANieFchhxM76K0v64sML5KJvTEBcllMmNq07Kj44V+OeMAJhSFZ
nCO/4BKQfLwt1aEh34Tt66Ia6CNl28oLKmI00hrAc/lYt/s1VaNaxstraYzXeJnP2JI95OtX3Dkp
3a4FFiskJo8DcWk3hfoyy4U1RQ/3/g8flTrmLnD8bDP8XoYl1xv4B1gjOqcqmbv31ewTmXdvvKQI
5OySpxvAaKBOzOdzeLnWivUUWBU82QhijODpFZGbeSETsB4VC3nsnTdRZl/OeYxhb/B0X+cZnmhu
CRrL3SAzLmn0D6PAeoK0jWf6V3DwIKRw9SBpm5klh91ULv0EWI5uTjO8JMw0c4WoiDpWpK246Mm8
0M+wzIk83tcJfBVz4GYmF5659FqCQgQhbSxdU4x33O0AlfTyN3VKEgns8Dudj7GMwLxYLOq052Vw
ftoIWrFqvrBxgHPyhr6jZbsymTsUrdfbkJjvN31dn6JQ+n2E4lwdgDXWIZdOtgIs4t3cRN8gyD8Y
7Gq49I93navylKrAbdyAPcD8VTHih4rHCJGZTQ3TTVUjNw5it/qkaGVIZhMrZxT57yL2kpbYzwXx
adjxKwpzs8f8aLvriYJh4SD7vzT3F/QGkoixRyhuE20j69KsR1aIJZN826tq1KiVPRnN1utKOoRd
Ph+5wAcjqlSZibLuXCJu6FJIdtyZTsULumvn0hUsM5yRk8OzP6Tuaox6wj1NiIBY6bH+bQqBG4QM
29HJhXyCEphOI5f6Sfl6YM5oQV4PMPFteLnQfT+NcdhVeXOw4aIVa4/vUQiAtXgGFR5uLeROJCen
Y2AFnmw3LveHxUnL+ZnlaGcBlUPGC2P+FHCDfx9KFpu1WZPgu5z982bixhM5fOifkz/GrZZFNix1
YzyVWrUsMSMrmcuR0FpvAnvON+8czh3UAsU7yTguTaAJ2ct1I8vQ6Tqu6OEQnKSDFDY1ro6MpCEd
QgoIDeJ76AzWxODx3BIvmqrS4IkPMmfvMZGxnxgRZH+N+qlIaIApDRM0jqDhE1i71dbOZsmVIR0t
zi52OavtrtbRoeIqENvT+BjWGhZrzn7Kx8OoW9wjv2fsS2x9tlOCi6FxBcOrvXsT7Yhl0m8MOwHI
JOb4VW9pAOLKNNqbJltKDTFGCPtgya0j9nRp2seFoI0opnt3jPU/BMMgC+Qn2djrnUdlEHIBSuwJ
0QUZr4zksZbi9PBfRobODWEQIRE5boBYjHLl80nqXWOyIyHUcUtRV1kJsYSe0g0ckeoqAzQfKMkC
NICecomWv4TK61kh8N83wkUDFRYyVOqwvNSpmUVYub+5RWuhHFpZnZON3mjS2vnfPR2spzy3Dhzx
0SLAvNPuZZQjr4panhM4zRMlJ+XruDtIvXWNQwkDyVNm6gsUoER78zUV/v+xzZyK6x7Srw5Bov81
uxKLSS8s7gXVTG/fFt/47paOIcWnLGREM3Nr1o0x20iFwcrRpjCfeF+Oy62Ojdflnuz7KgshA7i2
TPLlyJI+rp5TVvcMm6B2610cfQAmwvSb0baRO5iWvndRnB0pW6ws+thhbpoqYTzNNTTBC/3fy7JN
pXxw9Ukn08BXqqdVMj/3XXqbuulBQCiq4mbUhrmep10FZkM4Fg6oSphBooJZsWBry70VDDAh1V1o
9uMMjzUKnWcmeFIsPGNIR/k4fYQeCT+Da7DVCI/p8gwAJFE+y6iMx/5gx8ZlNH7yoqeBgYZoKnf+
ZDPXf0LnQ2X3tdehvdcruyhHXq4X9lD4n0+RVQUOqIM8B9DrISYxEDjcHLQw55ORVxHtjbgLkZxO
CkdefaiUu/5tdvNBAsIqXZhg1Fj0+ORJIzLHWUHtODSOzPMidZTfm2NTq8nTvyf+ZEGGyM78Lye4
20T7KrJ2tELYRiXFlCmGGfI7pHgwpndC4gh9FuNr52Qk9yXMaKhVGwNhxQNGc1oNYP1tXCwl49jZ
ntuw0NDCbWuXDLqLO6/gYpjLTC+a+yEfAQbA5X7+STl3gCeuU2/uv6L2pnUdRNWDoN8kHPjMAYMF
WbfnV4tayTSg2yKjOhCbEpDyTpSs39D60X6+6wGIBfLuqgOurXO2lpT8XBLZSVyggHklLdJ7kyQY
K7dEGyjWGyG5udkfHW2YgbJnJ2odCSNdRct1/j8cmllPKq8w3ucweMl00BU18I2Dn+e5EWb7IPbN
EWlSTnmjrKwFRlTOxRQNto1h9sJlVrYgvlNcxqWhBhxBe5+gp9Qnu1rAkhrU+IAW0aPrw+kkf0pO
s0PuXEFKEFI1+knj+Tev33l6iKQPeGjXjsLQkhebI8Rge2MnadauNqMI+LFToe7xgl1x1gDhVW4N
bvxIKb9EiSIvRKE+YUb205IDfN2bo6X3TvHUUjvC8R/jUOcM3U9W7jJVBSaaCAbiuiqgup5iHpQw
wARv+W8u5oqPjGd2X9u7guKPvZdC5ZjhqmYWgFyvBKI/kJqkY5A7rCjZTmEEPZu42Zh5UpWjE3x7
aytZaCTUEHqHXvhlgtw9sKk0yX/sJB8hwXh8pWGtz0zsfPefdECwX3UIBJTUlcAE5MGoMDRZP/PN
NoTJmL5X0ih4FJlK8icOCJ1gQX3v342cz50Y/cgr2ha3dfYjOsVa9ez88dIg0xKvZM7au2vdMmcl
GFBv6/4YIqME+f5ikCoBWs4NShZlIr77sZ7WzJOTt9x7viOXM6FfGoY1dqZGQY+BWykQHSGR/qGD
fauq7/2numWsWPOMVCDt3GEmG3aNRCsu5qhPZEuxgBjb412avoCCsaiD8VVeZS4HW2pxp6MRaOXB
rSdToryp1yOrTKKC11Iop2ZRIX7v/aDSj0zihd5xAWDuv6BT/9Hec5QsaTrhXp5NaJpZYESIhWEE
bKGOPlM+EZKtqJqsxsXq2BdyVxOu4+FktMuIZL0GnyUE6j2l3tCwHXWuZoHizs2p6AR38wQYLokT
079Gfda62mRYRT36xIx3xY39Zu9amXtpH90/7ayDusisOIIc/Kg2TmGBpRGkbPKm/UIBpJK+B7pA
U/M6izePntvbm2Tc5gibz5BugQ+nfYAJ/KFkUMIlSSfNG4Z338SR43abflFT02GGg7CRHQj/1cRf
XmtNjoZSzaL4FtJxc667yDE9Njy+L7iz7xZaBB2jyN9bJ+YAqICzGLWUHzuZodLv/Fx7SyAd49b+
4/izciCfarhlzUuBn3Uy8FZywharFXxGR0W6nDeZre+Uy8prqT0mOVWwjCEx0lguHCMJZPkVzbmC
h+nZ3txYmLsYu03bUPwEHaYc2zmuN22+QaQJftmzi6WcJZyPybHu2Kk+bTTyddpSdSIL2mj/Rb+R
S3o0+yp5SdtWH8o4TZOao8si0ctLqCeBybU33SjMQ06LNdQYjgLbh2zoAfXiHr9bdC8frtqwA69q
uaLI6ygycsDV6wNYaFR2bDBVV0Z+Z34jUnWAjKhGx7Y3GeM47HVgPUYKCQvnLBjQgRb0YHZbFq0R
bdG8joEPAATF3FmthLbGOYfhbIBJLgyvahWFgNSURppIaaNRuwTMkE6zPBcOM+l4t4Sc968HG65n
s04lafkinAxqS9jhtlc0sQnnd9OQ/0RwHopHH55hWY21P0p1fch2/fbu6AGJwQj4VtixpOk1rOD5
TJIM5VwiWCMhDbZPJiTnp98+5eHN/qaLzDJfo4WzAP+NBGJYzv8DDK+TprozYmA5p8ykJ9E+OMsc
R+w1zzLkBcdYOzsMnHPTb8TgkigkCVcJvhgUCOQEalpu+lPgTefT+8cuG1HXnYefs0KBHJG+NC9W
o37DeAizeyx2N3DPP3J1iuyTc0jhGnZ9pEl48jSRiV8Mqq8zwLBVP5llWXYNWaQHQOsOWRTXMOLb
uAEuyffaUyIRuCfk/nQvU3h/i+cR8EyRtdmDdMp2DqefJ8aUQZtPLqCxn/JPvRgYcSe+DmOneAmO
pUa+GeRlaIUhdC8I2bAaawl1SsE/1TAICIPk3Yp04YIP6Yxq1PekaITGb5GkH50aGM7mvlGl+QkS
CA7+oQVdQVoJWto+Jv92m5jWAgeaI0QIWCFskcB4m16sK3l0riOFFRVO3HY12SfL72UhTQQT1BQ+
gGHWel9uKFBM+Fijr749K1P8XCiFNyjiO37iLaSC978KjUu/AWqVncgjegCJ6nld1247xSuIIIny
g2QiCYpWJF7ubI2RPYiZAa0bN2rFZyY8QJV02S06/kHGmAwDEQivxqn/BKvNvtIDEgPGmS5SBDIN
j+gl3L9yP3kga1U0UJHGFvRNWIYtTC7d2y5h687BNoc1ucUZeiIJO20QLI79fjeHHC/RImU/NBNv
PcafcfLhMy5nLztQzeAFCkkUuM2D2yGL8r8Pjd+waj2x657xUM8n7xCqIhIIIt+l3lGH1gDmQMPc
nqCcvNJJhQpqEOWGjxvPcvP73MiI0C0PXC+VyrEl0q+kMJ6x8mlJIF0ceX1PrceZsHaksAdPP1+q
scZRET0vRNnQVDWVLDcHpSaEWIdSgQDyPm5XszGRY3C7zl5x5hiomy6YM2PO7RhbmVPW7J1R57tj
sbcm5YBnUq/cTKCtL/TOeQSFOpvuSL2LpZ3RWPSCP70RvJHznuwLiXA16p95dFew524UyCrb7IEZ
XyTxFGRvahRvPrTWuGq46SvgTv5aDqTDUF2+OQr3FUvFIPQT+ETQF7dvZO2gyZeOH0mDRH6vvc0d
jwH6QW5Lpfg0AV3AN8vOiDVESrirV2YjNVBr4LAL4q/y6ANAH4G/WS1N6f3uukhn8GCsVpu9QFIt
fYDUyUedDsq2xkVjEuH2M7Um2hlRzDGvAa3XSVuGWRqOFbEg+fp/MtOaoelOiocVYy8DwbzS2B2G
v+PLIjIcU+YDh+DTSE2bJkijkhwM1VaDfiVX1geW1ggKpjWk1BBu1t2saO03capO9QlfS5U9zW/E
nY3KzYqayo5gcPutKEW66uFHi9EnpoMZ6VV12m7O81dwFPfWid0DFB8pMSD4Nqrt4MM+CE81lBNP
jVM4UV7u4FYMQ4P92YigUbiPidN34f+/JhzkxKkpbGzcvhf5X93Jw4dH8a7ZTr52qGPx5Onjor7H
/gfBC5xH1XAWp8GTT55s5eiZvrVEWpPhyHOd8yH04oXzH9qDM/q+6HUlbJ4Rc14Cp/jG/dKurEBi
LFtB9hZUchm/Zx9naS7j370Jcxl1gYik8Jv8XLQJsodGa4SIOCCkwgNu9WbNgPHMO16IyBUcdMrx
EdGUocCVMoXG3iYyxD6DLu6ZLZ2WdNl0sdljnRKInk+4tLYZD6kzVgi6grxFdGA8BlBkauF9fkzn
CLgCidX6xnYwxNDScMb2x7sFBppFQ34eqYZIVCOH4IwuC4yNmum/lA7j2Iqb4zz/7A0QX/2UOkEt
A7lJp3wEb1wBI9eIQTHbBi79LOn8TGH3jMw2lPuG4VUdLrwovlklPaO1pyiiftVyKo+Bpnrksyy3
FO5hQkSULgu9oM3vs0049Hf3KI7+f5QmxZNFXfmtfdo9Cjt1iQLl2lLErfKWRbq+cGbb36Nfjc+8
p4v1KtFlsdccBC2tywOK6P5ZoMTNcpEVK1LV1AEpSmevnpdrz7pkTthtoQNEskjFlOxfQWz984uN
O1k55KSMKMYzVaWX2ZVYVX1hwQgnRsuFhzolIzsd3EljTahhKFZugZ2lycCpC+bDCYkiPao50Moz
KOHmPOBRZenN/4K8WyYgLu1S+kp99iiqPtQpB38OpnaJVWlqLQzfXff2uAh+lJrCfdO7tJpN/6HS
8AZqmh4O5CHU/CbApGi9Th+4XxMD89moLQhnviCu4kwmWddrU3uC4hA/YgjwnGWBpjL6K1GwxYyJ
IhvUf8kEl8di0qI+pqOM87raeJ/EjS/xVo79C9PNjdusB50tAVR2837qW844WZb7rZOAuiEzURMz
++L126x587pobFRhLHcPer8DCkz9Hq9Opv0ihdwfX3YGBWjjuqPtJ/zh65PICVd5igdZlvoIR2/J
qmy6KyqUwdYG+DvLDzgkhOv6g5lnHWCA4ZmRkyOp6GhOZLFKyoSRApWxS6JqsCaH0FctNw5SC2PZ
79B04wS7NVaLChf3q7171b5oo99mTkMnq0/piAejF7ur1tK5atef390zK2nQ71jkYSQkcXsCAAPw
6lyHBAvBfBDgyp68mRluQYY93QTDuZjyps6Grn0eCKCuR/pr3Ydh383oZQEUlip1ljToetbnOK80
PqagaMtUk2brIZ5yL1NLxr1KrCKpf8sUcGDcsmD4DhdEqO0Umad5if7MaeDlQ/+Z4agcrDVdAT6I
/PU/Ezq0LSRJVmUqg72NnBeAgOI1zsBwknr/mjnkRUYKlJMNVcKC5iQR2I0KR15egkrdj5A8Kzvh
gApLVS6gOa9oZDT3TP6JU0mVbFhOpzDV06LIr5OahlcxXFseX1QEA4fWL89zkJ4x5aPpaazmZ6Ui
/AdReVldjhAWJejMqb0iYr+81JKLVzUGEJFlSaTfVL6ftacRsCEeXQ2TyM4U1QJ9pQjFJn3QRHrj
4hgH5EXv+jyV70C8+TVYCLC/cI4xS6k9JOjGBp1T6VbG2pUZFBWHhFGZgW7jrYxyIqPXXQ7zblM4
vwtCFNcyxYZXH4E6V18c7FaDfaKLF7ER//0LIGWukp8m1km3Q8Moo5amYuDrNFZfHnKsIImZWaXH
C+YczDOAlrSFohrg2yU5vEy+h4cTaTvelGNKQbiYgZdf7CbRutGBTIMDSuxuU8fpni6W56xXg+6p
RLLwnXPBckft5zMJSo/pU3j2TDRSLS6l18orYEinD50q6ABhXgymwirqS+ngCphOMibZAHHJo0rf
MWMpK67BwRDf+3iYu0xwguNsdKq4xWRbN8fWhH/WhoESf82QVw3OJtDVP44DpMwVzOkJTEksyUqp
X4PvL1E0mLVblAAMo9G1cUP6y78AlQT9iiTjqP7fZmCxf6o/zdsN38EaCQcSMweZWdku22TQvy8G
XdQNuZYeHHjINBHeRThXTw6Em23SPeLtRRlsT7QFDrPn/YKYmEcRiNpcf4BscUBgTxV5I747xW5g
lhBchGiV5DMQSNIJdICCxKlAPBELpNivhp+K1Dy9EhO72QT9aSAq+lojOVbX3rZsYnU2F+zHe8NS
ghg0SFLVfFkK9PHiztzjvMbeaQnOI+E/r+KhRanTVcHOVKUJ6nZL4Xl8vOSCKp1bgNh5D4d7Bcdt
T3Elj1qYmVklHQumHyBAlC1EGAXbjIfh2yrb1U5pzT43pvqdBBMr91pxkt3FFssZr3pfMSaoZ6aw
UbwbPVz35P5pAG/Av7h/RkIGBSnQlhsd7KGLW8iSuoYsiLGIjKMJb2OeM3nPdHYKrlpDnvHNwijT
3ZTIE6F4xTd7/WljknEv2De9XUu5YVsJWbRR80d883XC35iW37r1oISa2sNYwuwpsUINgfoBmF61
KZuboG7dfJciDCTbyYUyu5oexx3nZ/gOE0NFK7tKoPqfiRbubXiwrSALLGrZusv7I+Y1gArY05Ng
2RU5+Bg+tHHWLoB4pdj0uMLltgok3b3NIdl9L2DIo9LDNZM00gnmapwlzdo3pIYi9GThxifHBhVt
pq0m3/leap4ld5SNy16wXrdm0ooM9HScaVtANZKg4QQqtvDM+yfkGiXv3LTFqdxWCqC293paBtKM
z5Tipxg40wTYLSQQBPt/09Fy0lzJG9jFOJiF5ZI8tvWj5G4hL3XlZbFE92bqSpX1MYMjGV9Wf/IS
RXIUVlsBERd7XfH06ZhAQrzlQl4NOKMVke8DBEKlDnl+5yQ3/iQmc59BNiDIDADPJiIf4sLiz7Ao
m2+4VUmTja1tJOjFxbLI/5cQcDpwXeSXBM23d9blwkVd4FEC2o2iFMMfdBRycHqsMJd8ntrb35Y1
kIlja0cp8uAPrQvakBxKoDuSFekvppHEbqnnYOeB/gITTv9shc8zhNnlphGGar3D/Y8Q4jQG+pVG
urY3C5h73gEHxTqNdixY1+B95D+WexBiUCk5DmBdZDJePoFkQtc8PjwwM0+O5IGgVMqbCUyQ9jzZ
49e3UdX73Li3LD2/OqDGkPlg5ZIPnkSlzcGlCNn5pfYEVNRn7cAHHnT4X+MEOHvm/KrgE0ZUDkq5
X9K/exkfkmkCz4noAkiRKSh2d1dsiEdVoEDzYYWcNzLRMbGtkd/5fN7bWIT4MFGIQFX6F08rdrHA
KDI4KC7nAohbac59gbeZK7vhLsYm8+oQPevbhoKBioowbB1Pi1p+47J15R6ZDdihvTK1RjRrZbcv
aKMHjACJYLGy43KivhnqPAWOw3MksVVQMfR9v20TGBqngUL8v+XUSmrg/amW2PZLIUG36yM49JSF
YJh/DeeE1ogv0/0dwx+KvJmT/N8z4nBLpENbe82eBmnobaR4jWpfns0b9IGZRUyvEhsUmasV/E3c
1jzdp8LtCdxzL0ZtOI8Xx+LocOJxidEsOjpsS+ZkMLGA1GPmqnd+cDZqLkCFhgZRLeQjlQbJIfTD
QQrfofjuyYQP1lFwPNbySQHB34sQIfbKo98vKJKjUzFc0srWuGzP9r+i/ImNfz3AhFmSF5CuL8/0
u1qIS+ozFDj3XfUp6YNVfH+T/9ln3kANV3ugrOgDHlAD/N/LAHkk/6nox6tscMVrpzl824Y64tAW
p+vldSgpMxbEupL0bBwmx2yBoMBA2ZSJol4pkjkcyC3z4Cd5NK7pkdxN44b7LNzl3l/b3tDHrJWo
09LE2eHG/PXvj3RO2WWlSA6TWxx8lB/wuG+S6sSoSrVcx0tcw0CKGOjtjTJoLLtzaS020w8OKIkc
mvO083SsNxfgcMlaZFRZJABMVt/EwYoa8/lZaaEWwTBcNDFQpdwvxdfoVnsM6zXZPmdhSq7USPf7
8QhRweMx7f21qI+/LmsUQFk+dhKzcBjiSohMXPlH4l3Il7b1riqIRQfmV38LJja1T42q0VKwG2Ii
4mo8p8UaO0aWjcdami+KWqNdEUQ2AkY+dhRFQv13qZmlBmN8FILtmGuait3gzkL+oBD1YdbwaHNZ
kBiiQ9OsOuiJ/AkT2vx05ucvFl96czS7AIgAQS+JRyPIWGCaNWCnfIBHJu0XlQnAVFqpE9A5jNq/
xgaaMY3U2D8jB1bhwhqTmSLuOLQUITZx481cQqaWgJDH35xLSzUU1Lo4vrOladkMBZeV7mCjtd4t
rywmzJarxh/01uYavnkE6TxEzX08uZj4kp3lbvq9uLbDl2p6837KcdZqaF67hOKuEpoGaJVWkTa7
UCQwYHarWEF67/nef0g8c9FxUvbus499XoqibIQi2IlsECBrnJmcq1kHgCrvMcAMQMYvR+n2QxTS
2GQE6g+PoU8RTri1uo28qYWmgcGaIXxgzAFODwbLe+4vN+6Ojy1EkTcaVN1O3Li87C1P/EGu2tQ3
L/YYbD6xvUruapvteQso0O/KcR5QrV8BPQTjfrZRKsQ+gSawMgCVzBCPFzi8YiSDGe83FxpKWclB
/dcKmnYHieYc2M4vSCYk1vyB8uDJgq9uYb0SmNTL+kv2RLQvPSxVSyj4TG7u2kxhjz39Yn97AxU7
2IkffjI+v9UJFLuywXI4qH3gANwxjrwPLl9+ZL/rjF1jkC8BO3oRzMVTay6nhrfGlTh/CGHnTBW6
fXVexQFtzjRGl/0pvSszto/8QCJ1ICE19plXXuvHhnS9Ezi5hr607nGNXDz2aT6w1bEHqjk7PU7d
40XDqeQrSnjC20XTAWJNCOJvMsuZEyOniMCyJIc8JC7TFyBRIoMYMYSl5f8Jxmsw4jANFPk+PEk0
AlMQmP0ipJ+TcOH874H1k28lMw+v3QrmHfPfJ2gBaixEFZbprC7d7MUIbBXcaJLqM+3OxMHWC69R
bWmPgcUm/eS28p8ofX6Q7losH0jErgUxQND4OPW4jED5Lz2Re1djzTsbmUoIVQLLBArDjhnBakZZ
8f/B+ZsCF7JvZ5lNIK9AR8znptCMyAFxQfOBlW9mnNvxsVID8Qo8s2LokJnOUK0u/XGJqmBMr4T7
5OBs4nP/9s1R2azOMx5TXo/ud4PgdaXNg/lsXNjA0TJ4mjiTI/nv7iEUJ5CrCglw6iW7cM4gngYS
jMpmG20kCw8VVB9mOPXRDSbAfGa1lE2+9/ntwcYsZUfV2EQpha3N7osYP84JJ20uKI++d8V4pJkr
gm44+V00nFGEmaKnrG4MnciqNnqpItbVfoXF4ztsGWzXU7jB+AT/vnt3M/Tlce16ZQjanAkEL6ol
QUThmRUbal9Y+tykX8K7SuJJSiOPBk41ywDGWZK9wQNmbv+7bZba5zfaBV/YrTflhqIFLCuO53oE
+OSK6e+LiZav1djZHCAzoHDk1J9NhbEZ1ZOl7XdU8IJ/Oywg/j+UVGJIR40o4EXue91zUC8qiqVb
sofxs8huc0hSeX26jfe040fwSCvgquL4IwpdXHFc5xZ2XZKwzBZ7Ngn1MzNaapSpxJ1if0x0IVj2
QcluaqY0azhxQ3FaSfGSEmUtKXhbbpWGW7Z3qYUrNBYpeYQmXZM2y99lzR9eNrN+YYkWk+7XO5Hh
viKO6gfPy04FOmjghHAfLXLikmsFwAYeKY5IuHgxOBWxWIUBFKgrDqxHtCO/Y9vBaRAps+HSIXNJ
Ztp1sIjEx4wvgr8CBlQFpLLNP6M+6vXizuHh3mTroQQXEP8qtw6j3W80rqvtNZ9Z98G6P1O/+Ruz
JsvZ5llCp2h7KXL9a02vMBbZnFC25jUwLS2Jv383WPVmp490KvddbJaJ2eEzpb90DijVhuh2Jm8V
cgpqjU3VpjK5hFyaJUVspdQlCjBmmPcK3F+SFozEnQgk0bceK5Zq7Te13H4PaLsFlaeM9BOaAj2I
gTDDBH9TngB32kMLeOdwoz3XrLti2WtxAgYzJ3C4PFMn0Uu1iUXvDbOHF7n0AFkexDnaxvxcGsYy
1tmFJ9ZJ7E0anIzZgB0EUAMyNQcgGXqeNd/PucDWlwf5fQsQk+EQcidyy1+NAHeSoVcj297DCRba
DE1ApyRGNeLszOpoMQ0Neikls1qD3Mh10gt+sOXOsLQxbP7If9mwe8cHUe3PNRBSOzRpEUdBrRIb
U7/kfVIGNyCaXNIpHMtzsc2YX4+5PMHGDAYr1HdIRAq7y3lW+osPh7R7W2RJu0rRVPU7pEDcLWe/
P3pvXnhI8cOxlJDWjWSMkFHjHQ+wddJtTc1LIgOgh1fBPPOL0/UYefMoMe2XgXrYJDpsZcVHkBVo
kQs7GCluaMzhzo2vWQKrdVajmsPndrKs6cuZrxSragz9ANSJl5BETLlH8+PkzDLjt3t/9dMQ635U
IEiLxXXifUJsr9yX4XH+KmEajJpYhgG7RIRrdWcSS17dNHAtHUo/GeSN1lWbsBXyRqBhktUOiQck
3YPqiSayX0BgA6tLc18g9/Poe71ae04yfr5fVOfc2usHnR84F75iJUcWKMdF5w530yRTiKOLVUU3
XgChPwnOgh8XHlIBJQrSjFauV+esRu4542JNq/UeVLcT4zo62iunK4FsXPHEZ1s+3dl/BCF6/OLt
WmB8PhWgubGc5wM2pWBXee2HDKVC77LJDPVS1CGggM8ViXH/n+8i1cPhx0Fgan6sY5/xd7H1XtMD
Z61D79heLDE95O+nIPiKsMpdT+3v+rCf55C/CTT6FjUCecMtYSwMDJg6VO0KoO+2RnXhW1Jnnm8I
73gT5vr8DvlGSvItV7nJybaWQUK4kUs7ZkyX7D9tWAML+hORmLcT7E+pDUTfCXDyCzprd+LL/5TQ
a3ZzlVYSAxULY2JqgeF1uRYzrhDQfrm2sbH1DGH1mOjhh/p1Z7+FvMMmh98IQJcc5oD/uOq11Ri5
sCArZj5isI9ujOGI01DwmsUQPEsnfWm6APYZCjRI9K+dGMmg2bHb1fK5ZG+lM3Qae936mIyyb5H5
GTuuniEpD9D4nXXR1kew4lMV8vO5ce8jduYoFX9kne/iMb6Mog1R0rZdemU7WFGrFqJod5wZP8r2
3eHla4ljNVdZFa1htqlScEg5TgOtJfNPW+8cTRJ0R9NuoJT6kzXz+muYko4FUYN6/4C8sOuVAYDt
yaLeAVSjobP1ZaHuMsXRo3XIBPIok8uaNbVgf9zeVC+iaEeftqlx3pADOB9vQNkJ19FdTn1lZzPh
ey6VJFCPbqC7mne4T6/HPY0pJpXNGWbS6BKVMvso19LOYQNg4mkAWFwcVbJBrSS3WiGbKGAnoWji
I/U4EyNM2bAE2GNdthX2J8zZoDZuJSlONrJ14JdM8YL6VQLgGPTyleEESGmJzb/4xmLmK73iw24b
b2zfFrF8L9bheWGGP2d4sJ99llkJ9upQshuYiwEokSLF/js2PL0ABTX1YJcHtSzFkBegV+QmDnTw
61b/UVVtjbjPE6nhngIvF5ArvHCKnasVqgzSMqOj+LbHSzJM8haIxDJtsBlVdzQQUfrz3CkKDbWB
tqBh2H8osQLH7Y6IGUdBa4TZdUl55yN6Kz1h0Dkn8qa5qubknn0zSNjVvsxvSffgv47sP94HAsLe
2FVKBajdrE/qObkPCQb/VZ2Lefhpb/lgUlvkJvVz2o3VRRbE2e4pKUONz6yI6AKNItYieAsPH9ee
rbHtSZ4GAv3WOdo4LcxwrduBztzh5mz9IHqF8otcDw2txvDOxmPFuXtlZdEgPf4CAbR1eT4KAShL
bn/8e7pKk0ehXG3omBG4wyR2E0s8TvRNVuRL+A4RJmIEElaDoWnSDmpY3kRLTHu3eAPqKHZCEIJq
MJ8vZLn/fHuqUrLxEAHXLmnB4W4NMjRLDKxuWcvefepom7dXFAu+R7NP4pCp4sGt373ipPK82bWm
Mwf4chABP7EhJuOZH+ewyyyGuFYqOrc1rZupMFHOShvpoHIme4MUmu1Pf98/aikSEFqRDB48ojp6
u1sWivEpTXdYW9UNN3OnPEWquB3fhm20i68kO1btBekDx+vXe0mPxblUeSPP6s3P1vCvwcYf8FO/
IGNwbjRhfqEAwWMgBYuGJvRv0KiRRy1+q4qlIlssVxhNrGKrLYe6C+iGoxcekISITV2OhZ/s9Is1
KwbobVIyIjsB+KRjfV0Q/fusW5VP9+Rgnvrr62eQ0BMcPOj3D+DdwE/CneBQQjugghlow4gqJLrD
mr0Iuty3vJLey+P2ELSEoVM2+LKDalUAJA3dy7BZne7ud4RPRzACn1B5lxqBo7SviA9NOjbc51i2
7rUFwzgxqeOk1+BnzoicfO461qcFt/HF7JOA3nI1OVVh7wx1vW0o1W/pwVceArnsqXUAfzKKOcCp
JNtFGrri1He2xHOF0tW0gyW4BrqQKijTHXCvjPE99zglyfyjFLM2MEyOVisUFexcP0H19s2vFZse
oUcililk0lleKv5WzK7ja5eksZ9XO8Q9sSZpqmBgqM/nPDRaXWX1mZRFLa9gRsoreSdWqmZkq2mc
+mzNDO/pLaA+1NA3D9YmibKxRd/OL6f2trBCLFoB/tcAT6XSPBHm9wKyi1sMwYXHsMtEgwDK4ZTm
f/hijcMilyclcQEObhC31y9LQgG/HZ5HK+qoQaBsAvrIeP0YGZgwrJKPOyE7FBnpFd2buMD9Fe7E
dt7V/bXK02lwR9EDnLuw1lXhzMJGQoYPlNfJ1mlj35EtXWaNJ3lKHhcZ+zQCHsF2JWHNcCtTBK06
XeIg+cwdwS6ITWl/0Ca/0cKfAohCCU4yE+Rt+6wfh8GhAvPmm8+6uwlvfGKQAB9ZtUyUfsE5M4NM
DdhP16jk055hmzKAO1KpJnKKkiwkaVqlVI1y3qyIx3NsUvlpYqo2NcXHMC9CSoifnzVRdXvp1p0H
LRx6yY5zOJua7fjhblLQw3KYO8haJ5CWyZFqdVxrh+seTQCdh5G73mqN4xfPOb/TrrqiW/U5mPxX
Z6anxqarIOw5NFmzex/0m9rAq0XBK3YGadWKwXDXmH5e+RXmmij96GJXBBBOx7vh3diTLy9iMgae
zrSuxf8MPcWMMgGKx0m1snjDPKxDa9G55aT6VmuV4BmXaRIheuYt0/LrrcCjBbCG354tuE6pyG49
gLhWLR/TOO7CzIMEMZCxuvHZAE+1dEgn9ygkMf8Ikgye5H8GPCt2SLoP72XtBcEPPcL0aD1cSRSn
9Y/FV6yaJOAA6oIYcQ+qbalGihXp7zNNSUZEm1bTGVYyE999W8AO6MHaZ6Wbqf4y8Ke/+KoEsvfo
Komii2fcgywOvY4Q6OXjJ/l+dVdIrM3WTJ/4htm7yjIiA5l9+tKgSEZflMo9p8HkYHGunRxxKM+O
sk35CRTiPvLJBOC5HVS6OQDFbFEmymTKEYprcnzlzn8d+vj8X60cAM28EFXVvOjG0E9LZEdyAicA
OGU6IkJcqfMQyHYCmLO+8rbqD3xpY9CpuUz3WfqiFKdcqYWhqZlQe2dhV/SS0uXLV6lZ71X9xG9Q
zokdHXILiWx523GyQnQGVbNMJn/5XZq8d0KjCCghucLdqnSv/IdSgAMeeqWnWULk07KZVH/GYjBR
73E1id44gBv6f2dI93yp7W+M2UHp5DsJMjXiFE2ReueL38PhVo4IqsT2Ni7qIZbYkAhYufUeJwgn
8TWX49rc9tAsIT2Xy0aVZnwifmG01xUivEP/QdYMKX9jR7dmmYarMiVn0nTIjHUMD03/xkAYTBlf
6X3jdRQzm1Bdb5sUod3YEbNQGR+lL3mephCIfv8GCzVcYc9JVg9Mk4uzn2c8scDuD3jy4MC2Xxgs
P9BngsBkgdqdoMsQ7gMPeP6WM8tNoNMCoDXDuArP+fBGjLdpXvKLaUQNDYYxwXPajh5f0G66or/D
Bx22E39ACuWO24NxhSGw6UO6qBkQN6gr7mHmukfGu8d09gg7XAqujoPg+/K55Yl81RudaC8ZO7Aq
kbS94YNo8BuZbdvhmo3YcL/a2uQd/84Y2HWlaVgG5HAyCO3RsmqpWAH/2UyyT3VFArP/FLdkBoZg
QXkD9rTuN7HnTmKAxW4AJILmOQMI7dksCgx7ygam+g5gSFSOGk8s2jeGhfFpTeso59KPm+ej7fnS
RB73uHmUWLQmFFQ0OzMOj2JlmbuU+tcaWu/iFWv3HzLqzxDThNFHTHzHbE4IjDlte9ylcmZJtIuf
P9yaOTpatkuKgFAKTdpFf/TXmN6+eVDtgJMSaLbTVTK/enaSF7j5DbUxaADSAfZDP8x62O7QydB7
BjUmz032d43dHq1hVt0Hz4n+CTi7bGabxS61ckh6/8G0mGwW42iZwS2jX3Vxmp+VP4V4bLXMv2rA
tAChxtGQifj3Evvdjg5ZpzCpti3djX3byGarjkD0m7QU1c4Q3cNGTgXTgSK699tZ4IIoDyasMpGD
QSa2MKw3W6nR+sLLFaTkFVObuwEANqKjj0kuX58QRg8YKsINwjq/oWAQdk+NQN3t719DeE5Zj3sg
IvcLsUmhI5FovbVyj69n0Auv0IHhnbFMBjHZ82WukxhqKT8KFnQzU9s9KeaQ/4igYe4BYp7saPbQ
KVH0/ue7QfuNdC1UDDAhpx8H6x64HPI3hStOptJZ1FSAQrI9z7c6Pa7Ny4rBPQz8PoSWNsdeCZ9s
W3HkbkYF8uvfBD3PVCC+P4cnIv+JtRV34NOSyy+4hQ93+rpPTeSmuhggoFKxWZez0pR513Asw6XY
/gIMt9pzXURvGca6Sb0OyZEW3TvpFS5z5rTnFrBxvWjS6bTjYdbyfECyUGBBh8DM8ZhwCMUgX0Ea
bNZDKMubPorZkMAhisXw8qoOosnMZfODxwUQz7e71zn8gzsihanSVS5nAlum/t2BEK6+qvqhdmJ7
WrH8yRTStioEi6dH9iEJR9TIf5LbYugsU88w/mCZKf54EeJhdman9OZ+14qojAq9v2CAC9uDKKVM
jit7xTaGYP/K0z2w2qWNsQVACMtiacrBLS1yZnN9VmHAUO0OnhjgliyB6HBYQc3D6Ub0q1cpDvef
aG5gBa34hj668yqMECdVxLZihC+3RyQ2vC8E8V0q7tgNjwf5VANTJZXlO72rg2tPi00Lp+AaaK+v
IyRAY+MDpjrhBGwO8A7KkYVhB2XwSGQAp91lQWtT9oGlCbc0XVeFZuAxwG3wZsakii+gTk2djLbE
k6u7fr1piSPIIn3QZ0BD196NBA+2zSZSmwwnk2fg6h03SZvgvbevI/rVooY6tPg8vzjvUhSUw508
mLNK5shSDmsqg3YKtwCqiOkpzJPajog6I9Ai5HlI6HdOGQW8EudolWMamf5PEyu4Fuk5vh4E7d6p
BdkoWNk+9YsITvf9n2KEZ8tgqnAwwF9ZIK0KIP5JuEHmVPTe/3VVZTqct85BOF2d+FDjZM5MdmTx
+PDGJvrYVDJwQs4bKZFc11im7zuyM54kuxevSL7AvrmUNSHe2qIgeWmEfvvurn9UZ7LB+DKPQh4d
/M8VMvfYox4PUAVOgMrLvduhs7KVfcpGn2G629LMsakbGqwpLX890mizNjA+G2I1FUe/u0Sxpcee
7GJPIRoWVH4IEMcOMHXZC4YBs1LaWPVXVRT9hhK8ItENtBGDcI/sV+GVqJiPB4cgHTXmky8sTYAS
Z1Z5bor0ucbq+DJ9E1YIXbjf6ouJVLAGKu7mLO4QPTQn6skroAY/ME27/tUExn1YcFG+KeLI8qEB
BKcVnENTblBlzZ4JaPAksZ5dkYqaYKF7/t5Mu6d9oXweexT+Oc1S7cuO7UbQzq9c6rgSaLmZJ/V8
toYfToXuXTmGn/cxqfgsGACdltvWSbk/ty6GwYYTRDvEQGxenwgQyA39D/g5kQToQIwyIUzXCIqH
+XIJHTuBxt8E8Plo7+bvP5lOErNIahAzL9vOGA+ui2yOvLfVTElBfa3UIT/yPFrC1XW8PcVdRILQ
GeBGVWwou/ei/Rk1rTCZW12o/dpbqx8Frt8s1qAac60nI/K1zCFGTbKZud7TJeHdur2cvNR27xLX
8I2ay1skPVzZxTa4Ipa3QltoV6mdVVwpdYxObjaABOwZib2MB2Mwa27UIyr23Z5ZZQTWbnnPZmBg
9a4JXuPWUYqPM+9S38IvRqCSZU+jE/Sq99UQj7SwmS1uc6PYG6c+yY7+GR/FuDW/J8mR2H3uEqOM
ixwKxb5rhshIUzVQD1DQz3XFixQ0FHGd60TOoTjGSl5I1lL66YpaDKg0286rMsqQurb8CetLDLDG
ntuwsvkMwdNCOUkditFqTifZz3kQLZ7kam3+p+RoYColgo4+qhc2nOB+/8wPafo5Gq21sUZQY3h7
rpwKTK+JDWED3Yk4BMAHFP5XX1/Yh/KpHnKAsNWEcbaoars1wC89Og4/KTYP7DuJ4vO1xTAHSxKN
xup0wU1OzSmfeqHIwsm3qCZrNVGEEm/buWJOGMeuI7I0fud54TkBbXpha94Jhn4CNoiHzYBEANyN
qDLLGEmLTd5rCTBDgufQ4AZoa/nLfalHWtvfUDhRcNaGGkDuX+5MIPpS/mXyHy7uD8g681vdPYgg
/sIqVf8A9XrkgjJC/zHhMGey0PnNPoSvgSTtuOtpxTqPsSmo/vh9fCIUokcEdgmpNhrh/6HfWgLE
XaWXhq1cEAu/ZQRVUeADK7p8VhdNEmoL083r9IhbPmzdpyXWkqDrvZd6GTQHXEp6MJu1kxmpjI20
pyEzLyc8PrbaGJshpWlKVVqOu1DCe3dsfWHtiLWuFgkrD+kSfJOr/TObB0Ahz+R4Geu5Ox8MnSUj
R3TYDzbQXX5ImCi2+PYHkah0UkcwFA3GBQPRkff60qdDAe9RPXiRjdbSzrcDtZUc+nhWTJfhmrRG
f4GpLMKV+mIfm5aKlf+uB92j9Te8w9I9d+7VlsYEyyUH85/O7dsMh8ZH1xpHWHMSqjpRztiOo6v4
Zh8wP3BuOCMYvZyrRRMahUSglmRy0XOMPCXwWkfyAtRmxaZYyEpIZHwIwzyu08hQtwZ5A0sT4ils
/H3S5RZ7lLoKfADJRGXditaagpRr+uZzhbf4A9dDV+EnT2lETh6b3YjFNhWmS/dDIoJyyYlQDBUG
W5ZtONTl3KYUd4S4ULjEjB6ZsV2hw/aG+bjOB49GDJeXO6i+GXXJkikLeaIKrzUntr6E9DtF4jb3
kGMocqZWrU+TRArnqsh+moLrRzKgqbB090wDKaACGeVsW5seJbW8ciY0Nt2g5+b7XDNIqr78M+OE
XR2QzAd6fZDO7fsNRI2YpDs409wYV/im6JeYu2sr+R1lkP/DBPA48n8TXvyrYatajaQUjyRJjawr
2DjF4B2mGX6OW5/v7Mb89D8ec9Zb1tS+QKaIcZ/tNazKK1Jcfg//bAWtmX/1mGvyAqpLQO2DR66X
SqVxvGrszsTio3yPDKacqtmeENll8tcwiyiZI5kk4kvWg7EPU+SxnllGhC93e31ohIr9V5+scS/H
ret1GdDsw4yD06zeZ5dfstZYMzhfqn+TtHtRSNmEuy/PqMKlOGINGqcJ+UZbt1wc5ZYBH6Cd2FWF
IfJ81LCu2V1KHnj6xjYxBJqq+HQbcPCKPNU7ElljyV1dnaHUrZBD/WPqEWa1uMdOlaOk0IqNea44
WkaM2uaShnOGmSNTWUycuZ8vNrKKX1zt1tZ4RIgD816qDowNUGlFk3obD9KFHmtOxmXOfaBepQ9F
hcsWuk+ovaK4HOVwMrUQR/st4TcU9MR8pdPMIeJGoe4QUjjcZpJYy1Dfavugx9ZHvswLQ6wrvtPU
6ZW7Ow6PUph02+LwYzzemztjjbxxlJtdOmsd/GcfLWOgyYGNwExFvRVhrVlhtSqaULEDfmqNcw7m
9rMKEo2jiet8MIE0/rDHJ7IhSHJ9nu+zhCIMR/dy8CWIdClDa3DNxsn+frJYKjzsPnuVY8iv/EFQ
MxlUA54kyRVAffJhOd2HdbrAes9Bu4ZU8TaDZ7raxNhgdBeyuKqEzIZZrf/dHG+TSNx273vNnFGq
jhmv3g5418qVfpH/EHB4rsHFUl2M8mnNUSO5aqQdF43UxZcf3mzIMEnpSQm7uZlDCz6AGt0hOpou
FG7qEV1tmy3f0kzilz8terPZ+3VZzlkqhbaGblEail1T2CQSl/SHcPSgv3TYh6zjDxZtFA8Z5ZyA
+/MT7aWAoMN86u3drSDHDWRjwnnbwDCP8ptKP6IEhevVQPPsl150LAjA2FdgpF29zY7PXPZw/1js
CEL/UN8a3C17koqxraFSZ+wxTMZi1m1kSxkdmAVJWIj2CISrVZvZ3s6Ys3uTI1DjH0XT7XN7El95
DgUJT+9wQaqcCnCjb8PWFrw7knnJ26oLfsSlz8A8IVaLarlk1A9X7ZaskTeww98HIMfkOX1ETW+F
nHwCJ8aEx0WXczag1m0r/GJwk5kmrNS4+RgBC3OcenMPXVzlgnrPkh5Uu6diFmyVE/RGjgP05+7p
Lqx8sSzHQl3PfiXQeNq10wkzRKiWBYWHdO1nZzPOyUq0P+ZwgB6aVX73wJI5lHVI0TN58Cph4tLb
3dULNUBquZ5akd+U896LTuLxInwYKViIo6srHVJ10sOm2NHjjRkPwDTUfg7QEfzc4noH/YsodsxA
XCUcMA4Z+8uddlbAhYtbhnzwGtvBIRmeQr27diuwzBvlVqjQOc5nNSimePx0T2xc5sjXmS3D3M1T
WscUJX3VLHzqPcADJVPns43pMS1v9N+9BxWJ9WLycmUkc8qCzdVSDr9ZJ8MNcq84pZl90RTAlos0
yUw9JZ6GawTzt6+ti0tJMnVetU/GMMvgcMlMLrHHANLpVI1ow0xJzA+99V2hzjGGbYXTCdQsCQGk
k0qvp+bIb/5qUiWzyFQj5SSNU6URh3g7TVadnAGAQ+Tw04rmX2sU3zLDCMSOa/Qrh0Rqx1tm7x+m
3YjAh6XpJesWlU06VuvI0cNysxqBmJJ6chr1Ilgrk/US8YZesQOmi9gLXRry78JaoOa10eDT6ZHH
Nqdl2u7Ow1pHE9Pb0WJ5AirAdTf+o+8z8ZjLiOa9CAPZkhcCMWgT9kP7sCBxqn5U/tg4uYZH0bqQ
2DeQ7kTOr55GOCnnNHvddp43u79xsB/xX4pI6Avlfwp5utjPoaCVBfyRRGQlWSEsXEMAj9HEwTyc
wl8qFSjp9c7Rwn8tprO8sSUTpnl+6lo8W7ehSALqALmDrgHaMHHP/+aXRKwY7MMQVMz2kx7UrywK
yFW2RTtv7V/4DavPr4shKFnxy2zb0DNSlr4z/n1M5OjxEghSqfqSj6RP32VpoYSuUxpC3iaUfbhC
Lo/F+cwsvCzkrFX6YRaM90w9BK+fB2PMHJ8aX7HfsdTe4J83r6SRuw4T9IJQFIbhiSdhuKrIrY36
SyQywThKHyMHAALophQjeKOamVOnfi/dsotLB9wW78Bg+VLIbq9U7zwG4TEgczGcvssY49Yc0g8f
0hJb+ijLxdCyMT1uX9nO9Mtn6acNd4OBxt+Hsb5524/22VJq5ky9cvVY2kAZvTaOdphXf9rxPoPp
56dUBTTVURhzmVjiLbPKPFJE3AddbzrjGK7LGc6ssWRussOFaTuB0K3aLSDiCqdRnvUDXaSUimZw
M7jjDblx2muVitdmxTf7dVW0xAvSP/Etn/JEV10uPiAxaI16ZMBdcqT/Y/e8p04SY8ls9dFs/0Tj
Fhz02/1a07rm8zogmuwFnfXmX7gBArDb9CRuSmDwEUqTTOtC0HbzQyfor+LPc6qw/ueZKU8aWgDu
k/0+5fdNe8N3WDOY0XWbpjGse7o4Zra1fhl2n949fb0A6E2agh3JgzRsw9uvLdmUdSJaKA/3tFzO
Ut92o/qbzBnmX3+AdV1DlVAekxmRKVHBgRAgcBYzG8vHlf80FcjwFLk6XlRWck5G5vmraO7WcymR
scHQN8RGNYgioTeZdkwTP0tzNPvzYjPTPQaxxohakswtSo/iJBtuKvlOudR8JtBq0ahbbVpNvy4p
2Stff3JbIlQQSXLA+V5w+YE71j46yV8QJj76gJtzG0UI6N1McZQEEXSyDx10i9nKFlCYdxfbUsIx
xOZfpfa8xEnkIz12P3OD/M4TM4PUctdy2jxd9o8DGl2fC86PBtm7LS/6/G1kUDf1UagOFaFBesv6
nlxVWbm3jP4dCLBfW4+bcpW7BmPKFPbu9zjRQfI20SdM34y4XvtvwwROfi9V6lzpJW0OGGdLanoM
n9WpRym6pddu9KPsiQ9h8miu9PM4EeF8aOJgFXeRyiaE/apEp7qCfgLFJ3/BKQAhjrOmcA3xEsHA
enoU8KUUKK2EIjPS8VikAvxGLyRohLa93YoCs6pQyzIdPOQ/SjQ8GrBNT0ZcGanOch0GUhWqcLiV
dr3peGOF0SupF4OztKssNEPJpVC4pTO0fwOCQx4/aGidSbPPhuEU+sE4et4PUncqr92M5HL48P5s
x1DMLHLkTPgrARzZ0xZTIm9GHs0kIWRDHwxuZCi0Eql4rBat5vvIAP9tYVu9faY8XoJFweX1vcgc
bKtZBo2YkxP1TKbns2kOOrS80O2YL4InW32D70IlGR8W2rysgGeIkzgr51xhUBKoxcdBZEsCRTkN
hy6U7TeiPg53WDWRLPaGseBT0MuCOmNaDq8WArnw86p1OaC/Ku204Fmnuyz/hC0D2+krr4QK43Bd
DXWZ7JZ4xEPpXze8QgJVNZTyj+80Jp8O0TE5x4EDJLwTmo2BJ1oflDDiRCPcGgEYYEgf++Gfl7j9
auNfHC3p8JBZJg6iLW3/RYiCI579MRCGkfplgwj3To8YVP7sYcJxW4SuSpUhYKxnOZpA5E9uoXQr
Y2hBUkXyaP8eGRhFHysC1hItEOMt4JO5Dxr3ACCWXgCkMBJv9l1q43bQCsnBlDJdmpJ2zFMRrzg3
79WjHLqcmx5nq8bwhV8UPR4jm6sPgzUGUTRcPXGOE5AgJkZNJ/D9mKp+nYZFbDguZNxvqRsOwE3M
C2tASU0YoMTHGW/0IpKyX2Ng+4ux3G9anpSIr+I/TaW9j9GJJ519HI6z/ZEcWzFNwpUMC+7y+zo8
x4pTlyNKxmGIQHnePT7zFp/8TMABAbqm1eCdbOKymEvY6sr/9qc5WMPomBxF4HxxsFcLGYv6b3uf
vsAPssg3L9sBZKSs5PdeO5gSLDFHYlUEzdwS0edNs+CLp4nh7eb7w/VYFwF3xhVvzLRl9/oOOHG0
4we0BaxKT8wb/A4nkZGef4fbSdWQLVuWH0gfQ77wNe1CZ+rh6vvKMYZEDirLsKTr3Tq1S63wWdy/
o5rVkQ3HDo/2KzuJNrWHOdQFBJISlHtnK5TIMlcO/80L/tM9YVhQ5b+B+XRupWjz7+jw+RYtf4qi
oh6iIZ7I7HMuZYsU+agUDs6ackR0/JjwRYg6ooBT0NiGJcJumq/Gr20W2I8j+EI/V1SelKvXcG1+
hs0zEIxql6HpZrQsB2fmzaqmbYA9GrnLIY7Tv99I+n8+KWXhcktwGMUZ/qEoO6tl4gKPJn49jkU+
tCr9kTKB3/7dodQe2nQ31F1LvVuVthrq2ngO+3IdWItcq+CjsCRwFQC0ldSEmN3GdbSl3SrQ5ty8
fF3JZw5aQ9sPBeAxPcvfw/h3oZ8fyJFtfZUUOpUv2ClNoyxLhIzJfpBM39EMgzrCK378Fqhq9YMq
C1ltuPXSmXLmyix3wMeAXJkDTy1YzNSUpGec6OZ8PBE/Jit9KyTFYcyTm42IdCysLpYUYIuB6a6X
5wGHyHVL5CCywhE4tM4GlXfkw/6AJmRIgBvP+mNk8yqynlTP+1e65QgC4JB7S73QCNfeaElHOL1G
vpj6ogjjMrFntGrRGoB4E55kmGzX/vd54e/g1kaflzg1eA706RrZg2aE94BFpG5MJRgVuzwfTMcF
Ut6DxuzegaOVAjVwFAQHg+dAAywgD5NU00XlVtIIyKVTzN714YVuEgrRwgFP/2/MvWE4yu1NCSTP
48vwxpdOwQBFdZfCpm77sRkWXuAAeKHnIIlGCgsGV1elaJkPNO2bzEbd8hAGbYLWRlyLD9DZw4x4
Pw256/rAz13nNQ63DWfh/N1sUm5cX4w8vuzUv/fstQgGPZLdWV67qGVfhNvTXT/mDrpVBPaoXMj6
RbiwyLlT9Kbg7+7NnmhK+ZnmlK+7T2X38gS2Inyc9/jEdw0w1+ojfEngkbhp3WFDajnFTNJVxq0E
IVNlRdtdJhJzn+8p7KlMnfXK3nnPwSvT3oH9G8mhNXvi9OqaqlcCbnKZaDUugV6bnDj8z2KRebcQ
iFEAFVmcSHxX6bdC16ZfOf7CHA3TuDVvFHePMO77J6/hNArxFvt299cbJoCjtjHDYoR5K6oQ8HnQ
JaRWIYrudMTnYjX9JMBlUEOAay7EII6DrwJvL2BAvvZUq3GFvJz+JEXY+rwLRMI8zAaxw3FahI7o
gw2TiSMsAw7n6B/rCJxyIed+muOkqkHV0P0A1FQLkZ7UHrlJY8pDgxfexIioeoAAu44Yjv5kdlRP
vDNvM5MRj9Q11Hk5wpaiIS4Zn4JiiAVDTqsvh0xRsL6kzUV3sYMDJQ1Rt1nt2YJqf59MjqILE31f
lrt1/5Cysp1x6W2TLl1gwoANnDVIKLpnA5r2tj2QQJOSTWtjiLCFPmyir3H1bncyQqHbxM8u+z3R
lHZHFZh7iwwIx0ATX6xOBMQG1I4U3rn89Egrc2cAam2xQhbyy88uUygDhxpYvYRoKs8lMgmTY7YG
t40E21FmwNHegNrHdxDgmG1shO2JjlR2iXSblV7KX3iE2xQTMGHY+ayThcL5JP19P8GVuphYtIok
T8lEvTUA7STdM8tbpUGw6EXbISgaV6bSgqh2tJMjFA47CGuMg1Bfgs1MdISl0nXLM7UlfRRRyerv
2cniZtfWWxwVrkkKAzMluHKPSiFkBqDHz/4jCEE8cS1HPZdKvvM0volug/Dkx6uLDRYe+AMMVVzW
xkNrKeU7vWyvjOi55maLE8s9zRY2kZmFnNId3nga8QxJXFkQDDeIULHA5t4uZKNaojSAPQ31RDCG
Eb8dvRBPu2fYR9aqoYjGwK/yLl/gwfL32WOdy9Y5C692kUgayuWeTtnBBE5UxuarLYCCESAvyIrv
vwInmz/0eSn4h6F/viiRKW8a4BO66p7dr8yCkIrPWojaByEYSNYs6saHBUQp9vEdwQFtD/lzL2e5
3xgjy+ygYDf0hx8nWUqFkZ6PoPMBPOLsgSFw+Jc+jib8sWZvEdVMB9jbK2aSLKjfoXRHWHUCHMnh
l85kHWnGP8soGs2j+FPjWn078YGqh5RPoOWNrcfcjyUbLRC0LWAmLt1ci1uFXuAxzOnzCmZQ/aPM
qWrbneX3i0aX3JhfA+Np3YAkUL0BD9gx4tIIwAGSM4VQPVfUvf4XjXAIOeNoQ1JOgv10fwcYcDYL
NVZtCjs/ONvqO7ilG7eyqEw/4wy63RUepi3sikMwMbNDNlefVnESCTs4H2zLrRfh785WFb5HJLWz
xH5A4trlsj4ajUvLXn9OeMgTbjrTV5YRTtuSEgoZLDN2VfKmujJ3H33xmeLojMiPlZvuxJD1bj2P
5QSt3XSZoqgh8fXnxWHyN6bGssa/rIddquCsCdN14yN1UL+nJnh0ajqX5lKWasZoaebI8b+gqq9V
KRH+yZFM4n3cpwZt1hrivK5bXcD09l+1t/r1fiOG1uLLKbAKayJq4Pnez/D2NMvPl+1UbW4rGd4C
PinLc9ZOw0A5eaQ3Rev871WLMnInUvfjFof5wEQRT05QoC7Z3u02MqINhUHfieMYX/VpWdjnsOxQ
QMc8WLs04t1KSnltILzcCOa7aTAJmHutbIFXKd5pCBgrHeSOHV66SvYVYjFjG8GnCEUPbUH4SXk5
lMPSvxVu6P6nFgjTzVAF/lMAHFGvRo3Yzh2Qol/D8C2ncRfeDL3MsXepFDlgX3xrU/3XDq+XMdbn
d/FsfQTMXGRsa/kroLKE1oh76J/s7ce5KW28gPOxc/ZHWIYNCb5MO8ndVVx6jjlVR7JtVbj5T9A2
VjlMsnV6J0oubc7AJALVk4BV1LhxUfnwkxfVHRpZoCPNadwvFmOmw8LRzlgY0y8ElRwtldyAkZ83
RScEWCddD4dnxhU+RBTDFFAtrXXzWY5H2z8tYu90K+SAxbm5PfIv5QWojHi/h9NmFZUhDPHYkukD
nXmmM7/3xYVqVmNrFcdHu2cmE8jKU74Y0cDirfnLDEVFTXpPn01QhfvFxSjFJjJ1yBKQAFgrbWCE
rkGYubFbxucEedoqN4p5npOSAcWY7Y4z4AEwxNiJ6dMIMUBIVtgP/S9lhGPZfFFw/beM1i6FYt+1
GZ5AMYLU0lQ592xhMULHDGaEQ8+6GbZOIW0nxwFxB5IsIgxc9iS7UI6v0Zto6cdzaYLbvG9DYRny
yqLjiTWgCd+fMDRtEMmrBWx7SJkb7PxI6ilfN2nIL/81Qldp8jWxVaea2L7gb5Moa6XiZ/qRybgf
5QuOgYCswHhHWzImstlEZGkEAs5pRWT89UqKl/aTpZ7hdOyC4BoGDtg7wVqW5jhtEp3JiJXD9utk
Gvo7b8cQfIVRMZQNxRCyW8/A1f4MlqX6ZZrtoSKEO/J40lLr1X55D5pjCdWOeXvWHAErGP+IdHnH
rLIt6sq6iAnIqSU5Qncv8qKZSj805se8cA46LM4M6txQzbpQ9f5GYTmWsh9O2mY9BaadVhZzJein
56jFbtrCbL1sBSygJO5bINVkgi7fr7lyrI9EsCeHMwMcZpSJW6li7oBEkIkOJjuy+CCNCVIiy3ZN
6WE07QrXTQaTvjiiJ6yxadfHfc2xsP4YLAiJPgraQhMJ3evpap7CaYQEtJhhod8RTUW+KUawWAqF
MfyDaoCCl3ru44sdpUnotzQve0pc6VfxvVpyE/H3gqiGVZKZ92MGbu8lb0dIHg21CQlrwU8/dkQY
jL3uwW/YetG045BK57kWa5voWSByl+mHXtbGCEhGA2x+gpA6WlnuL8sQwoWUgpm6rRF3AYcEfxht
iHdsELIY7xGgH/CiHvsnMm1tp7V6w2m93/a5hHWx+1C8rJR+cwIZD41mcn+pU2jjUuQdjIC7Gwrg
Enw+v2Dcp9njcUp4sRTSpF4mJQXlui6OLvn1M3/AGGbA1VZwanDcmhkJDqPnsv63560N/zzYa89M
n8QnpJTz2zxtQuDqThUwBPJb5nQGqcEnfD1CQK4v3v4jNAlUiSK2Ot8TC4EfxMvzg/1xEVXdnW+X
icuLiZX3X+QA33AXiNpei+hp5uJVPEjiJWS+y3PcwSCc8H7qJr1kVG2p210xwT1enxVPrxmZCzJc
q750aH+dwS5J6YkF0jiGbhLiJrMDacJY7cymSGC5brucxF+MN3uM88KhDRSJ6uVZz/nyXI7uz6Ba
DgrFIujhEIjqze1wX1a+ImWHsO1LwoTS8WS2q9iKvrCZU85PbCVmwBqtepo2k5XPRAAUE7l6fm/J
YtQs2BID7zwzR7cZf7+im5+NrqnJqfBdHA3zy9nAvhfQF7pXA0Sz75xwNVIm/bvlHOh3qwp+4JIR
FZAmHMUAUywj3JoaafjeyIGXPyeZrqykYqfMIhw01AmCPR2Qzce7XFRzd7BS8FPrfwjpSSv7xJMi
MldWBfUHTtoIT4HXTsFPFG86YynamY+5LyVsRhrVbkVB3g/wsY4jKTB4IJMXat5Aa0XtlsM+tsl7
WJbiZaoSVLO6/vJuTX9uHDfJFwqeNroxF/CVAvezqglN2VtdYoNeMsx1joCVdwMFvrDUDAtfEg2C
90M33qji+dYsLG/tNyFBRdeloKhg6kyGvoGe4aZoY4IVBDKUfBTEXQh6kkeQYFT9oVQbfaxg9UJj
O2+9wIB8zPYOOPudC+JmKAobulNgHWD5th1LWMKFinfVBCapb3r//cXKq+LGuP0HuLqq6vbItWQv
+5litTuVsBlkd0SU7kZS119tSqJA9jPad3oxhmGuQ36t1ZfYAni7Ib92mujREexAVOfCHEJ7LyRe
ftu7hriCl2zcs4msukqvAoE9Whv87IgWcAuDJF45Rr9C17n7DrdKyVKzA7H5xkE6DpsBNTIjTCff
QSgSMmalYv/uy6tD6PkDP+plTS7wkfuaKzTo9EQXTmeyznwkIytwe1LSdxE/XTsMqRsEioJcgmxL
LxuIHU0i/B72HRb71lgkcYEGAg1K2IQm1ktllUESASVwte+yoOxWcCuZkyN8dQQOA9cZf3iQ2rMf
jo8poxsoffyCVws/48RDuP5F8fLjFdJvVS2BpEBtfl2T02hCik2KZWZKywKobMhWS2UBy1lQIG/5
2iPCPJDERIzoQiwP1E0Do+7u1O+xWFjy2/XnRnSA9rzCwtSFexVMbnuqo6TNkMCjBvdHBJbFm0vj
X3ixgYoCqBzsM3ripisNTK+jySC9xqq8uRcxOhXzYJtBlvZAXsAlVQhjbKwYH4k0igaWwgq/vax5
aZxYer32HeDJdHzOJbnWxXn04pLHRA7f4W+Ym6CzXW/AR5XopRQmW978b1TQZqX8+TmfvBa8XSEE
e0+e2Am1+IDUbKl84fPznLs/d6FBPBvkr6dUrQKwoCBpIVTTfi6Re3Ppk1XUkoAucX85e9WRVYvM
a6H8kHsYAonMbbZIcQ3yiLk4hsRYIVFNhNqGdFJzU9Fg2b/hYqut2qkVCnRiMDBeKw5Lu6Ckra+/
ihUx8Pemm+v6kCPgN278nIYnWJkNw+m8fLcvUvfDZ3OUimg+kKonBrjJ5xlGjZCN7xDu6jdOgXlD
l0AqdCP+iro0Gssu7vimhoUmUqRN2211GAU/mY+AJ/9nxRhVa5gsqkF/KB0ijT0vBoAFZkaeplPz
YuUsPkgChZO/sCkzVLabwfjATflmvxITniPzObkcUuJo9mV4S5U02EXnw7gvMzix3zlczIgGgP/E
suMS/gf4lVS/JIwk5mq50P7AxmajW0+unGPYwH79Z6RqaCnaSU3+pv4WojSvc5clEfG2EAqroUK5
zt1lDkUGRe8d9mhVj5rHXKOLNljOb/0Lbl9g692ebPlGHCOfpco1BGFxzYGWRddcG7lzcYfHFeEB
cwPKjN6MDOu/PqzFHqyYaCy1chHWQHgod2GGEt3yh+Yg5NJg48x5iPAQ81L91kwEN4T0nVUmJA9y
1d5lwfS3Do5VZIszSaP/F03JdzODgBWp8D8xiNzLwl/i7fbFhBXGz/zuk/yXPIqidh0sUU9Ab1rH
U/DkGOpaHArQPt5cUbbfi6vAxw0V9YjZhyQTLbK4FLIEjWJq2wi1HGlabyNpnuKm/OHIUFarpEtM
SAf8t8qx4RaQ4UKLHzaQrZ3IaKc1uGg2UO/MZpxqX2Opa+UtcQxY1IaMSJhovY1fVyr423OWM19G
iYym3th6qsh3HPmMYXHQ2JHXTRWkQ8Iso2G2VELFdkuNRAl+yWYQQELdAleYIStazCILP8hYimF4
LrlUiN9WzeK4XANF7EBXsGPrFOWXkFPz84yezdrzb80kov1/q/+P9nEoXCjMWFRV7XgadQVafg4Q
mbNC91m1yZ5LHHc+1R2F6VH9eScxEcZfqI/86ZcmEwcyW0YuiI2uzpTNnYsgSFgn2rtdc7ZLQH3A
ckSH8m8gz7fy3ihaVto9fOTkPnN7pvrUt//i1coZjttifKKCUBlQHmlko8SJn3+TSKTeaKY7ZBNt
Qwj1OUjwEhxxmJ6LiCFwOOf4jjE/uQlccnXxWvyTxYYMzmyfQwShcV+JuKLPvljcL8itBDF4tq+R
8lOIiCzBUwk1wONEvSLemknLj8jzKrjaM8MkAojQPFjZSOIDpm9vwbcoATAAFn49Vz0svvhnKLbG
GAqaO0d48qc6hLfBgWVvtB7+jFWbpSE82GZmL8gayrDIqXQaRQoKDuHVY/+bRHzGtKV0Bt3coCto
dPH70A1Q2C1kZv1bwRDAh+uD09T/Wf3mtQoLLhaTfr7UufQ8x0rO38+BU33P2M2xXbEq/9AXWZZO
2E6tvtWSbDwqD0U9VyLqarEh/OW4Jtkon37an/5spcx6+lIRRFtl0DEbHv8i5OoST+HZSBfl66K3
ZAW3O0PFENpzajmy+M39IuyPwIzV3Vs1V3LtPfspDsJ1tHCi+sa9geyQWvLIUPajrRCtOZ/i3SlG
tMFrYgzTKaSF1R7ArNH7ISBtixTmU7luINE3l0xU1bPuAJU4YS4Zmv7zGP/cICwGb4Vv33VI7XCx
1P2Ww2Clhj1XsPSDx8FyBkBxrYgxTh3EqX18kRCOHoYEyDvth3XRxOu/TRuGFcg5h2KP4Uy67/eU
qre6I+x166NLpBZ3oPc+ANOhFF8KzyVHU/SeQyOvNwNhUzDXKx1Kat2pteLlsRvDn9OIGRFYen0c
mn2IJMfNA4wgxKSVE7P/YOn1OBX/co9yvIsyw/JA2dt5UQPURYv2xKoxQPye6teEej+ccfg01iLr
WlwZAI/r+Xgc1NieY7urxdD3cy5vIP14XX6ohGHarvmBoHY/EfyK+vq3EyQKdiJBhOZqcLiRFadj
oqI4maQNC04QXgcO9ZBfjJzdXMYVV0Eem+lbo6bLFXrdThd3i6+67kzW69eJWfqFeYjLteHsTEq6
PTK+UhkH0rSktgfTPDf3ezWH82w4Jie48CdjSa9tksBLaqLV6vrs8SIB1oxgp7xLiL77G6azKklM
gP5F2D2URiskCy6OogXt+ImjLHLCiJocSVFQhOwy4qCM7drmWX7RV8c/pFd3FQ5L5IE/KG5JA2Uz
9C2IrUpwzOnSZwk9of6UR7pOnvHC54QoloXCLw5cpEaYITIo4nVZbtrLOXL9i3LUeUVhhAvS8E66
U+kV4G9tCdLTlbj6b0TJ9CPf1Yzleoe/nIZLT9HqqBlDHJbg3HfokNH/ntYP2MnDD/kCrEKdJYiw
3jIWdNGHY4zMyxVvy9yf4ZeAS/G57J9gTp2s8usdD1DWiitN8cIsBB9pQ8Nmuie/8rslhOYXD0mA
tktZ1EtMwb4WAx9KBoOJVaOc7vV0Ofy6hCdiw0BJZf4Bbt7ZSA/RGBYDjpcSPa2AHPHI5LliE93i
t8Sw8VEkjLog1An94YjnlN/oJDGeKZ0QNPlXD5PSdo/j/FOLjCam1usGwws4zgEsWywI6NyyqKwy
ktnGoETa2DcFTvTuJ1t0sDpA4oyO81T6q9y9AERQF0fzWo8INEtjkZMVpcltR23Dzu5QFwgEs/eX
tonjawsOS+EHL+39NF+s1+5mW6jLSUGFCwgVAmNcD7dxlAbzFP6AYCNtkmobxOG6Pwrvq6kYsqAZ
PjA3/84VnbL5S1qqfhDjAzmHpwhwslEALzQC5bOT51rE9jcQ5rUqnXN0ZoIv1xX6kFrv+2gpr9m6
LEKpRRYseX+N/qPqIRO/EJWhWEkRE8Rpq8+r0bgl1VBm26x92LF+bGh1wm9m2Fq8eExw2h5yAY0A
byvfnUlUw/gIGNQvOcBlnITMh/4YM7Jh5g6Qce2GqviyYXkHgient0fBvCnB55DkuyU3I/vs35nN
MTRtIC7GMwR4CqZHwBkv41ahcbipL5H5cj+FCIf47hj09TQjr014j4B+n/4KOnega0g1pzMpMlY6
+vbOcZwNYcYrcdz0zIZhNqCy9hPALtGh3leD/BR7FNotoQne7YmuluDKVcCC2B1weQfHLfNj1gyN
ecKb83rvZ6HKIySE8stJm1UeqKn56461NLB9P5NiKhKaN0+FXMS/hSMiDBp7YtDGGLRBQAN9Nl0v
o6BFzJaJtuQ+jH860n9W2ZEGqzlNIY1f4FlWpIAufyo43/7khSoFTeGs+WoTqJ3t6PHaBXCDRiT9
Z8bq25S6qJ9lcVHarVrVSjwFpncGWX51kzo8GdNscruv6CPEdDjuiIuvZDUGyvESpQG6/eC04AwG
E4ymqIStWDSUteh08sUT49pn65lq0nKM3oszz3SGu8N9GyTp71rPozy9bC+ituV3mZjg2thbzQJj
ADo7jJCOFhUpmVpQPfkH0gPRN/3oGe83UKmsAKcYDSMuaxSmKHAn2s5u09JfdVLQjoV+cAx9QhtL
Fk389HJnURXgI6mz+RaytZadBDYuGmWIQiz6yww3Nv4YZwO8SNZeBot0Cje5+yI7rNyTk4xTdoD6
W+PYkTjPA4HWGYovltccPAie1klG9iWhTIqyVtdJrYfQXXp25zTVhHNBboa5CmqaczrPr3zLY4J+
xy3w2B/AcLqvEYbooU7d5Ug/ODOmQoMo4RK3qT2tOXOBGgAMRtkgkiShUnbwbNbFcG7CXTxeHB1H
TiTD5GT2lJ+tKIjbWstI72wlCsuaLKjDyjzKNQ+auA31ihafHY5RD0SOku0WH9hPOJXdHmcqgAeE
M5DsWwrNZbaCISJ2gIpQmS+7a2QKJ4pibK97me0LxaMpO4oElLkavxeZmk5Dv5OSUOYHn9Rpd1K8
N7CW2YJ2p8Jd0bulC51niIQqLSKFjbLRRRBKlYgVn3pFpcaEN6P1r4eeddkygfqd8Sc7RPwDY6kh
hCiFaA1iE1vmOB43odol4P9P0fTG4+6mWIAc+ljF5oTqQKFYWRUiCoSlO8n+c38YSg0kr0xoQrqz
hfs8z36zwuxdnP25Wso3z1A7h2NH6UJf6RH6jGJ7sHAlGwb/6Fc+t9Y4xu4GBGwnF/ElUmY1qff7
E0vSBRKwuVC42UN7MODCzxB8/HTJa3r0M5pTmBAWPuefymNvZDSf4UsU74sabSou5uOdiB4PnOg+
dEiRqreDwgmaGoYDupLGnriFXRUmGwssNa5rXiIoNrCDGG6/xUhUTKBsl/GVWoqE291rVPK4W3Vb
3gYXOObYZG3LH7Aioti7bK7luaJGMIyqV4AfCG/comuh7uFcIEMKWy3mhsWoyG43VukVJAzGZs+e
pz1z6857klVtIX0OrKx6AE1unw2NMc0EY692ZLWil8zngfe+GuAJecBzC0gUSaBIr3ycZCxesHOx
uPYI+zotOQpKZm16Z8JOsjfTcU+iK08qE0FWtKz3M3pl1OFprQv2HYKUF4tNFQYYREM22FTyI60c
MD1q1HUJ/du53L6QRoYd7Isix/Q8pJcJGx97qJ/a0FwXYJYp0zD912tiGZD4Zc0Xe2XwGz+XaL/N
zqdkNIynB5A30BnxgsaEIuhGJY+RdH2KthlfCb1CHrkpC0+HgPo/rMSimyJ0tg7rJjfP/twNUFTG
Tw87RSC88oia2oFmPlZ/LZieVwhuwO+Vhh8uOs+mOV43BQfuuoGGYkDtMPCr2FQ7C0/YR5jo8jhi
j4aYL09oCUsfq1q0F+4WcAgNvea2pAJzA1G8xT/RiGK/uGsNjvsEBPP5H5hGZjGsJdFZ5ddvSPe7
K5f/Bj4SDXvf6Of8iOKNd+4SiQTWjf+wSjUMC02106xw6MHQQ15ekWzqnT0Qstl4N28R8XzrT/pl
hL4n8Zoqeln0OibKHBU9/2Tcvb/cVmK0ectlFPqjFr3wTAuncgCV/WR6kSZl0uiJPC5sXN4WMc2d
TT+AZ2wXSk2m5JwGGly9LaSK7JOS9Q1c/x6yd6EYgqUti/nGB2znXrAVqXnX6krcX5qeujyKX8/J
y7qsq+/I0W91O2hcNeySjw8CFmT4wTK9bDpVjQE40PWSKEUp503EGKIqK8hcSghN65sam/ylQnn7
xJo5kOeCbfemQOH3F3094oixCWObM9vLZpnRtku5WwnriY9NB5LDwo++v04ADRfMQ9jB+r3+FYeA
z0Sd6XopwLWTi6+4sFBz6Cnt5Ggyh6069hZWPkKs54tbdi/kWQ8IxdIwrVRexrIuijkfduuGBWO8
HB9xjRlRe8+4uEvDGsmZgvOOFlxc9NNrAaptK4ndm/Nel9Hj36BVht2NoRJOx5KLq2JlUdV6mUKg
l8dFwrSzgH+/863bCAdx2TynIRSAzn9fJm5hmIYxWxBmn0DdYKnLFuyAlm8HDuzWa+ewWiLOqmIl
IwlPe+E6CWSCeTGjAUaupW5wr5kBSmTBY7CCWboG1J5lajNy2cxouwkx4IDXQ7LOWj3Ad2LArPS3
x3V/1VzJtq21EO0anlok57nA5UdJ3x+WJUcVTHtFqfYcBcDyhNQgbPnshHxDyqbSPhvQLTXK81pl
okFXG5KW7MssHJuprIK0gUK4S8cSBLB5oOhQQqEHD7us3GHX5Zi8IATIdLY7hwl6MZLRiJ8VkH7q
RPcNhVLMLTj3O2SGFCwdzTnL8ci9cIQEK3jym3KWBriB3o93aIghIavyMq6PWIfURezX/3574jwj
unIH5WdrvoT3FmDepDuAF7M8jlWgPtTOoc3Kow2+CW//ZX531eSbKq+r1jRWCLNqgSAwb7Hk/krM
/EyUWxlLu+BLru8JnrNcidL1ANI/8Ux8pcCxs6RwhgVTaa8GrJ2/mwrxw19AHZKZCseyXPuhB/uG
wkTov5imRJyW4k95Gl8QCuWT8cQy9fIiE1HGNjGYvsMKf4MZU3hB4idGxwSDiKMnA4fGg/xb4tKe
Hh9EDXIVJjPOsZrMI2+pdxWc/ZRwl+kWGfJJp28YCz7rwikfA/HB4N/IoVEW3MTr2oyxm8RvEoUZ
ho9elgR+ihJ8uPI8btINOmxd/GGQWp2N54szBH3aRDqbinj6Rj8bVpRiammXHJtYOZgiMjn+MZEk
Oy1LLYAvuyX3UJKhuvZC8ujjW27ykuGqkJx/Es4MS0pX50umFmMv6SKRecf0hv4oiwg8fAztQzsA
l3CxtGOmKqHXTqm+Rbfx3BeZLJ7B75CRBGaCn8b/MJOIuKjaJ+LBINB3RdnUGhkrSx/enm3RDsO0
7yko7ArbKZ6FIhJl8JbJm40jEyBphFOjVqNnqeSRgUyID5bjbI8d1oyIPg1c8F/4RB95v6T2X7MI
0X70b5B4KKVYttIVdIzl9ExzkF3uLMuvpQqT3e2l0Ikjmq4Hc4JfQuELVMwjGRzbfFuuic9I7DjW
AM+Saj4VEsrj/qqTXqWtu/yo+jnJEfT6CfQuzk7AwpQpFCeCz9prorSf8btYPms4oUikkZpq+Z28
VxOaTJRYJZOlcBBAV5xq08gLbBFBvmsr+cqSssr5trNNoGTqa2Y4NdLYmBCSAQyy239fbOhcMQji
2LSuCbntz/UwCdHFxwfq4mGysxK70t7d6HC8UR4EK2MGduPXb4BgpqaJnYHw+ZzJxeSMwHT67Hel
TSpgMvM/4INyJvGhjqc/gAOdtzoy6Gy2m7gqJ88TEVU0D62wxsw7KhqJKd5OwuMyoR0acB4/4U5/
fWioMaxtkO+8fa12QzxU1HfsKa/VletXKadceoxYZKcVDUghXyAQVIArCFuRPKMxDaEqDh8U0X8S
/qzQ+mbQnBiF/6BGgY2CQFifbBQT9TIbxa06uEdzDUCXFXckYMPZjJrydy9/wglv63NCa22wise6
S79LNK1kRttRTxv7gtvVYv6Q7vGdcNdVm2ESa3eIa1goRA8IKFYuEc+aRiArgZ1LCd3lBDAC+5W8
69pRuncAnzLKVTJ3/D1Olv6yW0KAtOZ8unDf6R/hpwbBy0mJH0d/jBedjmc4PWNjoo3Nn0/yKWKm
RJGgTlHaKlMlw5z8ZJRunbFa6p7MKuZTvRsfTjS2/tUTClyrfMLCGN23bF0cD/cVEtX3TOzJpWrW
7LtHuEn2OId5L1UFuFfGq/NVJccr6NCslkhdjlmAFLbd6iKEHTFZRkGwK1Yes8n2BnOZ3vmEiA/s
hRlh3D/RXrDDqCCY0w78rwubzTsVm84jYVLUf6gZnDYSLndES0n27SYpN1bmZvvsPDa77jZ3O4fl
vMnm07ImHDY4RAwkjta3ilYOP6BJsh/CcccOU9iannNf7Hs/jFij+6i8iDPEQc/ThO0rBjChn+z4
hYmRkTe8R4mBl+/LIE6ILiqIW4ykv/t+YWsf2w/jA0rKvsKlN/yUKaCv/C6j7Hc46Kqq0VF8Le2j
LuSMdR1k6HlaA1ef7ZNUAUT22LwzuUOZNy8ufjNMTTWVMurXuVbBkofYtPKZsiOwJpfHhygYxinM
rvKKlT0w7U/UQRvKC+fj/5MQg2HdCXiOADmoHHQuFznHXEvabLrMYgFuUalkBjtyl3lJLgJdRaBi
+ZqPgkX0xpDQlK9lYqj9tj0/YOpdTcjjWxZCor53Cb1tcnGPuqfsjlsfPKTxvhf2W0SqXyk9vCyi
CC+1+UUvzy/UTpWjeTKihz63vh/zAdKkukvs2FX98mUBDMsftUxnqKYhERUNZcDWFx44YVetjW50
GZE/znrMgPNRQpJYeRkKVQ3pCw0MuUGPCaOq7c8ABnEsLb30bqkjwFjuwKquGCWfNvYwTi+inmc5
5Qu5WWB6+4JsL9Qm3SEK1F9X4pT30uOCTDqvvoyjz2bqfdQcdUcIygne05n8cVBq7j6TWhN74Z9G
0UVO5/VDyK537qEQGJk/BvdTosPLqat9ePZ2eJ2loUVCKlBtkNepYXUWBq95efy6aQKa6ellCuL9
+cgBOpAb6g5EJ4/++qNT0qD4LCyT6J5ANHit1mJ1ullmoHYBNRjQYewgTUTOnFgsHCQWRPbMnA1Z
Pw5V+8/W35/EF6NTufBkEEhnbX9h4E6geJJNYctER+cFvWTUYzaquBR3g25UebdLx9C4l68j7oCM
bZu8PQLM6xtWTeXySf173mhb9ZkumLlRCgf9kYP9/x55d9gknxuVCvl/AT842FSc2ic1Y77WI0hg
2QMmLUg+yRKMca8OvdOvsizxIXECOO1c8ElLDz0aSqOxACb15EOrAQgFX5JbUQDaX7Nu4rHWb06h
mH04k6O1FF3hXP4fn0cDIBhSM/PiZswOKfQYcMgr/N192XXjSEggugIMoJy6j4b4lbSJQwShv600
W30SsY8dH8PbjfSvAzKfYAyNXhXvBaPgYGCbYw+mooNyuVB91Ku+P0D9Pm/Frcf+JQLGjgV0gZCw
5+GZUVcyt8o6k7ehUfzPt6lFdgk+sT8rMUt0cVt4oIp/dQqrAywKGYGtcrwT6uaDIr3sRF2vZ8Ml
R7GGp67DiD6pA64/lOE5TLtC1ZZXnnYjy4JAnAgAifgVOMFUqyK4Fkq/lZLWjLUzTIY5Mrw3dymU
j2+IV7TtsAFWjSF6CVchd5Pdkn/6BdriBIbJnTWa7M8Hc7giB+isszWBOY2domk2+w52mwN6txdh
aar9Pv5uGd5pLniHeRtIzAbKDJ5AC/z588SqDdjy/MfTHMy6JKaHj9a15XCDNOvXwj531keQGXEY
qla8gn0pJtizGoqhQke0XvOhj4w+ZjXMvPhxQV4h1RkilnIMQ2vgNge9UKVUjrQcsov/Wqgs8Qva
aDwdOd6+KzZE6g77X0IuTzMgoH1INuIqxKq4e3Vf0HUIxBzox3fJi72ZdeEJHQX9jLuFK/TGvoVn
fIZCrBA+sg7ZlhsyyRnGVXbq2UhGbRzAuf5ontEhw7HaeUXlUM4RDPsFzNGusO86HsXPEhQCWmpz
yAEOMf+1o/aQI4OVNFXRMLJzfKpZqXokach1blJSwaEvhtco5UkKg/5/6bhW9Hbba5SeITaFRhPv
MtYXMHq1Sna++6cTCIXAOKI6LMzvuT1/bgsOH/309va87PB0Zm98NhbzhpkCCm6KrR8PPI4s57E0
GdcDNtthrfCvtE3XaIEdS0nOIyrfrdxyhyLPQBkeGWeSxgaT7/3/2OWYx79q0V3b5OmgpiG37OVx
18+dSg3Qtm1yO2TgU3gOxsOkD9MZL6rEHWcXFOY3rBbN2TrwAKLcGDc9U9uOLbf7EEBQKBnguox2
TfW35k5nvrxnh5Q80HaAh04gr6FKFSeY95LzcfH6d38q3XV3f1Bfzp3eD9iKcW36o7rlpFTGRjTC
N+gGTXV4Y01Xmft4KQcHCiw13Bfbk0XYOuqP8ev30Dw14QpQgkMMHOCIP6Z5vT4RXaw1H2VsxB5a
GBelJX3c02FDd0sGXI8wPCJSIhTC8FmXsH/0x2dTfRyb1/ZygAmKI/G3ruczT7gxDJ9B9XdWglk+
2EFUmD4GQXzGybTP3ufj/YqLG9Lw+cy7n68cMexZywZ9dOO2zzrU0IOQrD3+IlYHOVw5Auc+qLB1
scvmoaCW5W8/ugkADesQJUKzZUokyudIOREdGofzSZXmQj9RbqDsdJ72IppcsaLnlJFulxUh8Fma
N/RhTLX9hy5x9p4Xrvlc2GgtaAwzATQaIihKpXrm68T6K2fDFww6XdwmYCe83aeKlaOKMbVdzk2i
mSuTLUtXD6P6rvQmdkiKnn040u8C1OX75oDDzII3xttN8dZI3ibpMDZqoKchjYBAcCFRnNH5J1pa
8aAd0li95GzlZEXe/LpCqJEfwDmE1/ralqqR7spLS5LXG9T6rvu4ZhuZvUuUX0CTc6UQ0Els6dX9
lJG/NO5Pxn/WNbSbMDo5woalw6Sd2RftRB0eXVByQAGkmvYT3Jpsvv/aqGyMcpCEKBY9Cy8Z4c1c
nQP2z+ZF51UpI31PFloVJb6G9lwpjUrbI4UPIBnxDnnMMuciwV/j10rj/X9Op9eWoGTPBtbXG/IU
niYKQrNOc+HDWLRx/n0CVsQgBhrAUMaw9YC0DkIP8hCv+GrCbehyzAuSIz4z5pkEpEVh0xkR1ipl
rElKdMQjVCPIltHE+SthY4bL9i0PnF37+4xDo2wMP13OWzdqkd6JqCmQV+TP3N6xdLr5Q83g0f/o
2CCVwwms90TISATrI4MPzeSBFqFRsqec4ietyAFTKU9EI2PlNCJt9xtFjAJFmnRyltWZKH1CTdNJ
l4QvrNXDjICypf2AmHHz4dKTdLPDT/duz1RZoycdih23dETa8mEQ7rKFAeCZI1QK2OnrChjpf7Ax
fJdcwOwIC6xeOsSkzejImEnjMmCQLpKea9a+J7Kgqb4dVmCFsSLx4eSYZI1i+lrW2cQubaeH8WsW
ZxjU/pX6FxEhQyhyDA8TAgNsSGgYLJvF00bmHzO93zng2s+YvmhRH98H44lxJFCXVmfQhswE89cm
rXG3xKUeikbPou16fsoDD166uvdierWa4jMEHZ1cFqGE+47glKVO23ocpuj8xavOJL4kKZ7pd0ix
erL2N6MhqENxC5GaRInHpz/CJ6Wsg27LHWryE3j/fEtTtyxcqMcXDOuo9LEKlGklAyKW3ju2fGu6
5s0kvovPvwSOZheKIun+yg5Fv2ii8mcc2VILSYaGTgXmBUrTN6Pj3wtG/tkhTPnCyM3I1++KDA8I
wxYdT6OR2ynMQ1zIFLiBo1/krKM03HdpGqlXiQF/B1ALrJrHunLdngTk17LSa6vHtEn+VucBduf9
s/lEtBsMcTXB9fvK/1TTmsDY5Zva+SzLs2O44ovqvr/IZzB2yQaecy+YiePqQIfGxmNA383tmzc6
f9VUmXBvUmPQLtIjQWN8NcwnONobLI5HV9be+SH7cYWsOdX2WcjwX8a9L79220ZBJ3y6HHfZFl+t
u5ajT/AYiwWS1sn5cmWQsIm74Qt/GYYC+NGRODQrLk5MXJEfDlQvRrq6xL0mnaiUW8HhNRg/qdKv
2JdQOa2nOZ5C/HNu7dvUINrz9/e7KJ0EG0MqcRaJqBswHT/yvQj4vuYqNZLjG4r6a7P4kOcyox+R
2fAdx7yVfdM7DPRkILSA0bQvUc+pdLdGxuQpI5v0PpwgcRc+47yK/OMOy/MlDsh1YPYmLXe2sBgn
rYEhi39HMHkM1Panp64E3BHjB2NI3K0+2j65UMp0c5s/CYW2zR3HITepmZMF1dzUksA9G/guv1dX
vIMq0krlOVtZYP41P/PhC+brRM07AjlWOD74iMkLNEA9HAkITICfh7Y1DdJES6DqTsg6tLyjVPc2
UV3hWWb+XUDHsMmah5ySTTCg8TShglSNsfJe0RzdTs7avSx8vNKhTrqSMs3XK47U9PTmAT/cp8vs
0NrJ+PdSy/GvpdM4PiKqj+tE0adkLZnA1x+q7sPEu9jB6ISU2uhle8UXCDDKvU6Vp+dAJm7Uwm91
bZbv7EfKOybaBmSI0eTupULVHHCHKQAXs5jVa0BOaAeiUp3fzkKjbMR2237k0tF2jiha7VB5+/TS
1LjO94Ex2apSayYiu0HNiLOrdXJOOe4S3kN2jK+WsA69XaSoAQNve4+2721/uSZH/E4bcuiLR+iL
bxRDPeKhzGjyB8uTQNFYncW0qedK0JPY/ucvXeeK0467uqfP3MMa6ccjY60hnJy/OK/oNWeftyxf
Pah1SeKsFOq66gyOMc7cRx7abr6MoZGsJ2uBy1IH1SuDWny6sscMjbzFJvehjDaubGQJGXpBMDkQ
iPZTmuFjhACfNbRvHu+15GjPrpjumNt2Fafau1U8KkVJPf9gxV16tJNGYtd2rz4O+R781cSMhMcM
ord9p8MaTxSA56Y4VJ/YkjF4g4J7thHqv2QIBQPAIh3sLD/NLjWCp7K1h2SRqO6k+lxtNkBfaY1V
qS9vyHohEjddPB0vNno+tf1Vqvth7Gwj4Qz1lIcxN+5+tx0H9M/InBu+Tz7A23REl6Xr8TwduI5T
YizEbr/xT9pCuoxR17Z/ymjVae4ee8oXrQEqirTlpziv7uOkrbwXh2pPtSmo4qxkBl9KF2oKLmxL
lh4fXrG4ropj0FvlsZq/RCGkv7b4B5ie3vOmBYc789cPYDNS8ki7psOj4zSLmMYc7BD2LuL7gyrv
66VSmiHIv334hvVwqkkLvqAW/HPIraNvFy0DOIut5yYih4u1YKHRFe+w4dyXbBm43YepfoER7baO
ipNYCgUOjlPe3vRaAjuUK0SaIZqCdabofB6p7GGt+FU3f67A1N8AlWpFBEVk9eVZuDE8FG5+zdSP
Ae1DJZ43iL3Gcuur7itFlztt/7DUDyu6f5n7zx0gBLKNcXKkd2kLozFANAAb7aIfL0TLMcgjVxxC
RjjP/HLKS3zNRdeCo3YGv3AoI1lmlTQKxzcoaqj04MtaY2dgZosg8K8PFukOi4SmmE2ukEe5gZG1
N1Efn+M5TkT7H3RijKVqBXeamZB/YFmuZxStgo2kXrtZyqeO8hnVN6Z93gxRlAHFQnuwwENhD6XC
Ordq27pfEcvwLfq1OIZhAVbYyPHgN5JrHDOEA69nn27Xotu5tPNfEg1VhetX9Ncpq9/KI4FGvx+l
FbbFKRTL8HlKNHPFBC1M7qF4kaplqETEVE/tlCFCIn4avpM9Ks/C0hbTk8qzhpAVzmbFFrni+sCf
soLKHpkN6pkG7HEbrpnL5/sZxAkOL/Bc4JyGcBYJkPsoa+bVrHnmz+X2bBe3Ax+1IM5EjQNNPKOa
1MrriN15OMS/wjegrUjbW9UJ9ivNtRHMbf4++y1UQWRQ5Tw2SbeSpxFvgmbNwYBtkyHrK+LZ5NIx
SCToUEO/inquu5LJv3BXm9YzdKcgBb+1ad4aJGuOb30xNI0dY2tTUQVpQWhP2khsLYs1L0BCCSet
kr96JyoqbHA76jcQYppyliwSaH9Xg1/0LA3wzraSm3TSKSixmlFv0z1qQ5nifiSN4cMfxm2lebJU
oMOAgd49MjHybC2+glSIDnGhjdeLkAbiSbrK/7InI+n1kbJZExnlT2NyVB0lz78AlaeZEcsSjB7w
XSLSzbZKirScb8EthkKUTbDeDqP7OqeJLGYgoyHoptQ/NfNOFESXjWoWZsoY8k3GJ3bTf/Xd8ZOa
L+Vzq4b+NxL76g3+jNpmhmYKBmjFfACUqvoKDnCI+V0RPYDBNG2vBCJbVnmLriAVewE8lKj3wiea
3C2qMFx9ALYo0EZZuwv4ooRq4h9B0Ed48TFunVJVdP18LVzNQurAClV0CZth2dMHBdUs0S2EHHBj
BF5wlsjoTAhRbKXblTkFOgnI/Ir07oh0eGZMwUiDfjFA6Nd7fknFFBEwac6LUGHSkdLIG1WUOY2j
MlYcmEoluFNBuBs8pKkCpQpxlaSoLw9qrqCp2UVFlbDLmRpyxIIAmWqFvEwOCX0/PSP1mp6uOpSX
rgWsIc/ejvKjXSgdQMaA8dNR9mF3ucO7J3qk9Y7hJUIgPWKwMau2xedJdNsu/yXfgqfSdPFLXIfz
XGovS8IiDJMWPZEXa+2FpBq0PXyqxgSBa8vkJLmPGPYK9Xm1Us5NVi24B1HDAe2ysNnn1RCB1ymz
UDXzyv/z0tPWh9EqDL2VndnF1VVSATqkI8KaVg8sW7T47HWB2HQtH/cdmoWg2SkLzys5GOvbg+sS
m8jRu4WPRNi/KYf5W9KqsxFkmwTX1vRwwt0VCYccV6JaB+UhhFY1uuw/cVwlcbxZT7YCis1T59A1
OJ71RBWNSwVH/XkYjFyoCHbWpl6zPDrRqpKJgO/SFHzqvncEtKx9cpexSS+XuuieoMHRVo7FnGQB
fY0BqS0K+xMUwZs/VTR0kyF9WYeRxMDYGWOeLepD4IC8f4jlCK+M99fTTFI6FeFFghAWYDGOkdDP
89+phENEEPJNanxFIQuEwTVWWqlB2mEMAj9rsWb5FisCGSE1MvhuS/JrS/NtPvXCqeWjS0bVzBoV
oVEWngrKeKY9GC0kKg9l9Inb2gyhQYvVa/IDXH5CD9HeTwLl/Pdd8yash4ri55u6ZzuOBFDT05SN
gtslASoX27a+z6lWvMG32bvQXKydywvzF8DZyzvxG0/XYM19Dhv2GRwtA/NKZRCP48KVsH5oD39L
JPycce20s8x6oDPuoLOnvOYSVLp0mTUCohzUyqO33HJrqCzpW92FJuW54MB3iJf38HCX3H/TIyrM
H/ZDcISUXGB3vy6zjLP0WXrSrtbSraoz2PPBHOcy4vFyRkvjMnIxy6Ly6zg8wSP3b76xGnBCRaPo
PQQj/RuUuqPuvpxxb1Qh/7GbUDTAnV4OeqcKkposP8U1kYcs2O5uaB1GaUKy9nKF5tRFU0RMoKWI
MgHICAi6nIN7Lur1Ah7PXGc91eqEkca4Q7mMvxI9NDlWXye0JVBjXyL/y8zANEoKPItX8/DLaTg+
EZlxIaPj/EpnyrJ+kv311rQT96xlfFSuFX9z1LrL5I6+0fL/KYdiOStb/XwCrv5MftU8f9tR/lmJ
uhGuu1I0G7Lufg0ZGUpZlLjggfIe60vwKixvPui3NVzTFtPoYxFuD1UKOqlQPypVpQg5zswXX1WA
YtgSlWRymbwGAtxVp4JRhJfOnVjg1qXJiZQQ7W2RxlmDecmwjRgW2d/tUilb5lG6k8GDPClhNIph
1KNUmEFBPBHqjBS0wmGsTAH8DDoOELh4QbSzbkfGr3TNxNs/uvBbBbJzG+rFSvh542z1TcQQn91p
ZGHKHVQC5eQ31/BqhE7sMRzv7yXaP3GDmeucukZMQP1QIBi50NUOSiNrLvDQuIHoa9amGqb4qEbA
DK2Kb47FNJQz/G8Wcy1ua4Hdf3SLz8WtQ8PxaEo69WqE4176U5z23kpBqbElFfWOqqkYBfH6/PPM
WrIQ38j6Li3G4SrweJA5xsS1+ro1zsXNkTnHH+Oul0pdXcnFW6RpKbIq5Gpdx0GVG+d6DKV59/z2
uaz02NWdyrlKh2UETa45j8YsLvG0urvGqAn940K1v69CG4TdH/0durSEE7LC0kE4uKesWCoGgxq3
sUzxG40xiPLNZ8iv0EBDa3V8+VuhIxQzo/nYKNNb48k0ylxRMac290NhVNQTDygxjtNIEHcd5CqH
vW/k1omv5MGqWwpN+gYi1fV10c8HEaJg4HZ5g3IVg8tEp/z8EYqhlxC7JfaZ0EKfB0r4C3A4yLa7
7OHrN/8iOnQLTRfiVfPccE3xdgfde3D6oyu0pc7OFMgCEP/6GshGcmzeDbaLHYYRkkqS+4HlTbYW
BYcGR6mvduBQ3cth5zjvzP7UmZTBzgSNPgsomORKDxHjRpUM/AygFdSxtTxm8+zSTttjx/hMxgfA
NoWIafl0k+a3bk5dBd6CuiUWoJrUNVaQtd6LuE5C94YP24fGiZO157CQqroPYU0FX1TloNVcu7HZ
AT0gH4LU0Vu7l+Lh6rwj/OLBluE8BCqyu/9aVr4PFb84kmzetHR0W/uBwT6jix00kZaV7R9aFYjR
6BsXn4yYB4RXAVbObPIyaOGEVKnEZENv1lbDnX9YM++jn022/Ii3D/Ekq+LyiO6VhxQK0z25RwYn
L0x9XCN1tFTzq3zyk5mVH2uNTAkX7glEEuJE0TU3noKrCK8F+pCjDBmSivBGBptWEJZOZciUkXPr
b23O0HPA3Xw9WeDjx3Ly7faimswwrAFhAXGuhCWerJJ+pwDuqXafWW8EEG6onxcIJA10OSroTti9
7tmTgv3OUwFEbNLvNKMpGWInhdtqKsKnsGQNpibOgs7wT6OgpeIqUcWnyzzhecLsL/YXSmGjVZQI
PsbRHeDFC2NZnhRQWQpCSptXtC9CsV38Qc3rPC/E1e+NmMoLuOm+X3e5hn3XbY5WFgThfrrwnDoS
Z1OVcoPWTH1N7RmCaVXSX9+sn/Ky7SoiNn5SCCDgIQv26IcqrmRTOmLPSghN80//yrborcugf79s
SheRl4aeVBEQKnK0UW8RogCTHb+wg3QVxhOocxwtIT9FZs3VncBO/wNLl9NFXeClkItk2sCYoAB0
49We71Ay+pnmr9VHK4Dxw6u+3fgkh/UvlSn3Ecfq65uxBKSndN/+7wddFUcBKDRAeKpNeoyOTfpZ
gnlAZOI8CqJa+U8PccJZhLn7PNRT+x0tPHQGoK6SeAScY1V/6kbVepW0eXtvsuvpJ4MoF1KYIRf8
1oo5h3wdOukLIpQph6Y65ySCCnU5b67fIWcEZrcx0Sq2oJvvqfDJ73ANBtaGAJh7IUE7O4ZB+tX4
1gOhmsCQT37wOWrbfXdLbmI+sXYl9T/7PF7y6D1m0Gd9c/C3d1/VhtxUry5JYE3fhd6y01MVmOE8
9yJ8TLnmKxqD8DB1NjqXGDl6Hura48Yu3bKRFPgJtIAMlBzsN7b8r+ALlno1Kdod0BSMVRZlTEb4
fz4BHerACINXea7m+TP1ICmAyyCzRWaoCNynO9VV5AA/LE2axvYPjm1Ar/YxyrYLLBLnKxvwc5IB
u9fv1noAYikQdu+UHDI/74aY5YnYN4ErDMd8uud+oSC6h/2vl4RzhmnhjhB9U0sAU6xjRZXJGNCL
qmh9hn6/7W4R1UqF3a08avxNcEO8ZQY6iTDRl17ynZBBrF6Ayx8TzxZSQsqqfeLujuTAhpbCZK0j
QyN25SAtv3ntiMtjdc0m6Pq/9k1TQTau3VcWlPiRJ85gVz/s27A5iD52WpgLrHz72mB73lK6TTEZ
j1H8h2pGoyeYGuz4UMwIqDf3MRLQ5yr1aKqrSWJc9Xpmpld265B6pWLG7UzeBkEZgC4NtE8Cv9UG
V5vZ/oZm7cvOIX745JyRyayIjCaEHoZSM21fjcbNJzgtrNrYi2PBSe6PA460F75uUUndgElfCCLu
jA0Csb+cwaa3LZDfp2R03swnns+xFIAu5j2yhH//IqW0s9FU9TLV0PsXpPTUBNHzmB6ihpv3wU1L
nseyfNlHclwTlBR19IN4Pqjx8r4FORnZG7KvAIHoLlB7HUcQ/EXJTH5pJQW7dl6AkSV2irz4HgGs
0L8Z0Il6Pg8beQ4/8rVJdUa2ze/rPSQ1JU1eHH5FDTpWBHZp39rm1lFFJhLY/74XpstwXjl535G6
8Dsnp5pa0Gcr6jfwMe7vOsBOX1XwWnh+HpJILk+8/APPV8xgei2rYKlk4Kgi/o0nJnSC6v8wb7ZZ
JOByx43MNLsUP6OQkl8XgKU+WZY3jXz+2MrrZdIpGjJasXdtLEh/7Vz4ZVuacADGv7NeHUSaAq+P
Exyt+lj67hMnlC7gdyruoAp0+9aL7CDYwUlEuZbvR71Yz/NBCKgpUKc0+CRybmXBOgjD0AIiLvbL
MunJR6dRPcKau25XZtkCyFNx/Mlyc5CXbABB++AbipQXzqiIc8v91WwoOuumsqusOHNAEJNIAGLo
fCUO1SzIvN+4dCQz2ppzFHDOMpthsHUtSfwR52l3FHpg6Q6mOr3zkMvfWPBZ1gXkcS6FzjiZDAt7
674SQqKYRXRDq2RUVCDftHIRSwXfSrcozSP8XYpmrUJPE3TJE8FlslpYfAsUeW4mMcY6Us3HWK1j
iwlIziAtllADNPyUfs+4n0jaKFq1A2Od5fzZiOTbEtsqOHpzDu5dEQhMNuD6c/jPX7I5+aH/KNXP
Fn2WEMKFiQNqeG4odwU1A4PNubJLpI7AhzHEK3fy4LhrL50EUrohoPEDH9HvuGyVP87Rldt1QUmU
IyOeuSJvHJQKnKTWQZi+Fgwt7WuhyYe7hNXij8SRGYcM5QydTrfy/iS23QYPnPBGJCins78HrTdC
6xuNxuhK09ZtTu1CQpp9/1Yhp1grTuJt+2WdkN6lS8ODNJ55l1dptGmtqrrjS9tvVi4ifuJRnpxv
4Vs2i3wg2eEBvDxNVNQFZ5TYWfCeCCZKVhkPyc9zyy9agMVdHMIlGR3qbBE8CSpZwfg/KwKJ3ARv
Y6+3Mt1Cw7KdnzDyDStaC2o0bTo44E5BBWiq0YKGaxZb0vNLqPWY2hI7hFtdMNOwjpvj/jenkYOh
mW3E9AdmE8EJYqPDS8YHuuadCBnQnxHmaGaTu32q1jbmKpjizrI3Ue6Pp3vby3LZlmMXKwK3MiN3
e32AxA6XJOY4TZ+GqtlleofrrySKeTvWshOGcfpH4zizwIoODsZ3QsB5eHZgj8olSuruOuVO8Eu7
sz8EIADmrXTjjkgxMzz+oP5nzRqd8V+UAzoBgM/J6Gbm2tMhym43SIjZQsRnUEqSdtkEf3HLGwez
QHy5hcsHJE4lzHBS0zDqkVKYgxI3rli+2+Z55XdndP3+2LTlO3o44nkQaU9NacX+unsTDBHSe8JK
LedNxYy3LMo/RnvEcLkB8/XbBI89ziiTlN2DiVat8HRbzKQSzEZ4tFnCCwnjUMeHeLPQuIfx2+qe
O2EEynHkVR3LK4Oq3w4K1T+nZ821Vi/knXXUbslP4T5q/uAVMctzm9QJ7JcFhM89fY1DuStSGnFF
q+qSxPd87vwiI+Dc89slEloKtbwVTdVeW4kM+cIOg3NtW6EW5cl9KrHh1P2wzs1eF/2gJ+emm7k9
Hac1ARyBOoGQnkFotSYqaybpxolhTxQdki9UvJ0BvB+fw1O4PEa0WLcSTKCXXiymR0MfD3egGJ7g
WLBq7mGvZ3qx91xgMu1cZ20yxwSFVdUjKbOxZQQNC1NrR7ZoC3aLs250RU/g9bH5cEHWdV42/XTG
fNdOmjk/XQvAQybBepFlXp3aQ/W3xc7MiW+YMfU5pGBbjcd4isxASi9etD2UoupdxTw1zbv7lLYT
3XL2Ukmy36zJBPyV7x0OZ8V/6lLHmvn0wRMRtVoWb/quhJj2Y6JMTt/5nXbj5/bE4IMcLVxpgckG
KTZTMVJpi86fny5Evwcry4AePn+rXcgfbgxqu6OPm3TcMak8nmXVXArl28XaTIex6Aww/iZ24OCZ
QwJjAK+ioR9hRMeMm4KamWq6YWnrRXgqyN5mO+MOQQfsEByYjFhO1gtomWYt76zoX9s0DZnsEdqT
emgpXl46Rf3khT0eB5I1WH0uuckbDxxLcTO+3a0Pc1g30O+0QwJ1jI8M8NT5KFyWVVCdnJt7QkLT
HCOhtotPsiNFRwF0xqTlBaAU7KTIHotQ9OxWaIM4WmOTDEUgo7IXRW9bbI2J01YyVnw0B3rG5IIQ
kl5WNbtpXo598/E+swTBt2YrW/0bvOV7/jotdwB0nxbGgfmhnTuw15wSLv2HWdH0Plc9uVzQN3QE
a4i/Lr0SJphCiRkWZleoIMaD3sGfPNX8HQ3vOuTNs9v0GvTOk5DwHLXvxs8vMUlVbDOXDqB1h8oV
dYSGmrXNMO4Rgp5xXrdDatlKdvjC7s4hy1O3+82095s7t8J1sPhi8sIpr+eNsiCJxW6036XqUHZU
sf8aBW6wsT7+aq+S+ZKey3wHnkTiY7soMXBzMxWmj8rRrQ05LPu6bRvkv9Ii9c+C4S6UcfSGbfHH
Re9OhxbDAy02gQE29LsQPzRIrImwXMfCGbrX2CadWij0pAl/tCK1upKDqg8OS3LJHqJXJYQWKXE4
vP3wbQFfMDkV4gxfyvw+wF1W9WlHbdmudkFWuZy5KstauACoArn2CUHg2xZr3gjDPvU7IQsIVysO
oHOHNW23ifpPhjZvf/ra0a4/PBQLjTyG3h96prvrfjyS/TjEa5ZaetgY2z+Bk7z4vcJxYbyWLor+
7ALdzk4P6PNUdSBjB6ay+eColKEUIAe2Z6/s5pBtPQYz04Iemam/HC30+pYALxz3pkNX5zquR/fE
twsbr7H8/Wc0tpLT8+hXbgi+PJAlnSuDFRnm0N1yspkG4J+GnjXZ/4OiKgrkgl5uCf3S1yvfVbDL
J0PgP/O/akAoGUGnw7Bci5o+eq7JuCJ+zvZUYtf5n1JnZqZMVmQkA7oG04Wq99xkTKUoWpI0w55v
0yqC0hD43IFWBdtpWeqn4dCCPk2wdGZwVohv/3mAidIxFlxpEW0SgFpW3ZYtXahIxeRgbNe2dOyw
g+LBF6PRj11/O+jK7FHoY2OqCT3ffIq2vDMMwx3X52fHEOsdyCoNkH47ntuZPxhPV0kwV0aZpIsD
f1AGklwX1k0p05kl2LNFdDLr2PYdpTFrI3GyN1B5RWRk6VoQtJy/MwICyFybTT81icejnGnqCiJM
7U86TdyVe4ELDYTuC6S49dkndkFDzEKDaArHpFdYVfVuNp/OYoc4jkTRUeAUWUx/7oavtXcnvnnR
92mFWR85CIOcjdsRLx//fZ5rmm01BkR3y+mj0CD1J3SMl6fYtCowrZWhHVYvDoK9F/5riYiKy/H4
gsLDdVKvC2w3WN7XTyuWXlLACLsyE6+SMXze1v7DgOJlc184QIBdZrkV5BSqDx7yZuHFOA9yTmqw
8cp0HMV6/CV3aKB7QZHF0X4vsiZWFJ1NX6W8iXocGJuMDtgFSxO/oJcplJAwYHaqcGU8yvr4tm3z
1emNk2ms+uy1HAKM0fz0R2dMGdiNohqmEkn5idrIxwpQr+u5TNc2liO2j5rxOLcm0Z8JDLBImkgh
Wxs+cZ4X2vujs14ANubTWlyOk2uei/lsVq19+yF4B2vtPT0skoDbLKALiKqLS7BS7ISB6c2eC1Tg
DRFbf6Bw7tTHTjUNBKddwnHUJMcE2Moik5YCMmgFkF4dT+xUG7EsJuRIX3q7XKwqW5sOYmCkG0aA
w0cnIqLoYy52Yfhv6HbGUVeaoojZP6yl0kjuQQfvEXBqQW3EVtgisutFLWcsrTdvWIhZQ6RRLfVa
HK34T73OzjpXSEkW24sGznMTcG/iZrVlYELMQRDXAemGERxYr32hKfjoadGVKN6BRMIIb1PBHhl2
TDbUUVMbCbUhW4TMiiyWlN10wIrRO/MUpT0e0j+DGOtC0nxazt1QbZunkXeWjchGOI3hQ0xbgucf
LRMAKzaR860597Yn1yGudyX4w7d8hFTKY+jiS1COEbbrh6iZFqscZig24U/iZIlwPzwU9Pi4XUrc
8YEk7UoQhKKrbfX2cDs/lXiSpHApxOhD12zstu1U9BROpPLJuYCmPczstSKlccZLha+1/nb/quTo
WMAElVLbb/yguMpv96+dRe4OWu1yrlwx5jax6uv7fmTaW+lFCIf9oqQdsE7o7r8nNYfZM29xE1WR
5ri6lmRHAT4YAtX6aVrmpgr/DKkfrHEr/BirbLYEImTyqHQblSeVqxfYhZRrCT/EyQcGkUfMj8OY
w+sLNgAcaPDgojK4/RiXeqgdQD4RPoZjRzFFqnTC0+ibwpCCsZolQgBPC/BEsetUwQ3HkTaBLzSK
jwB2KnR8cwwCwzFeIg2jQnmhsG2l8+6kcbvFAtJnLcehGk+eOA7EaTBQBto6Rd19T+qIeSGkO5AV
6s0ot/o/5TLsFzP2x4OxAOGxa/YrZP2WMPx/9/P7aZycOMEjpdmbYO+qH36kWyJMt92F35245ARh
1XZk2JVeOnSYWFaLi7aG30ZH+1GyOttF6YXFkWx7kPsecMxX1sqjIEjmdGoEg3ClqXbNFd6ZzoS7
vmo0eIxEA4H6IuZqXwR6F5PpuMgI6UFtoC12zAWd1XBXrtczEekd8VtpcvssKLxaeJCfu5iFfJPj
c1mZK/RFIZri4z55H3MB6iCZdyXEfKjnhn4O4/OOIjN5LjXk4zV64N4X8MYKN76Nmr5M0mk14oPB
wUs8o5hoCS5T4hNFW1TAG/dWpLHrQl3F7zdRBd0UGUwpxCiHhDB9ya9wXoSSL4bmYoG4xHs9tqvB
wNxNe4c8GeWL5M/o5Os6I+qPonR0YGmqiVS110Kockt5I/qqSP3a+5fwO4MaTynRq18KfiOkXySC
WgEBkCBnPgYhnBQae6+5nL0npUJ+7Yur+WraTg2jDCoXT7rgGycZX/2aLjO+pxoZQuIYzyJ7SGDY
FmD9xGTmyM646sKLls0L5aLkmzFi2B6+pHSXICbAbjd7F/nzbIahkXurOBbS8jC/gNUoNk65f2WK
ruBF+J18qJEfG+fQUN5MCqVheMNte6Q3vv66H7SqbLgx7Y7QjR48sfflGpOmiSeDW/tColpU+3g1
rVMmc1QC5zAivyw40PSJXxFaWuwXM7Hun++lcA0xBHXFa1shlbnaz0wl38g1iyrTs0FEVyeCFl0p
3GEfbts1qFjxE0KD3ars+xA3zi0fEjR6rfkgANCW/9ZcyzRS4GveZrKjf/oEaWnC6n+3Xam/Twu/
ZHJv02Lq4QO9Ez2qW6n+D9TRN46q3LFrv5r2ockQFXYRWBxIPdJvx/vQJaq1SGq1xbyI2GmkhOtM
iORoZ/DJFjH3M5S/7ANjUt+C3QegK8bsDU3pYm588eqgFRaMDVSbgDTAH5ce7w+mHvUcQtHFmWoZ
Ec9dYz2+6aJQN2/thJ+rMO5QYrBP1qGH8hFVGO7tpaFRiOUWiIuxeGhLdfeIoDoVkGcvCp8zJ0Xt
Xs3DrjBcjo1ZxSWQQ7lOxJ98W8Ep5/qvwPhHFk0eAXeQjW2wdDvUTkHIb7gg51sOhIsQ+fN3CjeE
pp3CBFddQHeh3glwNJIGdqriv8TTvzLa0Cax5uYrpB4N9T0B1l9yKhWvqeGdqLTjLDIU8c9JMuAS
Q29uJjyu60IVxxND+z6tcoEqE8+UsySe2WD9ypMU+aKCjdfnlFepLrdD90A/bNEmMKb9aR+DYGKs
35gf/dZTrzl5Vvene3t9kFqViJUDdEK6hfW4/KOUyPVxA7jCAyEjFRXb3jjqOto3cNH0QI3l8lP2
7jvhlTb0EhYB2QqxK3+fjf+jk1IIFGskq9K8aO/kbBhzlV5ZUvr/gKkzndfjcPHnm0OFJonBZncA
1R5IWKy4fmQKOkkgL7+G1dyGJB+PTa+Op1rSX3Rlj0VzBaTSnE8kJoKDyzVTeFcWhX5dqJMixbgl
I03VC8bnKV3PKvbD5SS0SEas1rWyvzxEsxeo2C/Pl57rv5Ku5DKwYp4naZjYZaJpQxViLdYAlHxg
P/fX5xv5ozn2jwJYoSmp9/Ho8cumk82rsWeXFXjpSrJYMzkae3o9RvkGjOnD2i7hh7c6fN0bsf+v
5Z8hP7JG73QUyxvXxQuGbmawuxZSk2Fv2X87UZRtZ8uXB2oypK+5r+sHY8hoTCUxrW01BvgSZ9DV
m9AOzJPwp6NeJp3FSwShqV1r/GRBqyzlsWRALga/zbtxKGb0TVGIci3/5lHYKItj0IlHFRVIfH5K
4qMMHc1mrAJFakxkelMvKZ3UDwp6aANJ6QgYnU1WfAcN0LYm+4CR7MR4RZB/RcOkOr25MlcINqtN
Dnckv3UTwLZC+JBzbh24S5k7yUb7E3PjmPZ2uwrvKbU8xKEKgJnPsz5o6JyLC+s+cNm/XLt6Q7GJ
2TOSos3duHZklM16f83oEGL/4I1Sng71B72E9qAXQ+JYSrknjxwt4QBHBi9MJD41tLzX/3AD6+Rn
CCK6h4hIPi3Ecxp93VX6RP4/bkRFuVMqdfX5KzoipUZF+yTx4UuD4uEPjovED36bBtfvxExb75YB
cLesv/1fsLudOll0FBzjuinzX/1u3PQBA8o7qn5Cy7clq8y9OOke3Lof5tQ8W0BLoFbWYQRKVX2O
iHld6LDV31j9aBp2ZIcm0n3o39P+SWr3FzhD6i3wNKXt8DXMDka+uM1C3PL2zfd6Yq5Y3LH1ZFTc
fzy81/vZ8ZnKEqHqeVhfoGvEkFzhVk13L3uNGKzPZFfbFgEKbEpzgtWcINZkIytYeIDfoQ0P4U2T
dbCvXejXsrM2KWZkpHJQYHP7s0M2eQhscs2xy6VuY5Jam/pZa6SRVcTGdNZbRdDS2i6sqtuupkrl
wbh+S7T+YyS+XuyYdEc7E0Su2Qj3TQmfuyVFa/iIvbNoe1USnk19DGhn3fySqPIdZl/EN0X0SpD1
hT2FlzVnFT0CLguh9FD7hYbSLwkxF2PobP7WipBER8f3zkDfxHvx+kmOCDU2hjTGp64NwhPCoaJH
an0I1lrPBvfhXq4FkieLy46dyxySVAN87LkvrWIdaU322pOFD5MecX2VyNSlmrLtp9gUL8SIoiR6
/ijyVSl+wfQpB6CEXWL+WZG06R0RR9ySV9jf/VwpQO/KDU/YvuFkWQXQeE2z0SjaVfLm3XLUAu4D
tff03/l2k+NfXuojuFzj9brD5aIERMCbj1pHspmo3C51iWqNZP25mk5Ek+yVsYcHU9bHMrdzisQT
vNEANjKzYS2YsGDRHnyDTQRA2wGU361ZlkclmFrUhSnf5dfrHxhOzl5we5/DKVw7e+3HUrfxUpgx
dkiG39VJhNIpmFebC7Ds3YacqX1y/C+kAv0TPZcHgntuG9jnYaXIEjr9F03rOS1dnD/MlE2q6x1w
u1tksTQFzWU/7El4XKkXMJpxaDyaSb7vvdGcNDkj3Z4Ct4Mxy3tXMYDGeTDsPapE8nyXBzRURVee
s0pi56nuS2Fm3tLS00NhcSA+rq6wl+PEbpQiAqerVd+pP7g3em/DDhIR2NsWiSMa21XlboZ3f9OV
X+AsCL6TvRz2BgPtxQ9UVPI2fIVGTRznHk3XsHZo49Avckl2eSPZ++bPQAEM/n2bg8A/0X7ii/He
8o7mtjHeyesxxpeMQiyS5aNfoART+vETEGaBwZlnBYkKI0g2SaanwPL64J372+s8Uyfd2cxh/2Ic
0RijldbMzTBITS50n1zieDIUJLixjjdqGz7bVwn+OgywzzxxiO/AKK0BtaUfS9rGad+1+MiR034i
SZ7VnPnbZv6s50RZr9+JsPt+ZaYYZfj8BH36txathv+KA6gaAaL8NNBzW1tfAyGazm02LGCIqEDx
1EZDItLEDFy+tI/06KUvf2caiSO2QXJfUHdfzPcmDWSczwylc7CZaIkjdpQGv2JwqRj8SAHALpQv
PZNbIDk8ErUnRbc5XvGaD2zDn5TZ3efAlOxK4kmskjyaL1YqAdtXQiy2n1+eCwViyYpV489ximfm
4+PvuBhQZU7ZAJ/4B87pzo7tw6jSsO76xvUhpGyiS6+fj/pv9/Tf3tkoRZJyV1Xq3rjJM2QfoPUh
VBBqXxOEq73GTtZF3VhYq+j7hi8ixRi91sATI508lwkWr6BuI9CfkOID7yLLk4H/Y/clnPqOZvZb
xLAKcrMThhWxvtH/aJVY0ufeq1laxC/0hJuDdQNvTF3FYkY6ORYNcXWF2Z+J7l/iZPJFo/4JH8WW
MSU8A/6W5y9PazxrLxtd12CXJXv8SccKvRwXg/EiSHi4l8mSKNHvAnlH1WHK4VL7yb+u1fzCqzw+
AC72kodL/4j4UfCv+JggiNMdiL/cXeziEP7nFbb6cYBQzvMR7cSx3Wits50SgfbkwcuUSPwYrrWN
b7AICnsUIWEl3LPipjhtT1FNMFmeRO957yWLie7T9dKOQvSAAjpHEXeeqDKLCKmhrM3E/oIn8LTc
aw1keu5Qnay9Imr66AwZ+rudsTPqLDpDBc2iGwte5mx0Q6of+GMq2EKo+10AA7qSOChauhfCA1a4
2XALmzOVqVbit3Xd4H397IyHAi2vpKChDA+b/3/FpMVNImn48FfxSxJXOK/ZV+ekxYfxZ80fSZqd
sDIw5my89HPhh+eo6wfk5PoVhnlwrLVl0ef0EnsX78Y1A5cWggl2jD5EZJICkPGUnC71A/7+q/Np
J+PBetDCqopjtg16+HtgSQXZPl5UuIg1skFPz/Wymf/Rw7FCIsWwVqwaa8loT4YMUcTQOLOwE+Zx
lUPVJJqOAC5Jdjcb1mXXR+4ndT3NIkBBRNWjGHqbLKe0waSPu2yanFxhLzQjOEHXByJ8uA7PPdZy
+XdvKHceA8vkqAm0wha91yqVRJzp4Lpb86bOs9yUaQ9SPhFf8OSZadIWhmbZvjG1WVcK/y0+kPqc
f6do6lHgqko2yZ/1H6AQNL9F82VkvDa7lqGhsmNvtPQbnva4lMUGomdRLxnPNn9wALw1gKz8N37a
Dgjuzc0AHsrjY7hIZIvlRuwv8MZJmO3mgQvuka60HBSPe2rJffKhsWWt6Puon7K/Q3QF3QoFsbn+
mC5oVMGK+Yl/e+KE47jSdgZRojE0RB9Qvl0fv7gEZHwF62LOeyWJA3aEf2T8WuwaMqy4sgMSKUzn
Dp94qv2qHPfgwChqwLTtBU6uHHTvg6pyUIP+an/9cfWh4HzjYvdifRQe0G3eW9x5f9s7h/+UPRzV
ZxM38UJPPD/JsM2h9d/tBTYuiItb+OxHTlnLMq1KE3Eh9knYUMBh8BYTAAWocuBMjDZ3t3FgNphz
iVOW5NpHFSGxhR2hsiyfW6XH6M8lVICtnpEIJAVWCkUjBP3r6ZBa6Q47I9KFMarjwTZIU4GSeWP1
CCMIC8EzMp09UuXPh8JwdUoOkwH8V53ddX/G6DAKs9hkGGepNrbJ4qaVGy1qEQk8cgLOb0l/HKZu
f2fNQcadBH5IwoKzKPyO+XjwhAvdC70BTx8Zn+yGDJLwnD5z/oK+d8kT4is4xSvXP1T7MufIZ7J8
LmXcHdp9M92g5oTdTqo9mJeIZrjyvE8iQXsre8K4bXvl3l8HZ3ksM1U0qA5rxAGyu0FpOArlg43S
icZaC5YJgd0ku/mNrDW2bKPMdDCX9cVUzO//SmrDJ9bOCF7qCI7CJgvSpWtbG80j4fFPag3E+xtt
qA7rJrIYjARGReqEykWHScKxSII+FH3lDJ+tnHJ967xFRsz5dz8kEmH6mBWnfUfXFpZmzmjLxypg
W5NdW94EM+eGxFYD1oqjook44+s0mSStrIniH9l11drehVrXSy6Z82hbJ73LsP3crvVquK/LuKCd
RCtNmYMTRfBonl3bjciwnD0FkQ7IRpBhL7lMmUZ/B3tNZckNyweJTF2ALHB+wt/F0WJfEMlyvJkw
oS9nclqw6l+6gNLQhsWAEnEyPPpAs20Hk23StPG+Tey4/9zfcrXw4uPCu8ThUyRGbTjj7wdR2pnG
UXx4y2hYHKAfqNhfglPlHReTKA9hEwKp/lEWk8VoaUHtaqxflM82/+VLrVQAAIQAZNjdotQaLBO+
Im00FKfmXxxF23HisBdDGmlOepydm5NIzjhtXTMLiVFEt3Yszb0TYnX8ClZm3jQRD3bh/wqXRzVM
wBsDErHZwT1wLWV6zvPaZfQ3mEWzilY1iaWgRInVYI5fh3jMIz4z10FcuV3oxKizGKiQV6MdHFHj
u1JG2+vGx7oe3lRypvKe4IHmAR7H+rxYLBMWEB1AYv9iJrQqFZ6g3u9hDNgn4ud3WGYFce7A2U1q
6ezT/nS/50qgzefiaWCQWjhhRBWMAOkplaqQqwdKAvrtUfQcbDrnkQX5R5u2T/VfU9LjPBT5JBf6
XGyGfG5RqEBVKCPdPwAEuYUcLjluRh2U9dcOcGikWlYPXUoquvV/TqRtMa+DDiLUTndebMHaM8xH
019LgY6fHflrzt4PTZJ3HicRqvSiT6JuCCEc8iErcdPd/RbPlcaIbv3xEn41sDqWtgo/rx4fc3j9
qUv/ymzwh6DRbaO26pKRcdz73cfIw2V7QHUNSouFfVH4KfK4foNBr1/qpIN1NeR0M3yuLps5UyfT
e0D4cdWSu8U9LPAzK60awru+sj6c7Ls2uvWiRq5fEvax9SNlFGc1KgFw9AzT7ZkdaAe2ZZ6pbvpy
bAPR1tOeWyUBEova5X20MQxPuwNrp9qwBu85W744YWevYuRADWYlLLG0n9cOY4TeWcpwrqlAqPPy
rp6LUyGLLXhE7Bl34wDwZDyHH3NsbJvyDM/ORnVEy2uf1c4mHS/OENV2q3l4dTaBGcMfpqavgo93
B/QN0GhFoWabNJQWOiSnhxHz9qQGLvuR4qAQfpK4mSv421P2fCNLAIN4PGIuTEYBk0R2hXudvVe4
VBmK4BJ/LsMHtUNoAJzbRxccAgxsnfOmzeRwTP2/IAIbKV8n5h9o98h9lGgAg9YgQHp5DaTSVclT
QU24KhhcdGkzvKLMYneX41GV3iwl4+vR5EfZH6hCfI44yjiX68wbYvpLWJMyGnp3l2aRleLyrL1U
tH58INSQr24U3WbAAKVtfPHsgjDHx3grJElknNZt4Flpoj4egMKcRq5eH05/cmZSnXMHBrJIMoSn
23VEpazo+ytSuWK7UGNKME6y9q5a6EMb3xidRbMSQTBcLfaoOr3u5yNGgaS6qxF5Z9yaXzSyq9SM
i2qHepB8pMclkyTixiFGeDuPqlgrGZA/J7XNaf4meU9U9rxFOQqF0Jl1octoLdOt6GnpSQi2l+WW
x7nuxfAsdu+EidDqLDvw8SsxTyu9apfHnMDVdkO6ufPSWippICgwfeHHkeeTVngdS+F/2ZdX2bO4
QZMSLod9zEfNlJE3Hqby762Q3RBCbZlLziDg+I6wqypNNwi7TAahJZimbavqDYO1F/cCltggl8IX
8G1B9kfXbYogcxwLR+ajege4X7ZIqqaCy/Y23zHNGyMnSQQxyUa9uaF+vsd1vv/qYfvLhHcNIxr8
0XQMXXDHjv2Tu/3jJjYFQQ16P93OarVJhggtOPUPSHbk79Nn46V8fvbOA5GyXT3KBwOEBznG3fmY
SQK5cWcgota/T3Fkad8SY5+0oiL2QSow0BH/gyEhYfSf34AARrZ/MQjwB9WA2NqfDp5x8QSZof9O
lgiOKQlwX3bJNY/OEYx1VSigEQ4OdaEWbhM8ZAUXGb3/m8abiqQ1DYI1yFpy0B4Qe3UasBRorxb/
gvRoLBD2pL3Yn2/9phEQeYwnF19HHHVYFDt9I0DoHf+5jn7sQIcYHuXE1gH5ArwRrm8S0dlwUyHi
g+TStNLNx0cK61vVEtuRxy42tvCvMvrxFYVXwYSeyeD0XLRGB9lJXJYZ8Xnq6n/Y6a2G94Xuv1sQ
XBo7OoQdblVjFNQpz1QlL82zzOhwGspY7zKhWIUYpanF892elbj2qvN1QRs11GhwVIyDVY0z9P5U
RG178Qyw5kAjH4lOoy85ZEDiJCHRbdbMBIrx/uMoH/GZoWKqHIXpzMnl164HRp50kuEjkJDpRfUa
9bR+loLA+CT7B7/1w/nxQezlt6Wcc2BcWLEH/VEvXcdSQmiOpRelL6m8LQsyZYxT01wD7ueNwwhq
PzKkGeLjQB9mIF4/4mCENx+oBYMXFJoHeYPMWtNKryW1NH4sQjGINF3wLUQ3s/6Jq+9n2kX0DSBc
t8N4QEvB9Wj0WqG4z47N03txoqmewaZEhbJstPXzRXy+P+cQfLoIPu3hZzVx7xju0SLiu4ZA8MEj
KVfv9o0A60O8wrND/LxK6Tlqs76CustzuvABFaC+JlEeQdRkZBeboUsZ7Du1r3EIUJNgQ2barafq
h8OW7g+SnuDTtXFM3iuOWPzoy8oKxp8ynyP5ikQlIg6VJoXV14LxfrBWP9iDeB8tm/XvQR9Me+jF
4elMggjX+g8R+DgBQIwM4LwmNjZeZCqjD03cIJ4Hd3ZF+wduwxMT9vAVWphCoI5T1hdKD5pepHRu
spd/9erFVtOMqv/32crmf6ZPL1twEZ8pA91P0HNTBYmRqiul7kccvz5leRHDsvzeXUZhPlgj+L0w
d/G9Pyg9pyeHTCJCCblDF6vd7X1Tb4s2lHN2XE5QlLha8vmzRSJSP5X3zEg5k5WobiqZ79/SEMvT
56F13p0n1EVoNajYmNNMCm6lCBSK4w5VLVQO9haIe1TQtVvTDEOew46mmxJjQDLLKB+8XNvYrao5
5Qj/w0HtasT0cdZzARJ1jd/FsPvyZOpt3d1qnIrQVIGc0UVMfTxCBe7aXBKuNAegJHCC7jNj1f+i
U4eiBOvAXZR6FsiZgPVAHm+l+usVF5t1YWzhgNshvJINwLOoHJw0M5LgJhTTfKQyryJt2gjKfYnS
YMtXotK/083tG6O13+q8bT6X+rdd5+DYYY2eRI9/r9bjeBQSeCzAn+Mt8CFviTKe9QZacAx2+P/T
9unhtnH+H+I4SGYY6VCWXtsMmypk480bIcRQ6H3GUi3r5QObyk3aGfpvhn0bPAQaccnxKjBrBPqu
dnz8B+i3stSzgDkkmc+27hPPZGYtY2j3tzSC1vjZYGjLzgwFn91vuvBGtm3LJOk7x1YqfI8dF4ct
GkXgfU9k3iw5dzOdDGKtoLrsFN3gIsYOWcmgyACR4o3i8k/QH2QYIgjXxdq8YNMf1j/T4COziTHr
kQ5Yevt4+gdeS45SndnO7lLdqBe4PUKMM7aV8z1EsDhYouFy8I1sAtbG0V0+TygsniTSUXIVo/O8
ZzLcCIHA97Ap9UPsIjRcPIAaBfr/TSH0TlOsJsla7J7SIgDuSYN8xupmPa4j6di2lJgNkgoCEpYe
7apBp00ELvkmK/LwGFgFxR+WErlQRjRbtmDnpJfz/Z225u2JptkLcF3aqDkXxn9loQS5XEcg8ZAc
EDhujPzk13yigkP5Ox0XzciLtv+LSJu798JLxTKccpq6+a870EX72sWLWolTjjokuB99+taOHPfk
/zIIb2Siox0l2jGITxSbhCmcWij8FJyxYgSw93Y4r3fAwycLE3ayS9StP7XJpOxquFi3UiiLwxfE
bmV68YrD2QOSdIgteg6gEVPGE5hqLzpJgl9clys2Ld0k/9AvyIbtM5FTKq1F8s/TPfEF8S/8legG
LUucFS5rFSE9uy4K0VkRmzz9SYfCkoreFDlus99cahxF7sTPBg+DVwIOWgVB7P8MoeS9SVRmcQQo
F1JTQFBT+wf1aG4+Y44Eow/zlMBWIkmncq+wQNCQT4xcIOpxPWEp4KWNloE3dcB+XbezvQCU3SJQ
ieQJqp987Rn3itdZc6hmnSkEvBxtq2bQFbvf+ef8mOjwOvE8reyjht7kFr2lyANGxM5CkiTwtAYC
ePlo5bZSSbgTVSOMwExRjxHulQjYok8LnCUKTzStl+1cA+zVFIChsx6IPacLUxX/2y9SmBLsMlIc
42Gj22DebwyPN71ZAqiLETlM6nhq4YYYLzxhbvvzCZ7IpR0gU8bQdXfK1TukYHSSEerc4XIpM2W4
Agnx341G5pOuUdMCDx029Obkjqdx5p/CW3aqK2X9k/vDFR3Qvv636okKfnMk7dpLVJ2hCcTFeDoe
DhoZJwdXtRQZMJyOSDaGdutBY4+Ggmnr89LoQmJzVLeKlO8dxOyK6hSeto1lCnSV8CM6opULfH88
4k+Y0CnmXJ3/HSC3+j/9p060r1TImsHRsJUIm3h6gMcEKO3B1L5zLCydzTGPIT1zBhDPBUWjvo1k
SN8hRuWH3ip+A2OqmBUypz3o+/b+zCTUrbpXGOy+pag0Buao2/JQMda/GnVqhAIY4bS0S5qQ3+bk
tiQBdbVcb94rpSkNDO+52ugAZCtjVd7oVscKHxih5g9sAdX182H/99jb8JCO8dNS7sgAR9Q1zHq1
xVDYEwU+keTvVAnyFKXBRQgotZrLgg2zkU9aq6+f+qslK7Zuv90elQZNmOoNTtd/folci/LpY8/F
aTl+cEnevf7kLYwNp+8HwLubGh+W0N78OqMrBcIM3ARLXtTlFdmXTwTkeIJ+tOryUS60kpBngmt3
/TIPexF6rMVCbXeZ1+wzKQu6IYMW5LCEYWOMVvKfc87+HpuHQsYsfQ/IV+HhswKhNykmud5Xd48a
HVvywtzOPiVBJEHLmhoKcchNsjnQ4cwCl1T9XYNxkMB1wzmqBgEDRDyW7iPrtt2+3XMoZfUzLs8K
cTcnYniFmJV52INTgby6L5rPoZLtbIlRrmvly4yoeiumrUYXHqGBiq3BzEdE2Xc8eF9w7M9BrCS3
rjwsMwppS3SAGjy+u5qAoagMOHN0myT01iLXQSM8cax2IoxKqh+bSoIC4jvlu+p5uB9+oYVjQilO
zw/V9xLS/FNO93Ra5b5mTGofa400dIFqN9gfXcJfVgZCTDPwRMvBytXSxcNqVGf6t7m08NOdHMwk
jDh/N8uFKYgkQqRsiXxNgLhjsF5Q4XVxtT755oSOYrxjH/etroSqtUdudgSZ6W5118ecpSs51FBr
UlktSnbGEwahYuXpkRYmlzFZPw83M7Bk2X2QZJO3NeufR+sIFQyiPFLpLciaCMLv1nweZd/ki00h
86Xzt899Y7MTgCWuBdqmlERAvjgk6ZL3cF7lNsh5QJIMdUlGt9w4CoPBCTWcTORZDGV7QNy5+Neb
kNvWr9fGFe4Nua8ZqXC/ngXoPNV/xynUtxhTffF8hKQ/1rD9Ql7oPButzpkhew1uIf/9TmVGPmao
K1mVAxu+ytW5MniDM+GYkUEzrPdSi0H6oPoR+9UuRrNO8/We/ZSH4bxTtvEIndjApUQrZAtutQGk
+YkwU2uRKjMygtEmleNtr7WEZEgalm/YHPKu9P++jM98jxiK2oMym7gOIdOtpWWNK7jn7Lypdy8Z
DbIa577OSgrj72B/ZnNgAeMMaOz4BN8JiATNLwFWMyhBncdFbF5Ug0EFbxNJQeCXA0amcna5zVHs
Yqn8+jMovzWuOamDrsLeTqM9Iox8Uvgg8vb01Glh/ZIHQUlvdTv7dyF3l/gT7HagWJBU7TZ/LGc3
h62R0CHZJ9wnAS/t3+rApP65sZLVK0BQeWUY+JE27tRrC9FBxtzSH868HEUFZ6Jt75hKh7qTdPI2
R2UCJpAKDXlx3B3Q1oFSO33MPvXbBq0Pw7c1ENnQygPtht3LlVdlKnyhpxtbXRUyOaTAO9k46P3+
OydaEHyZCzaT2J+McrA5vo1jVfAzTBdS+Jwigr1szdivblj6CsOOK/ngzp4/+orH9ByZKj5fx9/b
czdn9fe+PkfsXWywn4rp07qTfFTrr4sdioav9tSkP5rPtt8NZNXU4ta2FsXE1VFwOklGrgFjc3OA
kIL3Eu0UPbyOgmJrXqRc03SLalj3xmca1Nvaqm57OIW80N35ag1MNhGE4am0tY/Fm6iZx+nWD6DW
Hk/DvZMCjJiqVE2Ws3JEhb9UC+C2Ihu6hVLB4rUDKEgTv3wJmNaJfIrwxT0QWCfY9KYtV9CxuyVB
x0b0UzkU3Idn6OWjzZDBlQxPA/L6Pa6zqb9cnhYDufclh+EN2gQwcMJ7vMPeqtFdL5aln35YYwG2
GOF7+81J2WALx+qcVr1P3qIe79JQUO7EjxH3UGIRQ8MY+xahZ3qKTAKnnhxZr5Npx8A+0rnYpmqL
fS+4amnYAx1TOR78rVfvS1WZEwZu2BRQoZtRwKH6K+KSfu0oNgWL8bFZ8wT/lMUp16OHhR7RyHxk
IDkneTBFmxZfrJInbpxG+GogDFTG8359228nZdydvFn8ft3Tc7ATUpd0r+phd6wZUX73B1nPuKSQ
Tagh/5QYJaKPavF0QFFGFc6qFrr4+kS8CRBwNc+6Tu9txsIcyTS+ltFLpi+TdQUygGGoyDhyLgE6
NUTGjukNB37cbNTygNXrmuAWuI8njHd662pLNJkl/ZxbSehY0dVbJH2Pq5g55REvlb/clAB27C5T
ey3VoZnErQa51y4pbRANIEyGv3F5dbRGw+OBvX6iuDKcjD8y9zCLRphPDBHbmNA3P1KbNW9vE7vC
SgUlL9slGf1jJRSoqESMmwv5YpCcjF2lETfoi4dLDoMNkQhBKRpYv0Tbrtyjp/OzlOpkLpPSA3L7
DHGsf1hf71tjwVFGMvMkr0WIbSCIMbex5snsUHpqpTATQDsLQW2XVlWCUFTnegYU3sOJ8NuCiXL8
P4lo8M+dxEuxO52nKS+he6V2naOFRxuP8VdHmbO6/xaFdV3Flkouc6JZ1FWwalQEkmjXtsBPuGJc
+P9M29OfvqENpD7Szlg2UOlz05FQmrJzuzyGjG1gZJXh3Cqo/c4PcKGypGuD9H0SQX/f+5iucIek
6qmZlpPXSZDJm33L92henVXPDvgGSMh71uxK1bO7MuAdiL0LnXUBCVw9iTre6kIDEme/SNLGBoWH
ZrdB7KM2isEVFYtCGnhcp85S3x3PMjFF4+dnxi0tbE/vPQvp2G7qRb1x3BII1rRqgfqLQBfSFXqa
kM9EEJWB2KwA08hqnlEex9ooKXEw8EjAtjob7Z4n2tnx+CMSvvR3Ulm8zM8A4OgGSn95i2dkcC8n
Xu1lbRMh1ZqAII78DXsDTht1YDZ8BKyjG09dTuW3z2hF9eJK0lBv196M+rdjDIMrZ6KBbqb5RuRN
kKOY5fBVdTfHRJX1X9wKInpAUdRJJ17oFHohTPTDJye8oAyo/HBjozYwzOshrSKwNBw2k70I08Wo
+/pEsR0vAXauzAuIr+NDyDpP+qYnFwzlQLhdAQsFEJpwpeHpXgnqBgUNkB0mzQ/ZxwAYpsg/koJd
UnHsnoYMHSkSjtfcZEyr+nCHutbImn+mokX1RepCdijczkpGn6Ct4aiWHhw4eQ30brYxzUBD2ZxA
qYHjVAzdXw+M61tQoWBWhm2JcSY/7jVMQrb0rgT8R/E6sZme3CLeSA32SrKzf2xFPRgajXVa00Kj
YrECg5aftC79k6az8XKacCGeP1rhxcR8aVAlzzlcdUvEjDbShS/EFkSEdpZ9CpxS8f/di5G2B9kB
lAB990YiwYo9RMcCR4SgJbWkHTtMoXQ8TRp8Q333VehzZpuCCCe2Zg0+VQdDervcKA/dh4vwe5dn
f3C4Rus0J9Llxw8vZfEObplKqD0uFgUPZo4jw/PVeSxuXwtkLbdhesCW7vHnHC5uGNUoy22EKF1D
PaMBg0j591F82zA4J7vfvWDUJk1jpPRP5NsPKjbvhN8HT11yjaUtoNwlZ+/ixWocshGMxAlyyNPm
ePt1H82Jb8trH/+MBMcGOL1SeKUMgon3lT0xJdo5q/z9SB63ST2q9Ki9Mrv27wVvdrtWdUpMSfA+
sAxBEtwcJdvdAZkZWAfQs8kCf+qJP0g7SKeQR7Ettta5xrlF1bVO0/7EV75TIbo575ZOOK45z1wx
n7UhbiKPQqpCSlZqfbsdhp0v6pfd1kQ6NpVtp3Qbp7Y+4ojILH1XNNlHVY9LEfZfPMj5bgN84SbS
RHivTbRoe/+ZLigNVlCkipoHxB9ZRmC9M03KVvrloEAUYAQqMUfFDgTONnzigL+Dj+StcFGhp2T/
AvILqfBvRIWmYp3cKPHxZorabZx6rneg1kUrLsy2d0XYPlRcV/DcdfRIoD63ERAUdi01w6yoshn6
fUMZ6MAj/Uw2TTFyH7hjq8dOD/X586QrMaX9IvrP4FOvJbPipxoVpSOVRY/D3v5C2dTbg22J0OjN
ADZ8zj3Mqg+khVoLCFky0sac6yIVe2nH/xGqoHGue1SCu5TOWPQ12cB+YYqPtG6njcwIR2GhxevZ
hpdK6M4PHG1bCWcdgnbhlB0TFSyl8g6a7OXMO6z8yEZWQFkUdwslzvTV5nHPUHtfRVCwKED49pIm
lWtaOX3v/jLNSncF05TOzlzlDap9CVNx6C2LRyunbF7jedCLUa9feuhTla35fRcPb2y7qxFJfSSP
k2DBBlwPowkvozHQiUEIIS3FdvzFECFxZMk6MV1lUmejX6Dlg/6QR5Lwe0EmnJ4Ze7GSTvo7JE5w
dFJi1WHsoXd7WxLvw+6fZCD1/U5P7gNmwTnDYlGpXOaSo112MZA89HeRrM4OFVTzyZ3KSePgikyk
XH3/swiGyfs2YuZi8caEu/1Ley4Y6/LSXOzCT6BL9rgl+vyLQODhemoaNFhb2J5jFhmRfbVHAFqu
RXMcnWDLT7YtCfgzrf1GwTdRGELCDsSx9CE4ISu0c+FWVJU0uSNJAXqY/6kxszbTj39c97uZ408Y
xiQxpg0c/KN1ixSOPg9xAlbH6CZAbpKRyPokd8Uz/FdQlTbN7hKqyh6zqOPXCDCCsu2GzsNlmf6E
ufgYjxxrRleXkw8wDVh/Tt0rXKtDfKEYsiwEZm2QKuG0khi5nUi5+vnrDBuTRTqCPVHSaO2QUz98
SlVeazZ8N/RUDf4ca/nd8k9gCXHXW62xqToUf23DODjVCLzqYlEko6zZnIFuHN0rGP2NcfoTG/qM
jB42LHMQI9WNUcwGRv5C7CqG9tDU0ii6ttjH909+veUkWxxghbQeHofaf8dLwB9LcWInF26yF5+f
lMd3nUy+VH3SRB3D4YIHv9x6EVxdWeImsiVYO3nJWXu9kILG2ap0Ht2kI7TSSYhW6WNwL1zq6c/1
CZDCtBlTbp2nGYaB2ZG3zBP9FLZelA0qpjLCJZizn949OfxYakbE/2N1yqotllF7yI4sprYO5+Tu
/TCvd+Z/i5rrlui9It6M6pcsqRIK+Buvht5pILJaXGTHGjFS8cB3szPdQjKHNgerPlXuvOQx7I30
Ksr6j2GOve05uIAmIXcrHJ3idZybxEIuc3LmImkb+Su5gJ0TYuXqZF+pjEa6JcJmz4mbAUh39x4T
PNUF7+WO9UsOzIozQzMacPrLLp+yM8WaMn/D6lYIlO/KU0ZRgzxCZFRl/r86j9QXlx3imhYgp2uN
U/i3HEjbCIOmm9c2QxbQ+Pnvi/xfOORpM2Y2CnyRW6Wqc5WFZRptW4Fi8jEn/28OiYqDMgGCAMNm
6RRthG96XrMdwe4IYoKumNFu0FJWAeZS8tu3oR04dHQwx7EMBFeDUWiZ0nmhwjb8vf2W97MS9GV1
y6i0gkvQR3lSfijwHsADvgD0TLxlrKDyZWrhVjSaWr1KTTTz4cEUG0DCHGKGUI8zNGO77D7HKt0r
S+TWLAWQ8WSUgAeuTUPpzprWg9xLWbR7AwI/2/uia1LscLfiU2HSUV2Kbwnp0Cejc67gyi9cv3ZW
BVju2wmWMLa6bdV/LGPtrLkFxXqwogzIoZbCDqK3lsDcdHB8kbqsqNTPNIdbUGeWdcnhnY8e5sYC
tefWZPMaZPb922zmd2eiRpAGcL00PSC7D08483IlmhHmiTSmR3HbDq7+Ys9RwkHRhq9s1vsKvg1O
d/tTB9+kyQh/M/AGJsXCthJhaSttrbln8UT8vhzCX3Aj9z6nUaVe9GKYL2VvQ/oF/K2oN4q8Pyzj
+0DkpEpHKgHN7VxpW4mN1gqToDcm9wahu3QF3E5dQk1ZuG+9xe4AOM7ZMjhzX/9R8tCNQaIwUWxJ
njqFv6ud43TZTVx8VLbjexMy8p8dbHHYxfevTw10h1aqvH+poDskymPwWkEaUBrVZtCbuQ5e9gOx
lgLUk+fXHWUlZu9Rl/ajcNYtoqpvH3e/yF7ZMqP9JHM1p623pPL7zNqKoEigJhRLE2dq+Qrc4+nj
UTIGPGz3oLPUmvTEasLx2HXsRQTRoWnx65vVbR5q1X0VhSybl5doxSmkolms/HfKTabxzCqHUEdP
l8O8VyXoX/ZWcDyMCqmfGUcZfjVQgJTt5fz29HZ+XBqufP3BD+eYnXaVDMf9aifVm4Q8sjsiVrhc
ifFwvVfD6MDJTJ9WwwU5xrYDrJLEENjjAS5C+ulERn0bno5/N3LVGLAX6VeM21pX9TyEDWzpMK2G
2XZovbi99lhJ/BBvBIb2RbEyn7E05F/fKn6Omq82Qp7JmNLJ5byi8Epp7MSJF7H5low5zNEW7dj+
K6/PIvxoRyYdMkBP2dpGSpsOJiDDzCxr5MImmt/JH84CwOlf6j3o1XyfDnm/b5cITpzjUwpJFElH
BEGHIpk8/ZzLa1GdabLV6R1D8I1gdL0QJcXKRwc52cKIPzQ3l6TVx4VLCHTfe+cQKso/6Sdqdpby
+IrqnQQ9HI2VsBgTNjmlcc5BtWFDk5jjqUt4r1dlWYn2Xd0zcKo1XiXSRVocN0dcsUZXkxhyoegD
0ZxUs6jPcAmvNgXjQwUFfl9NN/+d7j932mN2n+FgYOpDB73LtNJ337u/XGu60va4rh8G45ee1WZa
P26dD+oGpOMJQiL4xNFWoXBiDn43g9Ro8V1fLinKsfpqToO9VbGoaY0jhCydxJZ/OiEG0DYv7cKd
/s9xxctOCzYEdhSHH42GLBk74B1VE0/I4aCkwynBvWyHY1B2oxbQWixBHvhpJjsZI+6Z8rRsjEU9
moMX7vp9JPLMAP8EplBFpBoKtPGai6QfoYePYkyyA/fiYyTqza0iStbR/JfzhogBJjwMQnYcBk67
p1qlz7mVdImQ4x8u1BxavWkq52ecxqd9UhG85j7F8byaJNER5pz4vkNm9MxrPcP073P1XFPjSAIW
h0We0iHEAIwJyZJAwFfHJ5QG21zeMBFVpdiYFNeCuVIVPmKtrI37O9xW+FY9oYbYEf/OfCaebsb1
flD66VzWKsQ2iGzVxr1BSXr2n9YAAlsZmpLBJN2LphipYHoYbeer9p3Gqt92mGN+deYGNX+QYR97
Wm1Zn0Q3rXDw7h0G2vJg8jtrzR02pCWGCKnTcs2a2A7rXTokJU7sp1dksh+AOSa6KOhHcDMzJp8g
QZnSi7TEywyBtdFKuAah33Lns24hpxHvbMpaP0I1nRKBHxtNOHXgtO+j8bcH7Dwl4U5FCJjjfbKr
2w9Qw+DVetxUmtftZyp7vX5z8t9xx/+FXZDrNYFzoFKM9GpNOx+JLGtxJJ5fNu92tafV2IeOhj7a
6R15NZPH/uycdhU9Ldk45hGel+bwhLM6tM73Gg+j37hqjyYB4sgUmYaY2/u8MYL3Xlg8SLrRY0KD
8oog3vRtdR+hUwMfoE3OYv6StIZgDMbWkyRwFi64O5nV6EDuB8MlXexgCHQ8R2FL2RBuO+/EDhZM
v9FVMV1PPhU3incP9JjIm3lZRcw4I2mh/NszT5SOkzL/XVHVtMWDF1r3pzkOWeaw9dssn6TiTB6u
PtX9bUyjckzUbLhrsnqi2+RAvaopgaxeE7toF5SOKE6KoiR/tna7ENlBN6LxTLQ+suP3+TEpGM4v
n7+oUUFCsMFJqGTmjfbTzOQrKraibe9fbyv1Z4vlm1DE99BpvaiITNEoFg1ipv+c5bs2giB3B0dD
S3OxLwnJKz6xeNlt4ybcKsGJ4MER4aJT2nTD9xcppleh3tyzZJNHZ/imI5A16ZgYRQ6Q/hnND9mi
yDb919pYpGi9D0A2X6Tzckx5r0wS6mq+WNJ/711pAKa4kbb68h7NdvJLu80J+PPGiOTHafFIs1qu
KDgmsGeqZb5fQdy93KKyOeWHR3rLhY4D/wez6lzeZpuA9ziIW4E0e98vNdfFCbLHi20yKQrwxZxX
qrNLOORZ5diHBDedrzU2SIa9jlkMFidHr78KGbfO4Do13fz5uD45TyP9pMd9HBV54kycffIoA94i
EWNrd1Au/K1vpUmygM4by0r+6Pwm6eW8y+m3NM127iUJ4YFhWHJzDyuTOgcQ0rCTJeeEAjErvrtx
1AvIUur2ZJf/yFhsVljxXVXzyo9x5FP0P9fA1FCRMbZzChnz52fxhrMZhrvMKoRww1Fv5SRupEuI
5haGPBZSOKO8TF+dKEQD0TPFRJdeLLrWYDwbYkUUp2XKKP/eZZ924IKORYBRtOw0hIEXP/KzGa1o
48jafUDCnTEPK4Zc6Aa4XFqR3SsvW55bMXtQ5BoFFhDOX1/m4trq8mzCbkqwhdFZ+e6Tb3Ul8vZ0
HAxqM77zyBYuuG1HM/WCduxe2TkAb6AnkFl7lsB8N8OWM4Y0Z6augO4UzLG1xNcAdkuGeK2O0IEH
7oWIOr+g44PuYiBaNzcqKH0FTdqPzvGkTdZ0E5SnBBgsbB34Du3rIgr8mT2iQ18KG0yZe5cfgFdo
jzwFLTTmPcg+TGCIMKCip68d3PovNRAxWsqH2kHW6dDJ303CsvYRh98HQGV3yUwPbW2qHqVoJ3Tz
8hCYyMJmt2m9EocMK9tpQv4Y4CgcwEA2ucUPw/f5L6IgkNI1cEmfBO0Sv/viGVwI7cIm7ciX4Il/
Ka5Gf/H04hRdlmkwe4PnZCMU19kxJTmJ9amd90pwDDEN15LOgkOshJ6jsmjKO7q4K0dJPTUyi5BP
kyoMcLknJbNhBU/ABoe1yRwcG1TasqF0aStJDP9DAlnxGBQxugbd3pRiGBXov9Rw9bQBr35Y4+yW
Qju9bwY80l1Md30YR2K+1YthOd9jhapXuvKcAfLFXaI9jjQmJK5mxx5D3q5w71/+JIlDDQ9YhMcd
tagtJFOZnrtoyrq8DRmhH+RSneBybuICi4MAfila2BpeyXJalymCYqvXlIvDlGsSqCAHryCHaTlp
ucgz7xXvplztJUbPsBCv2BAMkbT4cpTBH4xLuZkKCJI2ECz0cVL7PHy4fDagu0lDU1D3pVoz5NGv
fGlZFpiCfJhCTGB+IPe7jcZMF+qdwvP8BTyfcJLVIA8Q/l3jyVNZvgiCO7UU7D40ic4MfB+tDbRO
HqTRYna7n0JbSSf81ibBGvpRnHt9Aj4lX/28aGSztT3XPI+NSDAwcvdXbLmXez40oFNxXJXRhlnq
E/iuOEe05tqIj/wIBGmBMtjQMzo63qj8PHOEcQKHjfqdoKhP9pj6U8TnkV361hSj8qgsYAzNr24q
q/6rPxGC5F1Q3tHO0cApo2CrcKWn5E8ozvQykUChwOkQl7DjPUh6xbn0kr6k0X6hnNp5+Q5PKits
LGIJLbXJcBdsgFFtopncEGlxWxIcvbCC/rBnTgkP1atccZ1G5rtTn2gGV6eSqZ7UxkwFRRryDXD8
86x6aScxc4A/hH3XygvWJm1Wphc7KPaC9Joj/1rLySNfrEGmYl3jzsnLAfVnjMeQEg081ijFIMB4
STHc86QlkWFte1o+dMTIc+kq7r6CPBVS1XxYMMRZua3nlO9hJu/dR8MGDyNnqwatEZRuO9gDud08
nABHLvjw4pa0ObGUfsied5HJRw5ON72rOO0qSGiqrmzgGWOsvtjBW8PoWiLzvc8ukTbDXXVqVll3
A36PaeQ7wS58EXGlWmrbK9VHukr/r6WhMsUTcPo92lSWwoHmWeFvyPYxQMYu9UdnyGdl8NzyCDEf
XA73WneUnyd5GlBFQd+LVHJkcnRgXu4usptF3c+FZ2ofv+z4bBiJ8bQFqC5sPseH/NUKMV3UUFLD
cH/EX18Ob1oNXr/2SH1Gq+3XQ9Ri/aN/yKw2mlIiEP/E9W/VHQ1Gu2VQblnRRJ9Q8wylvE+FGxEs
zu5MnOB+jjdDocs+Y27ALh4RjYwiU5yWPrNLzB5j3ExaJ2vUUNqyrH4ty5RCtTt/zr2NTamIV88s
ZJYB75IZFhRcMEoVyvfM04qnSliYncGk0eIQhAPn+fnPFxqUjrR23nuhmLuoJ6wP54dau2X82tzp
MB/W8oNd/NT91ECbCWD+S7eVjkElRsXYTydT9TUzQOD+gkaz44Ag0NG3v3uXQL/ESa/VgUheUoIS
6Ql16SbFFoJpVMHmfmndZQyXIFH6CFiDbv0ICJL1kv6OAP7DO01zH33NbVei83AgYjgeLNwv0Nci
dK99zsN2mfgQT4iCfWZd3M/Sr4Y1kCxGVfrT1GAf4cuKawQiC8reP5BVPHwEuxde0CjbveBhGRnV
hVtX3QqTePwuaKDaqnzPIAXWLxkzS0Of85NdnmELK3MSG3zNpNwOiIfd++K9+haBczt1bkfUE7KG
T2QqbeOLeVzw6dKdGsiWrh/YcWK8ob6Cr93dYiL4LhBUnaoAm+J66zAYhUzIdNhcLjx+HLdiTDe/
v+lz1b7j6/6/prhz4GqC5TYx3siNhLFzSCekQnw/t+JW8Yv19OW1cd8XzNpncH3jZw8DDY1xUvcG
ektR0S0kxgfwPNeQO4DghMHjo2FAKH7PdYbFNonA3yRkPwGpdIRi9wZus0LSSKc/vMUJ7U3lcuPW
YMI4k7voa+/J1Mfebv5D8P6Y0yR59LoC5wLYjQ3OWXLuzLGv1vXFIRCEygvzN/MFrknBx/r6qHF3
TjMz+1/vKEiet2cX+GVyV3hHfeR6zFShW/geBdFZjwbZ3Tjs9O5ObY6LDqiPK2l9Xcd76ZwjndNr
pnA+IdEwz/5PwPcbpvwmhBqLWvIhyGHzR9yM3XO+0QCpN+FIMh5cwMyZWotDdUSpfIA2DFx2z96A
Ea08lkGfw6B3SDL3p9dUzfo3zYkNEkVDNCLAc1nMR7Bx54CS+nB2XLEtyfQKvFMw3sJqemLUnBTH
9LwkQzSpZwDbiIT9t6J62ZSPZgMGYv3RZriBT713o6VWO9ifyBYSAZ7xFU2mT6l7alrG1a0pwp9H
OeK1QPAkJ5WJv0nYVr9mZiZcMZCjiRAYBlXQMLrXdkGb7kq3H8Rg5PRqieBMdkUs7RvFnQYk01LE
dvpL6NjG2qgM1yOKDnfVhCRsJti8d74mAJcRRrvddUFXzWQtJs3Szs6NSadKzLmn5wVOH7/hdqgN
eV8DdVz+D2A4JNWaqxL2D7dvhTiTfM2R5w2IxqcZVYVX7nrxUxVkDZXjsPaXft3QbAjH3dEsqlSW
jv66iGdRDBahW9loq3wybnl46PfgpLSk+OqDwjWrF1E8eAr5DnEhSWXp2J0Mvn+8ej7hVzIDl472
6Kb/NDt6IktQdpOeOdWAX0SsHt/DUsxZMoEY1ckaROHlQGQ1j2Ha77pEQiiFOO6nQRs8QlDpCSwE
U/W3XaXlsHbMDcLf8q96rLatyEy9LAQndDB/F01p8LmUtqp+UIBV+Bm2C+8KF5ATFgQo2liAudkJ
nOGXWssDcmwoLblcAxUIUfqka5SLoiQbQd3/AkgAO9U6JgU/lwL1JKxo7QzcTd1bG52n4Lku2Ouf
qNqlxYuoM1MBugHbS7jj0InYqlHNjl5HDca489Kx7Rx8qoXR+SFd0GYgkW4a/iBcxVksNcvVqSgI
Coo3hBgljAlFUbgdrOz0L88yN4xKo21w5B2p8LA8Xcqw4r6rlVCY3GTDH90rR1+sQy61M/L8Vq26
ItZR91ua9jWFNSjdTbXX+/UIWq9PUj0AoVHKIhAd0ArgfAvWnFz91TC2aGTy9Z61r9r0C+l2/WBZ
pZ6IDEtsB8MJYzTwS9Dzous1RZKqH7NIL4HJj4sa34KQhySwVX0b1bDin7ucifO3QObY5wJEAVBY
izJOg8zVbHjR7jV6z0G/9ZvZ8dGComGJhLQkXIw1QGbJnJ8UgWFdA1R1UYwJuZ3K1Q2ND9lkSdxA
L2HIfE7GbparQ3Td3e50LiW83D784TkjDjlHBRxEodP5leM5wxmobTXMnkDVUIzX36kzWItD9V/8
AyMcqombIg8N6VLQVHpCYQ2GqvvIQPympnpXDtMv9s/PylrTFyhNoLVmXadpHQq+oiRL75gAV4V1
0o3veYEW4GVIHDYQM4DEiFBZMKaLrsSccmrN6af6V7GtNAdAnCbCfwv7Souxhw9QY2CVzPWlpv3x
EWwDJWg/CNr5Jd+0CStxRZL+JNtYbx8Nu9adkuRHTIu4LLN609DRCfDm2zS3DiXzTu8MFhkg6P/y
Gz+Un5exTaS9ZSebZflLK+jRpALlUt+GJzZS5MGTbLFelprSRyh8hnrdB6gMOGz3roFH/87p+KeH
nsjJq7ewdEQ2jRwBqi5w8YgAsH/VIXvgzmohofUw5qxjAGvMX57mim6ZxHwaUIyk15TIkajFs9DT
WTcuWEAT0DqY4ieX9lLy48P87JOHiGjmO/2qFj+4XGXdXjMd2uY9V6coQTc7BMovpb1AuGg64Knd
XCpWmh1q0pL3W2P0yjJp0skdY6IcN2oCaF89k/gd5I7somhkSYYU/v5SholBXvw3U9VweigG8OdP
anQNFqo273d1Yg2VfkprSI2DFYhI2KIjueQfXRCiFN7q+vyyqrvWJV0me0u70a1UDwSqXalV5Hoo
Gm8W7zBtnoz3QJQDRf0TgOf51MOtKX5UrAzQPs0FWd889c84rJotaMzG+uq4sLw5d8Waehw7A/F1
zSVkTrtBhlbIkcy1KG19FRt6wxO7WCfUWXof7WAbS2onXuJd0iNzv/3K+2L4zOaa3Ndhv58JG6pc
TpVTIvKBGrWl1v8V4RhSg5q4l0ZYyvNsINaZkXaEqbYKXmNLC08+bBZaFZdv57SCfbfrFteugt09
uDZpRSnhiT7tnBkxr0ihqRQVI3uUSxanKWK3RDToyzn676DnYRQFmgAVTrxrYQDtK7ZbFOVqbUw3
foTZW1CUNbkepOkHMp7q0pdfyVjZWUGaH22+PNC8UPT4uqFnKQe6ZQNC7HRfBwZYxXD3xhNGAp2j
vCv6BeC+laf8VQnKH5D/4S4G8OmJ2qbjcWqCHC/P0P5B0fT4dk+9Zi8vrw4/dU1QpBAFS/cPzH6P
62pSA/tGPVw6gVXxvg4kbUWr18N3wuFADk3+LBq30lVdzVau4yrl4bZP+5d8aGpb5POfakBrouDR
oWUSei/cqByTWxcZHlGQuGb3Js7RU6JVZWkPXTGdLz6aiclaSxBhgsKks+Uw43brk6jS262juf8g
0fQkXe06CnCVVqghbLb5ZJw4k1qF1JYcTBrTRaWAlgkMtDjxSA4r0/NvEyagkTQsBnOW86CsYuPl
2hkXq7JVdiBAAj1PmfviQsm+gR18Q82dkmHJIuwAypKuuHG/NNRa/Ij0ubwFEgAsS/hsuBOfCIgh
tht9a665/efz4EC7GKOetpLT2/xM9K/UrHOpXwcrAEta5bf/WuMhYdJ0aJr3f8VfaxHKM4QaLOvw
NQGrNLNrfHQ+G205uxqGo7DhCp7duuDCz2NxWeUcoLsylNG979VzunjKja8IP5I64WlVoRpjBOPU
kjoWlZTc0WyZrnhgxSVqxPU9raKR9fTj44g7xtGoD10M+k2Uxtji/5B9I7XNO/S8OaPSDS/t+ck+
UmF3Ul0Id+RuLphPizJFeIx6qMpM75tPQZAwT6tyhDmZxFUeU/sgnhkjEDGbbVathzLsufJzRYTC
ajvS8QhjC4BREo0dnBMRU0APT74I4Gu4gkeBF9i36QY1svBHpjKnvEidyJ3DOrKe1+AeOGwFV/Up
Y51b8MzfK8hl3/SBgWx5OyZYH1zUZSWXK6AyXv6ebL0W4Ed5OZztLEpC4z1LjUKS6sy15yydEJpM
VR91ddJ+s9td74xnAPR5fvzDiHknEIC7ryDPJgp2UNU5cTjV6J8DHavsd5HyFXbnBISki4EGbNWE
TSh/Qea83MpL0IFYm0vGOV9UjHYsthmkCdxBAqe3iy+h2Tyt6LpdvNjRP9i8ZuoVTKTOB0MPrSKq
kZ3mg7r+wVMc1lZUEJyoWKAfEk7KYfS6UlpPjc8TpKLY9yKKe1ZDD0LqrFKycHQ3bS35/4Cj3OUA
6BS+TYYGHNQTYzvdJBh2r2iBewX32JhO4Zt2nVe2dCkR055GIgdNoMjiSyc1m0WrS2fZNMDe05R/
FmlJh0jpq2IyoqNUc2F6teLAEybDrz6osSW0F60U7YnN72ZHyNj4PU/bPOBzwMHMHKzzpF2yUGcw
beRuHF5wae0tDJ8HwVavRlr31dxToWJAJLHTFhlzLNOd2J4HmWgacC9q5C2+/KmJM3rcoeGNmvFx
jZ+ckKWQ3E480S+4pqySPkfIMTdSQf8drCHn4nJRpvLMgFgHkQOViI2Z8Ov9raVAU+PdvXFfwDrg
oBEFrot2RPa/KWVsldqgWsBdu0fYYc8YzlYkzwb/Idqq2V5q55dBe2L4ptNUzqAyNpAzoESDEFnC
FB6Y48Xfd8p+aLBh8QioSCVvixVhEMwD6+r3qJJkObUF8RqIoa7j4T6cntSs5RiaWrLTfD6IaBIp
1L/i86LNu7ThMWRyWm83tQNNhYsYfAcxU3RC/El+MDwZ5QdXuiVfNEIi6/Js2f1JN4GamPcypPOI
oHQlRhIJThOk3Q+oQQvWKkSQ2dJ5kj+slC3pp6qn1fxQKYi2M4+HIz9Rrq7pMt13JI+1EnI9kTGJ
6XutVvw6WZcg1u249e95R7Qoy4fjO4JO4fMyk0jFBAYXEmlc55DzX7HYDpkvw/5IIvsb9EnGo1Pv
sKDG3nSnp1eYmHxDpp6iNUgEMlQ4rQX7IV92TExf7cNbyqK7ZNXnHZ5OUIhqRjHtqRDHofavAwT/
kbTAWNRNKprWnWdFbIpowxPMvqJFsdSztYQ48DJm28fNhyelmyan51faZEkqWEnWysZC71MIRuOL
ALgP8IhPVqrBSPORmx+wG+hw/diR/yJ1EnHFhGC+3fA8k3qwqiLmRd5wOcTka9fUoE58bVCz+c9C
de3CrQemdEppejWP1sHQGzxTCh8AjrDStVEF0wRic9UKDE2g6+vZVZ06ko73alUgsGl3+DEXbSNg
ElJgi62VhJdHw+egdFPAMppZZroIEaEem5COWCmLPqRxhiMEMY/GuUrUw+FVTJv0P+G6+WpwmpfV
FnOrMoX/LfMb0Hdw70VZBhPn+jA6nv5JGeS5XjgAgbL1Rc72nLnS6dNHMm1pAw9dlRfjI4Ac0MaH
BQn6pf4PL5V7ThKNcvJzFKN8zSk1Z3y2+w/2c3WS9+9bsPO8RBIMOxBxMVRSuaaP19OokQ7EWdHp
tNQN8LdTmvQMZOCJaVoeMuRjVHOTXD+4hfL+tt8qkMpAUAVVBJT1LKtvaqsM9hHTMUIV59jBtBX8
C9gpzJWAGvX9cYk2wVIWaBtXiu+S4Cx/nrjaP+MBBiIOCHjZ3QVMRHtlR5xl8s64V9TCzoxHzOgg
YAlcNRrKU543Bj8NnqQaRQ1dOjOKl8ecTSMxcxDX7mA+IP+yb4gcfjklU3aThKq6Am8Gar1bfnFk
Cl5DxkQ6zBPhj2xoT9futz9mhemMhu/69IuK7FAsbHtvHbflzJ6D5EIVnz72/ATYth7NTYf59XNW
6gCYiTPmRgf1ouVAwDzZ2IZCO4N+7smx9a/z5FIvkAgyGk79QnDQBGflN565mSdHyikfQ9ahnRXI
Qe6aBSZUhvn2Ju2IsXTR/NWQ66x0N4ObK/pIgsM9PGtqMKYpnwz720CjFVas10IUCAKzmkKcPvum
NKNo3c8AlR4biz5sV6yE9xK3j8t2aG2I6X7g6vv4kJzDoSQN/AA700KZc9hU672Q9fPXZTM+q9Wq
sYterjigY8DWAGVhrFaLHSiSMckd5D6W8/fmAji+Hdl5xFhnLhvWdpVLf9rbPyI6SI9KoaF43cCk
zk/XE33GRO1YzZziZ21ZJKhUvfJMo5kciiux8E6LleZDNdiF9U5ewX5SvYRAs2qWlLT87O0rM2Wu
LXJVenZNXjXweTLFL8x2WZhg4DGfgt5YUSgbhIQWzZ4XOXmzC69FVXnbkWzMPT45mT6EfHv7pE1+
/MOv0T1adfDvNGfLVgO98IJVqExmQ0dXfXIcy7JEAGtMx+yYGCH48SwoVS7N/Xvv+7l+wqUMqyTu
k0haktTGAXricRKdMQMs342gTGoB/7ZWfIZ6QL6Ts1C7Wn1p0vmQxN3LKBzdAmaRAd6+XVlVz4a4
iaTTJHoKVmZJ/Hrq0fEJX9XaLAEf3+gOx6LR0jJrR9rQy7G4pvYObhemjnQjIyjR9ibuoskoDyHk
kFCcgmWPlLlEkCFgrekC1PZT7FgDQerni5SvnhOTzYA57BDtjWbV8SEXlKJ8FEZPn1Epp1zJ55+t
SP7je8LC0j628NV51g+Wb+1IAXK/Em7Sr/Lny7NYc7EzxOUZuBXWeOGgWVb9jH96MwtIm7xiKxKH
pjqwhrzYy87gI1Dt5tbk+4zpyQyiCJpXnJ7igZkNZwUf0o0+AMoIIgIAKEWa6bYsJxsvZjXj0MjS
80DgPBP2LtP1ohuDZ+rqVBJpxEdODN0bAzRGGfUuKYnUsBqoxC/l1q2iLzKanTqJXRUN/GRceBpJ
f0/MuaFgPmE1Ob+D4pmsm74++LC67wVrs7go7ngcMq+pirkR5nawsayJKonus19C3GLNfXRIK6Xq
9VPsxI5X0AYTqWI3WOIdykYCjUy3peK0eT/5MCTvP67UggiECzl7HNveu64KkIkxYKFkaD616DbT
mqx9qU4FVSd5pLMhkCez6akA+rSvAT5TjdEGt1/jadsswRS8vK9IZ4GZfRnlMl13MBicSj6aHqko
4UGkFxq4m2hP1wIHVkSQxuQn6nNhaZadKzmdCrzbNgd61hi5NrboK4QgZxJjje0jpcpxocgNnLZq
HZpSaNtVIr0aVwPzpwKUbxjTYBXD9CwuCceVT4/NhpbPb6ACuDgLERre9duShN6CweFSUxEGnG+6
Sbl4mTHZsFQgEwbzRlVpmN6X//6b5tac3T0JcFP+TroYPc/sjUb/MF2PXhwfQE+bc1Dw/uFLHRs5
RiAcaytkqg84Z9TzAfYNK1WNZFS5FdBnfPaDkJy6aYtFxbG+pzi5mmvfxjzgR7CXy0aH6AtQ/a5R
VLcrCYAAEMBpSFPQ8eNOq7xvHTzYd19Kx8mW3smeH/tjbZMRMjTtbKrmvYgqfEcYSONycB1y11/x
JlL54Txx3t3MF7E7E/83oL7pZuNS5BfF+XWdYR+8cyNBn2JFO1RdQtQz4zOKSOlSLu8au+qxNxES
YRROdp+YHFy436k7znAhF+4SbNrAqah11oROXrE8ZxKShHWfgIY5k//KIuTot6UqpYQLgz8Blf6V
8vLbIy5qUzbLfsgygmZ70O2HXxfehY+cBSBhw5ZEg8OCfFS3acon1Y/fzlhsWu0I3D7HJYpcpVdW
5KT/TSzYRN5tF7wW/hNRSRVHh1bAW5N0S+2Sq3AmtQZbX9FTPst57QL28QrYmTKbO5XLvr070ywZ
Bjz5CjwwR919g5as8E+6t0Dg/ZhxH0LRsHyYbqnK8j8Fg6U64S0wIiZQYWYtDdEZtuQ25ljwEXZZ
MLpN2fJeQz5NWBZeGAT/HQ5Qq0Y/YkO3sR8kfJzOMqjJ4QWxca6RFkX+Y0hw0a81A5B1mE2Kygqa
tiSMxWQwo72g3fyVrIpXDWEW0W6b+vyLVV7v1d1JlkHxIOvSla12kMt3qV8D+EnzqK2Ep2uLaXRn
ERLBhxm1gZExeJWj1s5XEavSLgRxInCFZpZuYqvNLAF3mnAsyRSny+vRrPyV7vDJQv5Riea+8C0Q
A8DXLCD89Tw1hb043wtTEhctlj6FK4e5HUOIbVWzRRzO8dk8DxKMeoDVq3ru1f4V0N4VwKM1AEUr
TuUcWJe4fNlj/Ql5E+oHxXay6bJcZjUj9y7SC2RbwSbes2eXPE8c1w7HX0hx3OGpC8E8GD6BZJJ/
V3sgFGu5UBGzBJnXGGa6IoVdLT5t1MqqLAgqkeMCfCGVFVfYe00JQ2BrnmDlm2gUUMM29qKvYL47
26+8gjxwEWUPKlaS3ce9gIHrtfAF5fFu3kK1/EUo6+cPIbULNEhMllvhmPd88dR5xfvXoVAq+ixH
O8J6Crn6ZUdi8uU8kdgNoke+RULK10UfNLD73t4ZAkz2KSDbMfqKwmEPNq5an7U3QDTZUM4Zy6a/
sVqOR/AP49Z03NnInOPdLu2xfLetttZ4Ksy9vZjH7Z5D1JFDgHedxVJesfxwzPJbKT87D8Qtc8LW
nXxs1RveAD3jRjQF1PR6IIJJCYhzF+tcIW8JJZxNlCcPpqDOSrcs9US7YAEvkrd3zYNQsvPYv3qO
5b7CKAPbJ5A2GV2UMV5hRZlJj/L88+2THeeLF4/iRc/3ojBmSWB++cArOg6PvTixONTAgh6Lknpf
zEtzYZCDE+4cGoG22bWpp1hyQVXsII5zbfNeVrj8FzoMD1Fn0YU3f8meiK5zH5Gh20b/eS7vIPoI
yqhtBTh6T2HjtTUXpetnP0de1y1PZVH/Yh9pEdiKnH6rn9jUqCZo6FO910qO9Mqee8oAu6g430Fz
QjL/zcWfLDSEhRpkVgv4bb1SldLit1luJyI6wQSJ9Qqk1VcLiMbeGMulj/9M5JP+lUyFyEGHQMhx
LnhwURyqDi7GL0zWEDTMplhF+JhaWSpnDwoGgPVKmS/6lxzgIR+dc8lopVXxhmWiVW/+Pd5wCvM1
ehDppz6JOAdKhkNu0nGBCe3pi6BOkVZ1BfjRvswAJm3LuJeA3br+nbMcZgHwe3pFAA/i7jf4maRq
F36/v8kG6kKCHiLWj6jFMuZ0LeYNLFi51lOhvfoL4HxYtNYvU7mAZ+s2JlyIgsEayp+Q/nrvJ/DU
/PgLuu8MklyXDVv5XW3/1ZuQtdN1NV4EqWf5d+rY29N5mHVkeT+JFULyNUWPKmPlsVyF93ZLdU56
erjdN5Jg+p9/dLn0uvHEJ1cYT+Tr/TyuFdSYbNE/+J+gje9qoPCYdl81hNajinweh8zTxrJUe06t
QJTpY3aJb4fG7RxABXz1/RiVadlUei26rJnA8FdTrwFlPSv5pw1Hyjejpr9DsmXUMXu7hh+iNttA
rtJNKD2lpS7zwoQTW1vGB23L6dEMsVwwlbg8fKtzh4A0fs86T3ZCuZsWCDif0OMFyzRSBBxbFcuk
YnJFR1POGsoiTLTxMgqbf5kYru+A9sbgl9aMj8VsHcZWe9xAfcpOvvf8/1AivL/ZY5TAYqrcZPH5
iN/5F6vSo+GF5vGRBV6l/anBDqokduzV+pUqx/Rj73flRq/AWYwk5Vm2j3Whs6q4+9cBmzsbQjvZ
AQ5qcCuRVRD1L5DQQzhGddJJahbRnSLY7QF5tG2swjn6p1mLHRK+UKfLpHRbrWSjaoxTaIJ2FfUj
DZQsiFfw+Zf/rYfiEio+G0dCAykaqtFoV+SsxqjAAZ2EBEO2D7f/7XxwRRXBftLdUko/FTM+bGNG
gHRb5o9s1AfB4SVpa0skj264OUWvKYGYQpAFE2AO7qUYspybDTMt4SFax3sxlKzYKtulBmuPDn4K
tpgTsF38nEbldWTkUTEz0WiTNHKXUAQ6N+EU6FpcmM4i+Cii2X6SXvtEuchi035TTyfbC7r3GIIE
JZ8Ql9H/VIj3n3TTLX45IgN8mbc8GB5l9IL2dPZnAqoudsTfosJ3LVA9wi6evZqd0fSTuIew7/lq
S0YCOMGFKM7VKCbh4n2HfLZk9k+4a5VRxs8LAkI6psw6m2ym3M0CzCV8ksaOP5jsRWs/gIcFJJcH
JR/ujrM/jeKycjjrWxggfpiFOYMBQYbOBt8uhqTUxacUv8+1pVYPNQ93jvk/zHvjjTTURiwSCg7D
tHUsii92Z3epVlbbt2HIcze7eWsn8M2qbyau6Go+TXwsZAVvKHyiwboI+Ex6AuAvtqWU7bOZBP6p
Ili8Bg3PU1WQl5A5bqQt8uNnsMKeHnIFNbLn/oASz0JOuoBPIunkHmWPkJXftm/Tm3Vf3J5XTR4Y
5zjBXCa+EOcl9ukVm00K3T4nFwO6UiggDZvhbg8nyG5D9+b3QraJvep5203KVfULNos0pWJmpwqi
s8xgPZPws/BUGx3xJBRmB1w0dCUjFZ5z2M0wzz3nc9XowyvCAav3hxaYJtnKjb8baF/wsU5y4JY0
+5GakYtnoitCRfkFIrrFRzt82KSWjF75omMEBnVaOXHbVnmLaJRVvNlHW/neQoygjGEpROMJA83F
YZjUNLXYI4h6NyhE13lwjiPEiaeRDDJqs5WceHIyaOwxEF/OUirRLHBKEeF55a6U1UNb2CZZOKtl
zUYBWXBIpMXV6qVvsSIxQD+6ALMC3fR3Zyne/oOZCDvMnfcuJRvPFiyh9INWUz7G/LCNmLEtKRq3
uv/1GIyek0ODxbK6hot/VCrg2e00ocJiV9+PJCwacIKq1mMBv5SEBSkh5bXDP9jG/VNH5rei3FzZ
0Lo61lY2HxtIUMJkSfc/LMJApy92eVMayoyXI8HsHn+i//MywJtp6C4ZIgC8Rd++w2BT+1It7wV5
ODrb9RnHCU+qXTNu5jRpB4T7F9jrlxcvageNn81MYV/jYIas3GJY0IuDRvTqGsOluD0cd0aVBpUc
YydWb1/PoYPvB0amxN+Tk8onXRpLREIK0QdJMtglCoxAA2RGYzfCaLfzVvdBFodKYjZKi3WOYMX+
0SI1+fa36U1aJuuxPpnU0teaNLIpHf8+nqI+LErPg2gcNqU8N/JOh7mBeliGmFjhxnSpNCJOIJvb
5UOGyFNkAvYjAN3hGna/Xng1rjTZgWdbLxMgot71LdZMu2CTWgiMleNl6E7iy1C5ORSmMy3nWzgJ
zWfZcKsub0X1mNGaEcN+Oc0RE+R7fTaLXV9yTrJLSt7uLE/tEIFPulRLiaNKGxTkR0GjAqR6zhEc
RLupwcp3BxAwQC7n8d4wIKB1Jy+O0t6GtYBJZXTvtQsWwlJ9uuqaRCLEmV0+50IH/k593jrsMbEs
85jeX7mONj2C5Me6QkzTiFvVCzgkJ+H4KtkHAqlI5j0/LLKQfhvc03/Sd1T8Tbawl488TFvNV9BM
EoTXWsNZtC4q4KuIo1p4Kl56VBnmcjqfeAj2IuoNCsCtkzTGAY4BxZCFsFZZ7wGFsfxPjA9hg0Nj
zBDwagGV1t2RAYp+HOU0dFMuCdrWe4rKQLxw2HH3waw6C1f7iuWeWQzBFUjJXSjxupzzyWTfRnXr
Ff347HniQ8FKDCL/DokEpT431qyLbUmLWyasTa5zdUhYS0p2uve0lV1zGTBIeAdzJELIL5g1l99z
h5eQOF/rAA1RlGM5RrhbS2ZZHEsGFj4njAO1V+iRKfeq6AsImmvU6cGjl6B7JbvKpPJfjxOZBVMI
/LIThSOriGvZO3nhDkoxVd/OgJrMKR9J91mW6RZJRj40To7n+yN+2+WgwNIMSFSwk56kbT7LB90d
dPaPmTKyoMRnzkx8JEq8leOJikDktpf3w2U3wBcRZqZ9x90hAbTNLniEtpK0VoXgZfbQuTRFtVuo
OvLcjKE7mm28VVcIG0ZChJJDQJ+KdNU+fYdTrLcqaIkbGg1k0vNG6OZyKq9aWc0QME7QEbCN+gwx
HDoUCceA7KIVeZnZIm+cIoir7J9gOFvZ/oAlUKmM1ls9/AQU+5utflScaA75jqOJUjCwuOol/3y6
Oc6dMv0kQMToyRipbDiQWer4bRxm3q3RuKkfC3+n/zrOPF677WUCWotEQgg23vmqH07HPpVBFZq/
AGrTwEFeZPicVPaAH7lVEvABUsNhyprYOLh53kXhpxEKVt/WuE7V7b1yz6MPbA63CfAxbaP7o41T
ovfab0AV3fIWHEnQHQf8Av++kZsDYjPPVVMvbUOVY5TI6M9LzneqRKiGgEBWZ7d99gQT2JU44LOJ
MIenS5/uI8B51atNdfpsOkM0yZ+A6lbbFPFggEnmJp8SNH4CIez8LHaTG1zPkah4Mv6XYPn2Zu3W
1VsNfavJZISXde5juRjVAy6Jam3wmM3fUgfZJisKgPyPR5NLnIENtK0Fjx9lixOHV5nM2EoPK8Ot
1njPnrt/k87y0pSJRjEn/KQw5FETZwS/2eB3HECCa5/DhNzOFqX1hGP0h+JPY5s15xVn/g9xYEHc
famHBzKCDnNNaWW9mRNYTS56w6gVDBRoM3tcxw941JIP0cLenYCho96F5fR0m3KnGG+UMQl/Xl6E
3MkTkGBsKLVdMFzwtBcTJ3P5pSH/Ycy4Ye3eFXvU6Q0Jo936fxmoCoQkqFFBkDlH8U+zy1KLqnmm
Lkx2nZFHid+mpX3tA5rBSXeOZmJFc8veo7jVar4hHr3Tq4Kv9bX11piDfZ594F/KL/JdlgbcBQgG
0VtnrEQzH49Pk/Lorpg/eOCeL+HswPEThNjqlGqTpUVRiIQ32Qb4UfdljkUfZFia+zqLGjhzBWsw
tM+gPnkAPwSO+SklD7mY+fySX8CPPAygQzjBLCkoPZhsUZHEtJFWU8Pv92yRYVpB14CS3wxF5pXj
vjtmyHY9XbUqadtLDo6uQvtDCDU807gB07glqHDRn0/6jbZqCDLZCqSafvh5tLzWea/FfYiVVsq3
szEol0crV4l9zOgX58U5K3XytMbJSmRfDehz14m/aX9tXyxkFCda9izQO8sOj7UQWeplrJLI85QZ
nXGBfzG3uHZW8x8bHx+G7s7CXbhlueT0X8n3FtTXcJa4nbxnRve681V06kJ/HYQREAsrpk3mbvkt
XiAnm4sEdAB7sGvjB0eBhyZbyJ+Kv4eRf6KWMcCPXHnm0VYuyj7Tke9oalBMsDLPClhrteND0MvO
nbYv/OOU/MvWD+Mwdc+JfgaBVmtEYWG9AMJ46Zb8hlSov/3rAWf/joyjnnS9l9GxaxpidTcDyUE4
ooalEY000r0N9PsiNl+xFDpqqQR7scIC9YKVOeg5+jcTOF6YtDpfU7PS96CuFh+Y8X/8g24GSDsH
9WgdXe0pCwoBh/mO+LFcjGQArxYfo+zgMjvc5q/cr1Or9i5vulO2w2SK3pkBwErQGkCqVh07gRG5
G5s29rMe6jnNIwS2sKLT8sdeMOIv+VY+GHgvIlxD+7nqBDp4Fu4rPXjSvyn1rcO6nlIusLrk6fVN
XJmhPznFQ/SodtqakxBefv9mPoOqv6EVyO/aN9WG8OvjgILwrJWOgbrJVt2Pnfp5cxg/u6F6op/P
EvsLgO2sFM/wUW/cY22kmJn4NSO6eNITkrUGVzUZW4cWbGcSqPsvfEAavb7kKKhfQPqJ2ks3y7NV
jkmSaRKNJjikj1ed0JmV6+qahG0hSoK64wONX3DSYzgccvVQg3BYfJof2JK48nCL9faN/+YHjZPu
KEmXlKfjB2ynSEEJ0GaVcK3AG4ul+iNUdd+tcp/GjlkT+v4f2g8K74dPjRxpjrqAtgiO7tdXETwv
nXRe8kEzEySwRt6GKjvhvM28SU9LQpBnLA1LomfIlQAVbd8DaATWMKqmAUKHnxr+rgSjegeq3gB9
tgmTWAJumk076c761z9LrsCeokkPuj+g8fzVq8TwtGTYseMVEkWPWqrlVn+QdawjOcEouuhsy+QB
ebAOmsSktix0DFYnXCoHyqNr0wxiZX3Wot89lsv/MWCTDFeePlCjD1L83F3co+uWgmlFQKgFNB0a
HNmZ8aqD4Oo9TBPj89WsPL+CbMxE3aUpAedyY+lgbtDXgIkMTzOliomi7BsYIxbiHF25SrU33n4C
17zvvyTBfcJS43YNIk/gpH5e4GATIRcbmcCTblWVjxk1b/wpReKUt9tXHzJgmYGaI2K3t80BIBzl
2bXEWYULn9cKzXJ880HIIBKzGNCqwX/6rQC0lszj75CNRbxE5elCsEDnwRcY0iszn+Wz/kqGxLi5
xC86Wvw2bokWrja1PF38NM3YhWfa/T9G514wvHBeaxnfP5k9eH+0PnFhlXFCA0csHfGUBRlGOUKh
MalqOrXOkk/z9AlkXB1mp0MnAUhFSkjT0kLdDEgr7xD5Zr15yx4G9MKnJmDNSsZpuxJGS/cCJs2h
vvjkfBXGkvlN+vJ+C6cbi/VTWWPTqX8kgNlBTn6KGHFjqmFYAn1rOguo9lUQQlsOkZAWSmLOe4gw
+Fs3EYM4F/DxRHr4bChnohUDflYwKm4fAquTgfcpjXFzLki9sLxTp4eHkr+IL7JJFpf6kD/Wqi6B
ClevgWqqwexhUxlRNs9dqcMVSuP32i7EGxNkb2NpFWvA6IZflLC4RekQ+iJNmUubxipk1wwrctRL
jmOExIizx622EXYGB9V4sYX76NPYBRfFrwJWsWroXmMq5hZlSe3GOsihcRY9/tHfFCoqeuBJRvQi
Bf15X8FXNVsdc6RQgEemTQ9vgz9T4dVCG0vrHJEH46RJMjLnoApYiLcJNGcMM5zNOmvKOwqxb45F
p1dfqiLaIrDpxGJV9oYKBugfTJlC849bwAUlDCblU7vsMw4RWuDMrc4USzpXe+KmUOGnboLy4Ign
RfVl2xcmvnp8NsN7yJSlv7KWi4JFtCP765wtt/njxhuMP1V2dsh+iRVOuCR+fAfW6G1L2p3L+s7T
CP+Ss8GG8ZZX2NqHZt+voyYIx/t3acbRjRQIX6mq6wshJhxOxBLKe/B945CwZEb/O1r04Gv44Bi3
buIPcRKuq3UlM//YrViZtiv090NXevZ73x4RGKoWg5DRxpMEZNTJRGbOf8oRWe+1QBmVKQhyr5Jl
uAhAvrss2u99P4k7e5Afe2xSlgI/6eUSA+5es5OmJEsgxDuM3kk4ja581t2w8JnpAaeKjH3z9qwW
JM8U9K5VY7IaRq3Tlswa5LqkxbNH6GUrc98TlVjrg8TCCjSffOOLoS+Zjx/9M1G7maJ0wYz0KXSr
XpX9fH2FDiu4WLilqQVGANVIDdSZKsZ/IZBP0yYmlcTpi8UI53yEGakwW8bTkfuv1el3comjzReo
cpfILgrqmMXuo4jb7s5VcupC3ZNh8vN1QwJ177jyO40R/kO47xsnX6qxkuI3EnRS4hFcHqOfo2AA
iR8hE2c1s2p0blD2QRS+0OdpWvpEtzK+WbHKzzbF+wAlWJgaIdpMEq/f2pfCj48bKT/IQpLnPgw2
qb2vLcc9rpZOcwoe92WpiyNRG5MhrSQwsowtJkv+8+T3Q+DRPmF+OIgMjBSq8L430Oig9sDK2HT6
O5veGJwuFS71CbfkeXXXtEQz76SDDkmvwNnAxbrqFtucxh/bFulmpwuePmQJZP8rmQo1A6IxiI/2
KOr15uEejtUEFD5WJLEwinqqBqzSz2WRU3D/iDpbbpM2tm1nCvEsArxFlJYVcmESalnjXcG2RNge
8iptmPXOUo56LR0mazPhDUwtTqHWB6KNfuFyE29ak6PbaiC9dRjdxOtdjih87BiSdeCKEYxa4uwI
9HljOcWj2WJvM2BGn2tE8q4LummfSpuSW6urGeN2gJCUmR9oGJW0fXVqW/tAY4KahAmWozZr4IF3
SA8JOoOiP1B63u5ep59/vuiiYocSaofFB8M/9tDbHrmiGtJtZwMhJdCGLXEJd8boBGaMo7AdqE1s
q/DUPRj0IRwIHICWuyAf1Ep1BC92a1YOneXDxaN19lSQIIVGqY+zSLzgextFpzmO+gj7GIWpYdbs
H9STI2IERjlrnV18KyTJaKbwm2BVL+gfgA/dwlbSddvasAMr7uUg6qY0FmedwiM9duYL9sXR5io0
XxiENUeJszlVfroyvkU2Tg2JMrEUJ6e7DevH16qF3Y7Wxk3bBTNvUTMZNdotYn/4AIcUPqub3bXN
1PSFZ4rfiDZcTd9G0Y11NIpKD1iKBy6laaSOG6DszSDgEqLGQZMY61m9mn2O0IxmK5CLXoSQdFWO
la+52YI3OCC543p3MYx56oB40tilfo9MOAga5IwHAVnBSdJU0IyfYnPJdWInPLFGjxHOuolIFL+t
fJagBF+Tkcu6PXrOZQAXt+dhfQoP46GwP7A3/2mFS2+PlDFH6CFu1u41T2LBa3MnQyURIErfBdK0
mL8Ag3WYj1UhZK5gTKdIVMgEPVD19zUm9TPzs+SBwyshjyNoww0YAOcv04J9+gcXz8W8u94rMMWp
e+oxbzzeZR6LyCVlxsKy3FtUcDvzPfNpzVRhdt8lBLedKR9e2eteekTDr80UnOv1AwqkOPOf8jWi
DcXdTSxTh2zASzUZgZfndXJYeBjQKOth/2WItquTjjPXpWkXvO5dRBG2JEHFpivAOEvWbp+RsDrE
bYjJWqltb9UqG2jF9jfXHAwKhw7XR0f5sECkgXPm8wKP+usnJdBpPX6TJ/FrPQj+RDW22NimA8l+
0iGUt0SEghYgdSn5oaR4i+hAzQxd8d3vs0abz/j5x7Qbcp6p3Es3/RmXTNKNzEHkZcSshbiTN0lq
D9R5VwJY1w85CAY6HrDbRBdYDDCkI4NGc4sL9KBEpq47v4pkXKFs1GVkpWPzlAxF3q0zF2RaCKhr
1FBqUdzbz+Jfj/HqJs0URvO7HIIcGZxUmUNquZqBlBtbOvltK5vXo2Iq0X+vmv72b2rakFThw8bS
LbBs+DMLJ5St65hIMpi/GEx/Nv3bGNUZrHoo+R98DfFYdNtXTRHzY2g/oKGjFzOvFBYrQSY5HO0L
lHfVgZe563y7C9lKiltO9gXXpkE3s+aNR5o1LKv34WMmwBWtod4auB7d7+8chRyT/fw4sjaQBOxk
L1uRNxGmmvVaHbL5+zYqk3JFJ4acTkQCTFHLFY1i935dEyc48oITlvZDIitCVgg+3Ou2qaaqPt4X
Z6+vCqO9S/oXD9EbZvTEZwoaNtO4D+lAJL/MZAnYimdmetC7JUh0sv3goQSWks9jMaoN77kX/Jh7
/yTo/eZjr7PxylwtmmLCZ+PpVAYRozzClfIEWCfb3GBra7Fq7ZLsxhKZsVRu1Jaczvh4XjBHER12
l8yV0XWr/t5wwWjMYC1UEMgRAFb6iZ6l/z3qJgmqou+df3eK8W+9fOqg5/3EtDzIXdH1w8RBvAaK
cr0MbhVe4xcTAzOiiniZW9I9LJpuioVONWX5yAzgQYf/zkRbWFcz+PE6WFywKGv9Mz9ialPCT40N
bFmQ0EyyqbgoHt2Hh16ZZAuONOJ+k1FFMsVxuXavynGtSmVmGGobB7pzmZmwBe9HvnDYseuoY2Xp
ZzJJtf6aUVQwb1i7NgzodIJGLZNNEhqX5QGulRXHNJDivxrLN3xr6CY50oxMdi8WjGjflOqJfj6s
A7KuWeZ4CHlu8Mg4yCTlN5fqPirB/d5/mUodcv8pR3InbIqyFmSMaIG9E2uBqee08++25Pm6VIxj
+XAFtYkwxoWsmf0cwSyb6vRONRnQG6W3trcYsfAnMZxOXE5IAlV/T+CS47YlERC7NuqJDDmCUSKz
/s5aOYVizptdsfCY191CjIuy+CVzs3GcsmO5qeXNEsRhk7rRSKqwsu/BC8jF4jCTG41izsIuZQT+
vDFPlDTfDEuzzNQDB888uUaih8pH7dJNLjvjo7HxYxHuTV/jDH6uVNscoA9M8jwgMTXY/TMamVTK
WE7c/62Oz7/nsyBDshhX1uzZeZmHFJ7D/URDYe2j2+ZzW0JSJIKCyU4brcZLKi6RAn+j8cZG99w3
UzZhJV3sUzLnQRs5idaIbCxR23y1ubqNAGWxqmvnyKQha6AhFOnEtB9DQIkuEQXmVlSq1vpWUIeq
JHTDkomP8fxWGN2Na2F48ZgR7Dbt8ezD+7Y0FUiQgOlfa/n7ENz71nQZefeidEfJOlmXLX17baaY
eB9AwUN0O97r3QScBk5xoPJssEbvZHldHgjQzrytT1iqBXk/DCo8Tvc4eOOqpk3nS1mnKjwTYxPc
1qlvvRn9fNQ6HkJDuvZk6K0tXhycaYSz4KsxeKmL6ORIcg/qqZUKqQ1Qtcqo8mOYjMtA9DKHvYlb
XHnCsZJrK2GFV690uF21Lm/UIhbAmNQRm5NT6wFUULGEHABg0n05rzdv2Im0AFollXPscB6NzodS
GB3t8G+Usy26JJNeqb6fQGSz2CM/Uni2f7eCX0MUounzbldAyaE5LAoBZJ1H0A70KYBlbDEH9whB
EVm90hTuyFhYMm+5fn2nbxCYuTeHZO3BuGVNQJuH5QXf6/MPs7SQjaRoE+a9kVx2gmIO4elsdOWA
9PDt4lYyWCHLUB6DPvB3i78QP73LanlhFN4+TU3pVqRKaHZwl0RP85zunSULbs6DpO+w3NYExpx5
0ggW6ciAE4Z5BewjLjkhVlI6tVbYzD3UcvzxmMkFqwqG/r11tupXhrGyRKwqfpOCjCbGr7NRiUln
Wp9YUYNdah31dRoDqrR7FytGFcZcs4zP/jn0Ic/WvCYBqIjCxK23T+Zi7qouGGCKrt2MXmLZmuzV
5zhfzXtsHICKunN9dm7hbNqVfSQgOQTSbGMAMCdstUWOkiU/GvUnKto22pXy26qeDb1Vbpd+CdHT
GZV5mqt3eZ83Bymk1aFHN1GU6NNSLNP8IX7gDgVNb4te/dLAbKmd2VtEYRWqEC2bKMKekkyWCLMT
dvxnA+ToFg452JsGebBC5XVTuYUG7T4lQrbY8PYyi259ZmZmann/9HWfTSLW+4Qmvsk0mqAMYqBW
PEJp5Wmqfnu9I3QX2BUm9+Dumbw4teOGz3tUynzplKLiNknqSm2Y5ZGsYBBOK8tart/D4L9fCooF
VYTAzF5Iub6JR8uSqgjcIDRk0WSVyP8yslmqY5wDtAXGkXS7Yw5YA9MGhoY61BkKEvSwySb16df5
jN6ZbpKGWwev57NiJRkVfK6plIPwZk8hgZpVsZMv2TBz4x3LFXs1iyksu72pLcx8pgSIGOSyKWpn
yaxfkA/EUMSg36brVyK221TkcX6YB9j/7bLa/+IB6wvZI97A6NT1kQaaJkS11KSBy67HhcluISP1
71+CN5ktwkv7G9C98V2G8WrG82rbsoGpK3Eb2Kyn5VaRQ+WEuUwYKYhgzFJ+puz0wO08Ss9TIy0u
Ij8F09Bfj1ng0Gk1yRgPJFIOc7nW4ZCD+haomyExZOoXsjHjet+kGJ7qVcXUkz6mH+zmXqFChuAP
FSdCnt5lkuXkk95c3k6DXd7yyH0pSwk+YgCJLPdd9RcFSJi9lQ0JjTjZ2uqKA5A5axWE4GxN07Vn
qm86AxJIUDw8dDYuTA8UvP+jOlYm+0Uvq+Iyc/Ea9PerGmbpbhuLQipoGixqARnd0/A+ELpg926+
m1R0rmtB6ywxK9Kg+BNlrSgbucLB/aNfS+LFii+zPx8XAE3f76BfDnQ7Wz5aaBbsVPyXd+lzpy1w
JnZ3R6Snyg+fDYVnIBnzHSTcNv1Y+Csd7GdiRmiwI8Tm/z98lWC2Mm6ksycAYhIvmlECIg3z8q9v
7QMqcfArWfyyCwUzQAz6lEH43BFkw9vSYQDBET6+4fW48nuUFd5BlDBpaBU7JyGiS7b0bVnfcWuO
nxwEHn1vRLgP5rdgbvMtmqU+CDsuWtOzap+card2w5gyySIAnvPkApUSeTZKe44Ndr+TZ54LPNaz
IfbMRbbr41oCDq1VsUHg3f/vmjYJkF+78+WPnCT9thBGhVGk37ksRKUcNwgspwa8P6vjdVMk3yFH
T7WLW3711QbrQFJRvCWglQ4gquydq0icdIlUqiekHvarF06ioiCre9NANkbywK3qQ21MFn7aIaOc
Kd/IE8gstNuTnLHiao2qGeVoXeo01dsUbS8ijL5QxWsdzG9K7t6yQ22GfHVXUAlHqWs8Q7MCycVx
APfhwUYoHDxljhm/+z1MGGG9Mw6HITVPGJKFWPtG/qeVNU/cdQGgyphMys0E5EKWx4vg40g8H1+r
oIqo6vS9uUs4RJs95F3DlglW9Bnyz9rBL1v0WsE5zy8GxnMmYljo+ZksTEuEdOje/UU7bp3Z9I2G
GZ2P8VNx9VcOBHdbLNJ9DudEnFkdgonCrVBoeRyrIL9BPnNsqk49zWbwOOezjrRwq0a1d0Gp6Khi
KrAiEoh1vbnZgY/5PlNnVogMu6jGfsH0gqqBFsN/FKeNvrvd5F5BVYuASEr3sATNvgSMT0aUl353
BSEijJ1cV4vYDvwbhFpdM7YRPKap7QFstIqwSv34i5SBjmSSkSQ2vdmK8d685NpeEizzcylLbyKH
wILYQvIPQElrryu2zOiwUsLUx49H7dp0idQCmJ6Q2XfeyGsi2rdU68YUxX80JLOxolztaZwvlXln
FwNxgihu8V0JhiKeub7hDw0yDYawz08tu1qswNNwDciIno7BRsckYKWUq90JlnmfU1exYHG+TyE1
/Mx/s7Xivam9Ie77nN3gxLvy3H2eZiTIdShjhTuUXSN2SpCarYzVcRi4B7y0Fp2GErI1ECoCIJZb
PzA+mB2QKjOcaqDDu0TQnssvB1dKcW3DB9X8m1516jMnO2bMtMfBU2F1uzVJx9S9wkbtrBNTkPS0
gA0voqk4tpK39CUrnQ5xWuHYcOxaceIMcq2msfwx2z5dP0nkIDPrHKLLJ+rZBVwCW8h+CvSTJkXg
sX6SDiTbCTrDjR3pppy3u7raHtzOQksaXiBigqYRIaRACgF9Cbd4kPrBIq156TsSoS1ClzzShPkz
vVfurKMD8QPzBlumcXUftQTg+FN+YAoaozktw4iZjwxFEuRb4dQ2q6LU+Xkul/Kx8CHZZixK9Tun
uNqBjCp3xvmbgt+CulKmlb1GjW48lmfuzEPTtQrD7llBEiqv2AtQXcq7iqa/oW+Eu5M1QVY63qVR
NvLYNmCOpK8IUnIwO5u6Y9at40xs8J/MBp+Bd2Xp9IyiFAdd4f4C41852blnP4BKP4n5uOY9eQAV
0R0bsY+/sKLiHHjPdp0WFnB5O5SYIqMcazjsJ+J4YZGz51LPV9U6YFZZyk5rgVzx1hSjNvnelftd
37NE79en5cNFtT/u5A3dhSNXJsW6ICH/PyNTXdtJHrWzWxMhNf/GVRYresmedujN9iwvXKwES6JG
tXoKs8F9oIjut73d0kd4b+zgSlPLwTYhhHfB15VADpFJj+5HdcwSX2OuiEvkSrvBmf5HpOVqNWal
gJXg12tag+FewuXyFnA/5aKXMTN8Y8Pe4fJC7/U5B+ycUuRB8IX3TyAhNguk1XIkchbZBpSkwnrN
QKuHukJgIqnTk8sp6UFvOJ5/fnKCBalbe/KXjzlhdJF39V4rE51fU1pY/JTYE9Zm/+tlS8jclDQQ
x7ID2rOl8ttq9d/i7q05MjcXiSt6/AXYm3kacItbzWyqbjtjVhkLCIofGSK+fyDxpMwx9v05fXF4
H+rIQtthrid7pLTU8l+Gjk+F4rQzu8Tr0qKzniWKbNdlnMUBvwhDwdD3xBWjIWyVlhFf//P4SLDm
rCNJ7+BZxm0+SvB8iI7m8MMffsbu6uPfck1bG0J5RFhHfM6EmiQnRci+F0h9tqYKsQnjGbovuwH3
6/gQJW2lr6e7+HprugNqqvuhfVYtnEgn/aOUs9dcyDruvQvbciA53Cn6nb5u2ETV7AUAv1MGVvqZ
epB1ReEJbTplUfsrYuM2QPavRbgMIgFbM4UHD7/FCUmq/NXwnjiTx06zW2Ur7Eq9JhCDlOd5oeHL
gssVZaQ8JqyrXX+8pJclMis85/YpFpuVxmqdp75HSzm47cuQf8c6nwr6us0zOlHhiwmdZTo2FKKn
zglM2fAa63BlPZDSvs4p6QnXkUY5p33lSyZQ2FPnx1Q2csMrgiZnNu+DLCnQQRNU6+a6Wfpn+62I
3GzN+IuUIOOp6oOXjK2PvoXmoW1DHdIIls4Ogw8UV/3M0zv5BN3gpBTJ+vGdEkGsD3SzCujY2/dw
PQk3zZk3987ASm3a71HrwrRMhDfG8EI+DugaZT9M1s46WlAr2RQJFff2hkXqEhVc4F1RS5oDS3zY
Zv+r9V23WZmRmdvSqqJBtcKzPLbQyvbR09tJQikWIW+XB5XnUHmu71aB7nTvAA6pHBfVzsZ6DiB9
oS3l3ncpaTjDsCiHAagAnP0YvmrWzWJ/ZyQsKE1A3KrI9FIujll9xhI3FH3IMx+cFn02TpHDF5qa
OC7AXAGcj4y4Z8/QSHEsmJSR362tOW/jjfiK9DVwdP42AljO9v2f+rr59qYMXTbZLQ4GkQMT2Oyh
KNRyQm5WaCcLFL6s+RY4quCmWPdA+injTPq4mzUx6G/GWD4xorBTSlkDkNHC5PeC9GJCUsMtzqgc
bR5TD4Octb1q05SiJEXRLfOE8bR4Rh4t10RmjsAtYh5Ol8jV/0TAxGrXZSd0nIAac1SKVdw/Agat
PugYAh3eAlfXm1NkQjgti84nwhnGn7tCp9oXJgehdp+Zyxv3wwHuomctfubF0fEdefekwPSwcG0K
xOsg7Rxq1OH2oJTeNRSs5cQE/aiiv99TsWKVz0yMubLrruDHSSUwbH+an2r1WCIQZaqAv02C1rXi
aYZhr6ULtO9hOqz1+Dj3DZ45qmhAA65xh61LL0pLiHtt8AndueFGXz1A2VdEmmojJgV3bhSfaWUT
zpFb5T9dl2DsIvZxGJPGK7izH58i6BWgKassUSe6RlrTNI5WzC5eXxXN0uELbja98xASH5jO4a9U
A8ZmCvydeRZV17H8VV1yoja/V0v0hXW/0mO+7vYlBYP4C3HYVx6OAzgcg6y1m+euOdPRzvbDqL1d
5aw+EgLpgQi0Zo4iwA3SzSlEPVL+EdbMFT99A33BuGt0Kph5SY/sXBkmMqV9XqZWHCQrwWp5uLZU
vnYaI5XWSA5uE4yAvaOL6hqF+aRw1KI35vD3xQHqRJJJnIm+/lgJ97itDWAPaC1jRWlw+4HOB0an
W7U0aeT/SSAM1TMAGpIBztu3r0uPp5HCk+O8bidfE8wWBMT/5aFX2FKDMEnV1dovwXemqW5ZCqPW
YJFBu4geLjJmNsORPYVjaPSu81kOZ+JmNpkYtwPrwDMKUMtK3VSyEAYdAChHeyLwbqetBtnvwQDG
kshSE86CLEIJEmizcP/MGYqycyIFXxHD6pmKKIJYG/8SK5n/WVx3jJnWAqYsabhfREpoCCwXr7Hb
yaH2GZkh6UtMNOlMx3gdxazAnIM/yOYMio06h5TIMKvPflC+RTkS1yFjxv404jbf8tL7jPEvM+93
pMplwggFBqZvBsbFzscligGrTu7FGSvM/42rq5ytsUIjncVA6CrS7uswUyYRoMgmeQWPDhmNqf7H
smYuN8LtneyvUWKobqbLrE8wqIw8gyaApSI3LpaoT/QoAAQAZKDKyWeuuCKYzbSdvTVL8S8wLKl1
j9VxXJwn44T3vRS+QQIduVaRqF1mQmCzcVCjwSKmXN8AiEpY1uAUSF4qx8HEv9xHVTdzyy+adoPz
klgY7dx+1D7CQEh/TsGcEImuiiG9Y9tpQ/G6iAjoNsd7NaMDGIN30sahiem4C3sncmI0kPMWxemu
f20x/Wx1f4Z6lLpALO2hgWOmizEhzN8qeVMHiRAQryygK7xHzDa+b9jibQBPrxhO8QchXxlFL5IK
11HZDk5ABsaQOgzQJKSO7NWTAihxwCRwpRci6VhNZz28jTIZFo2mblbvbX2xpUhDpJtaaZiWKiOL
Fo+sbTmqPDMn5hoY46C4tWjyaYvxjIm0H5XogrHtHvnzPD+bX41eqetEadX/60vEIoYRILjf7n8U
8lXy1A7DTD1h4R3sy4V0MGD0QdKSEBlXcoUVreXh8jUKXuaSOragbOY0uNQlM6ntp7qqUKxH6TUn
Yy9LEahihfgzT8U43JkNYAx89YkIpTJyENqGvHEswqZG/x2SWzKLvlkYd/4mMzAaYUUZ4QZBChI9
vK0saw4f6xn/8do61l6w/nUKuLXFfa89hKbNKORafRfqAJ0ToBBUEzbqVh8Zut8H0fnH+zVH0x/i
YvZuMhttJZOhXwE9U2CG/mhQHK40ygOwLS7e+QeZfNz6Uw7qVpeb2L5zKtkATu+g6+CT9dnWz5aL
0rjv3Yxzbcmhb4LOOkzlkGxMaMBHONKgLs9sgC/zTUfCChqy0zS3wbc93Bl+aBJSTcjG0PyiN7za
9aKnyilHs35uQFBNQnajzC4dbLXYIuc8YNbfraNiaHVSy6VPrABp3V1QqNiMbSrntg1JbH1+AGwp
CQqkIfw5N4AzQJg1x0cC6Ob8EoXgqc2HtqpSNQ/0+l6amkYwtBP2VXVbRjPKvsgJnplsFKv8NcfW
+rmipmmAOagtSssUH7I/xjyfdEegttWZhTxs58oj7uLvcLmKI/G5/s8Xotd1CrhyqgUciT5Nf2NP
dt3PiFXs7Tyc2RhRnk6P0Jn1o/aer7NQdeWW++1K5wwN/MoThoqux6F0H+ZR9ATQ2o5sLU8j4lf5
Te9m6MX+Nly7PFLtANoSx0qqyW1XUistCYJTGGmKSgV1Fo/xXptOTwpEJk0FboU/A2xzR/ZpTc7S
k6IGvrQ4EAv9YjKrVqzSoiy281MeXZkLNOVYSWhYwZXUoKBGFBQDKEBau1uLQELQeaRLnxxGl+y4
P202HlGbR2dlJH1X6BwAccMwSSoxZkUswMW3SbePi7b6kXODhNzMXlp5PH3EsFo8bjZri5ECATqt
blCYqRHL+029jPjDhRiMx8UN3iEIGEbHEyFbrA1M6KjOYo+TonGIzZjImgyns2r+Fl/zETbIefsK
MjzIRy4/V5sXH0IHEJzBUQkFkKMdsuepuhF8emOMW/zBEzGfQtZVZZDC9K1+EPguMpgjMmKKOY3u
H5LF4EkBjXhzr/0rlRWpybwn8IfTte40zPsq+RinUmoSsi3fMG3gGpdjx+gx/GfF+xN8i1Loof1u
WVbDaAL8odEwHULRdkzYwrDPxxQoeXsmi7nGWL/lC2mjKq5/qJaz2UxuQ6mCmwe1fzktHSe7dmu+
vCh2ADR2Tzcab6R2jfD5+SWfWBEDL/fl8p2hRkNAiQXaahwE8S7GnyylT0bJA8VJZeiD57hjIjhG
7bRXQ7bZNmVnAnMQ7b4Oq+mR3lyDB4DMO+fUcY1MVsPpAGud6LMIyLWlOi88kNOJioffqHH4QJ3f
sTdu/10QLLlyf34d5MXwuouBCXh/9CdnVtGGRxdtndMkqTIlbFr0A5kqpxhcQU0sUxd+9A5+0YKJ
qeXH+WXycMR9uMcne1FIhUxGIXboR3zKQrfkVvXcV5zWZaVvDwyUN3ZKa2eO2g/KdfNY9vApahA5
mIOMg0f9Ig1XKd2cpWYU9YmHLn3KPhDXN3E80bcFYwe4FASaSQshJivlefy5d0FZrEf3zdKmPATO
Oar0Jg4AFK20NwsXv4HQfq96ci63gr+h4pZBBWeQX6200y4ZHXm0tBWuV7H9KLNx5KyEkK4s1evZ
9LF3PsXT9fN+cd2ICY/k88aV8r+RAUhho2UtEXM7L1l+2JSBzHnG7ztS/SjObBfeGw6G/kAvXrqI
tJ1qK2+lbZASEqdJpYiaZgnFDb9EvlC/dSM1nRJyOf7f5wm2h9c5p0b8G91yIBVN6uUj5QjuIi2A
AOSfLaziBYPG+km6aPKzDtlC+av/ATnZgDl2j/zhxFvQ/4Z/vuRDUJ41sILWE9ob6/SibRCa5s7t
oRWHrNtJ3/d33rAR5HbuLJjeFHXzNorJ9AuZlk0KkpJ0NH33cqS/lTTv9Zxs5CwOyzyygccMJt8e
ZxWDD75FFgQ6FZycGyvKFgPMe/mka8DavA3FQi0me308KRczYydNT4wvhYtZPOUZt2moDsWCMmsD
mgMI//Vqt1wFrW7t2YbTF5GKhXgKPm1Nsp9HMju9HATd+bGlBjMtPMV/Q6canr7IXSOQqo3raXon
uRR6bPJTjM12hcNhPbfPASMjaoGADCOWKUxhpjLgKgT+iotJ7d2DpwButs9xY9GNQ5i/2/7VFiN9
V4yspzOUzUYApRJ5SEhqU8a0qd7bqFjvxFGmzfs94b+FwmAiuvCJQmkAZh4WpxBsv5ZzbaLHGXA1
RYEDtwVJY227ojFobRcmsxqCHsQz+vlFYTvTa9FJc01eJZQYEX5S1QMFRLfgqnSx+oD/ojKiWdZ3
1OOTwrCsakzQY/rR25sebRBq4wLzi7v5KxJ58tER4ROhZR4A0jqPDgDNmZ80O3W2t13w86rxa0Ol
9Xlrc5kAUqig/i+OkaDiXyG/GsR+Pknt5jSlviXYwttPBx/OKgzuicaY3I+Kw8UXS91sxHW1QEWt
rsKevzl1iHZXzEiFaa2W3Ixk69qlJqVHCqCODtgp0qUFHAZJMKxCn/A5ZElE+Fg21Bc1u9nRuOMD
BO+WJO4K75RUkUqa3CEl9cqsEkHnBtsW+efwnVweUmiOG/XblDf330Tqha8Ms7BFssw+fKTQ6A7y
TLwfmBzmJthoteg4hhUyevAPGmR3nTwyrfYkkuDEB78KdzCVpl+ZssE7av72qgde2DHPzZ4Mhbg3
kdI4OHr9Z4XG9c9XRFg0oWsiaHMZt+Y8kbSy6SXyopfYBS5V2YK7481JThuigoSgutWOP/y9ujml
dm2WfGaMJecNQCPoGNzH6/nZxCzymVIL3phVXL7lw567XBzp3aM/DhAZrabRgyRNH5FP1tgG+Mqu
0CDEx8N373TTY4SbVXWHRQhM/C1eOa/u1EFX045bca4+uOf9qNMp1lSKPpSOSE/BK1OP2GGllG8n
gzPaxieldPzguScWul5BQ59V3h9XPgQ4MnVGhPXfhq1pKLsFjwmLfaNHGIQ1jq6CqqZJ8gfxbH3g
eJtDj9/M2mZoDjZ/G4Qa1Y/jbDl6kzGRJCck+eDznv3jo6uOmTcj+jBK9kX72UJBRPJumGl+VRqg
H6MooKwhZKre7Z1AZqj+EglY2afv2q4ZtX08d0bby1jXtcfWUVegppbeWqb5QenxH4M2zNOr8qOz
YCDPU54cOqdFLv75iQ3Bb+W1/8LUzrr0MHGOSoihQFEOhWXaMoyZbpbJenq5M2TLMP3h5adXUi8m
rKya+cAvkCntJUY4vQ4cgU2BLozFMQTGjArimDmibW8XHgOuCyWsvSt+JQBbr8CHMSLLXaT/ORFQ
Gm4xTgIJV4DXozYMufTE2ciRl/X2nC5smxHh7nxHhuJmQhNQnHHWfJumb40w08mqCo4vbap/JHbE
enSTHrBOnTk8OJyoPPPdaDkD8fTTKnorH6EuYw/2KWHrQb6nybr7nLZyU5Na7wYEtmY8MJyiUgiH
VbUatum3Ae9HCPnd4QRkotOatW0DvbOD/ojWqw2krIYhmyRoPaYXx5nwS+rfjCyQLLfmsnFlY+j0
0EzI0NXeYc5HarxScQtR/3WEifEzxls0w9SCfElX0SXx2FmNxef2iU63KvsLuUPnDTsioge11IJL
v50RMIDesb7LhBXQLNTENnkBjlHYV8IMAGSRADKe1TQM3VpEx5Opd7k46rAGsZgeYCAva0UJm6W7
MmWn8dcLGkYmr1DWPcJZS8L2PFkp5PIv/pp//oN90SuEy9cFvdwbArFnKvAbY4BGVXRuZbbYcRwO
F6BfEwTf3vxHnix/Eng0JVHbcJBQQ9WmFhzGJrMIltcjeZ0j6m9ch8x/bUJuRI5rYlI1v9f9xrGd
UNE46OaEClj7vP3DRvVApkCqDjNHetW7q1CXNkMEH+RjfPCC8GK9l1tGN9A3Jf1aLvP89MIduuyV
7Vr3+LHiP+k9Vif6doVnEym0mP6hkyj5kCdDfWU7alzcXdJLSzftIIuPrYsY3OplA5mT+Oou9ZOQ
OoWsr2/+P6V1jzxD3zMe4Q3QsSIeUR2lnnUE2MscS83eMx4kkrrQ1AhISeVURhMkitX8thkT9G+U
BjKbiNp3R5a0H+KcmsgvCoIORD1WtIvtJGsLmfbER+b9SqM+Ad82bytS9mNeywOe7AHAuAdku3ad
nh7ka05V4X8rZkiOzRBU2Bj0+oAg0y4HO3tzBuHHERE7dti0eucUXtxGh3g3geromvdege/OTcdH
1KpXt5xJVHGiJARrZDO2JqqK+6OgpU25uZvHP3W7+oY7punS7FAq1rsyA9ouTHzG/eKxJjchxMdV
34FtpXlDPI42+74ZJintcOeUoVRKFXChoaJ97xevkapppLJgwganSwkuSh+RAQhes2tOcum+FJZb
dSY9YmXYKoTZcVLs079cYxRhuhWFI9E82luCO1AaTHmFvez2WpYowVlO8i5wh6s817qbFOevJsRS
ZiuibtqsQTj0c28f74kL7M4sUkHeO8GofV+/N8VmZnadxqqLlzBXL4OUXCZ+G0trx2utt7ajsq09
7V+LLhMbCJIVe92PLUPSkedKLHqt1t4n67z7/BXO7cDNwiP2tcwhYrcnjTj4iThx38XRHdB+Fg+j
KIBQqborqyClUgaAVMkzb91Nfgc+Rdy9HbauqDwsX5Inm+VYC6zxVW+3Vwzl+iInayzeTTKJ5EOa
hQEVxK2h5LgnGtc2++Q4E6wL2HObLC08uMGfJt3V6fh4pDjmGjePIAxH6U7A1uVL7W++CLvpme/C
wrC6ROdD1C0i0XX8Bb4y4aBNjC9ae1Lcni67XqX/P1F9lbBQiI8hjkkkh9jfjxg1vlOsBpwDtSIP
owQmZlUlwIKbf1HU6N05mr6agTvT2i8ilWOSpzloze88jHu1ckZ+oEJRfcuCbnZpFUknDeQB8iEf
hkjtLrPwrOOlvVL8eRd7gkuOEpGWgqiEW/476uS2pLBq+8tGvDFrG0CWIG8g5PlrKj6sMh8GQRxP
YWgfeUBFqsN1oGcxwb6sFFcmrQlmXpYOKUrQII3tX5qyzEkDOea+pYydoFCwMJfSbm0Egi4X04s9
Scu1V9+ycyL7HY0TIdOSuAR/szre55wXW7OSZSGRtjfT+PMJ6hutSeIpp4rb5XNsVM+m74ns58Mc
brmnB46mOEjOEZNIkMmo9kWNd3P0T8NEMHgvKASkzm9lKwGEl7I5Nj6kaFLxgtXJxmp8KzcNFaGW
LwrybZzuQem6QK/PYDAY+Sf7wAVvXGySFpJIKHGtx1mIdCJg2BGESQXR7ONlL8Uhr8/PNyngEaVG
yzw8DuGgOEfmJdUVPdSPqd7xI++E57b3IFeZoyPTgycvVxIeIzAPy4R6Kv43Ns+8gIqa8T2VpFo6
PNvhuF9k3/td0b0zuYDlf7eqZSKDPJiQTIGSb+7mQQw6YE0GT/v0WZiHGOmzkSov2iz4VQavTAjN
QGULJjiHHn4i3gNr2gLl1Q0SjioH38tV2NGDmOsIuzwxoXxiwavyf1vxnBDdkBl9DAGxYpdV6lF7
b2/rEguhyHYc5VccK9nSDfYg0qNoZGs0buC/rL7//7p8x8yiFW0w6x7ZKDfaUUJGJFJxc0lDnP/q
T/q6aTJTEFYvFGnIU6um/tKJimXYls4astFZTpmIoy9MOdWUnFjfWlKrYsNqYXkOUPPwCixBXFiX
tgEJ397Co76tVVAwqC5iRXIAofrbYAbGCcWV0MV6zvQbC1JOX3IizCNKIUtGtILJxqcvguI6f3/U
W3xb3BurN0JKlGNtyhyy9RrAUqAwBL2hqx4X9tMciTfvhu+sfHgJT7sCIGzYC9u+UdcHRKeae2/A
w51p/iRYEHAQmIB1p7TySLagiznGo1v4DyuRANZu00JDHAPP6WeCl5RUSwky0q/u6ttdu+bMIKuq
C9cT6rNEsUnKK6GwrkbWcD3h6XSk+OEvKvu/BVvdJ7eN9EXbGKpncJF5Jj34TGOlmmZHDLwBJYHM
olCeMxKQMwVxiEwQkYOwyTz7mPTrnoPR/gGXvYCqMWgyf9sD8r8/68ggogAMI5f/Gx8ca0KYu6u7
xkVp4/rSxn29oTvTG8X85+TvB4RGCHDPM6CLg94x4IOczEAYamg+KNZQ1/R9Rf89a6eV8zTRSsiE
0fM2FUI/3C+P59zdg70Ja1mucMPYjNSA9dWqi2bwHNgvaM7qbW9FWK/nLMSWpWT3AhOynd/fgeUf
dWKF+2y2jW8bMWdbtCTYK6IcNmXYncklq8Eo69xs8P/TKWY74NJmqeIZCbT8EXyerS78nEs12Am0
oTE+EAEURfa892Gc+ukBu6bB5pkXoZVmXSYoNB5leM7FrXTsZRLQrbJh1jJtYUq+a2CHfzXS0OuB
JJ6vIGP5szDRwNlRB89pW5aOE3QwXq2QjP8QhrqrzGztFGbsMkPNKiCvZv94beYE6AXEfZPf4wHy
O2qugO0GE8gm4SWlUWEIi+g3+pAYBd2dVaqsDaXXGLKKQYszRp9ZIN7mTyWVvg2uLNp9JvVpezA0
WU5QqB7XKL5XKqBrjbQb4/DiCzVmsoPXBhISR7Kdi+SaakWU3QGd+ykUhqalP24p2iz6vA5q6+bf
OrmoiuQuR7VJxH7qoX2elLDp3rcAHvO9kFjXq9K1pO61ux2i5q0Gkye+KW4CZynW2kUXyPraurR2
uqr6PpaLAp5C6kWUK5XA0z/i/pwYQNVM5bVWSCduNdwufAOTJij6UvYwD3OcQl7MEHb0fB3vypxX
ga2FUmRxsRycgaK6Fu7AnTT9R0Cv4S04ioJuejzTe5VeQXqlDLs63lDYqQAgeGto7z4a9wAeNIHj
CiUufg4+YzUqO66ntR06ylrCoe3pUHc3MR/UbDbJBXAX7s+kVbSAPHU1cJA55nQBuGJb+wx43COj
5wflpLQjeBbP+epiBvNBTDZxIcBv7V4u3BohpDpOzbiU7wXcIQZss9KkLUM5a/uswvQEzBALCU+S
dAVQFRuaMekgzP7pN8DKU5H6fgZvFjgkXjg0y9rhzci55y1PRyGOe8EZukC3kqJvR4rBaPsO4xSq
9tErBB6fqJQwaHByrhVRR3JRlCeWhqBTipIBhZ6JTboFMQ4aPs9LpobPpAjavTINqYEJFlhmh5GL
SuL1vWGZeIYLskAX/ly1AwBV3WsmEG2bnW5FCCARj5l1zt0G9IboALgfYqqxjiODMzrK+xVth7t7
bi15oNuYT0wLh9/ODcTLEIdECMzIcF1uTUsLItCFSq2Iuy0hTrrxdp7nabeZ5mgdmtVvXVlgPKnx
ywc/oU1KeGdfHZP9+kUwGnXwYZPqW65UlTYWy7bgDO2pq36YD3q4GMEXP3s5a271cvlB/9cODcPZ
oCWIfuauFeacl59MpdjQwnwDhnUxuu/VQ7wn6sbOBx1qC3DVV32i7lZwEcgDSWW4e23l8GMdlCVV
mdyBc0r0HAcVIpmx8t5jzDSAhHrjCh//aFrbU432WPzUNC+/M7S4ifWAn3Pd090e52t8bLLHA+Jq
eINRg4wVhWO8Juzfg+0pV5wvBEUn0YUX+NQ4K2Dvuv1JdXz1iFNYuXkAf+l/APXMEGFRiitIGdAd
YT7vTgy2hl3J5hyAQiKwykWplaGpsqMA5G9qVs4n+C8bVSKXTR5wdMFjZrnN9KrNshV+Y25R9gUQ
S28wxF7hg9JPX+kctW+GO6TEpwB2WW2BGrOv0F5IGG0f5J9uLKr2nfSa/YIW3RdmBN0XOAqdWz3f
zEQDdMlX4wW6fgUlx65SuxqkVoZ6pKmlBGlxykD/W4GHNFUm1fzWrCh+C9FnnNuU5qgZWmNGgthS
mHwqng/JLN0o2fAQrRN0DibUPiZI46wr9q6kNzzwJ4sdeQDKs4Leg+xzBSmiDlp/D0HMN0OL07Gr
C0lLNwWmj6AjtGtqcZK51G4p3gbsHLi+wI1tbjC2QmiUY4qjICWF6dpYX3VpDimy0VNcj8g60sLz
KELtWNobEQisF8ouHQAEyPMz5PjFA6P6YoBMWaHsqyiHUsPWXSUmauunyCwtwcwvcDvRSINhBddp
zCxvc+SCu+2IP8L87/g8mq6dTCV/5o/Y/XDUJqzxUXZz34443nuIoFACN/UjvOZPbkCXPUnYuiOX
UQ4hXRan/X1JBDWMVh5KWhzZR1lNrKBizK9y7K53cu3xkmRzIiffCnM3H/pIaZxgsX9TD7OlRpj5
nb7L+76ElPLjmH6dtzJfctMUChqYphLZemqdg7ZAakLcws03g9v+IeN6Ds2NgwhIOJ/rIFF/YBoL
K/i7z+eZZRiqTGnK1yDoGPxVrTJQr3FZADv2lojKyyJVCfqRT/XWzW5oMi4zyjTBUNFJ8X7Hb996
q8vRNUAJerK3RP7UKAmHmJ4F5Y1krmATkvWzu5aBQsAJxqjxqs6pV525bSVpwq+0rnNA5dm48dXu
Mmjp2MNaj2TG9Asxl1VhMc4o0ML8jYG6Efbkp7C7JbDS5c+d1lU59Xy+LMDqJcAJe4AbSSIqO5oM
oNeob35uSbU1IxX6d12akZRRuDZEZ1gmtLj6mgyRSyrYh10fXbgj6AeX2TbgRFX7MsKFBbq67Y35
m4tPKvMyTrQoTEkc8jmk/jmbxc44I/xfhapkp3OlvnvrtFKBXy/JSTjdmGyznt7Y3SQIWCwR1+13
z3vgBdHEwzqhhR05+35liuDrQ6UwxxMxtk3RFIPpFDMJYewDjna296LrLmallD1cRvjDWvX2DwbX
ZhzYVJYcaymRooT4j6u6MpjgW4zZNsGOUYJalQz+REbW56kttLTvJqJFILZmkopa1U2n0p+UeWPX
bmfVgW5kDsKKhRDJtBLQPYdZIHNe66ff0L2Y61iHIukNBZJZZl8XCFFBrnrTFlDzYFzftdnqXR7v
k5Y2NHPF/dCy69BJjXG2PDecfOu6+JTOvXGUmRidJlMZDzNj2X9VeFwDYbUI0jKvde7f7OTv7WVU
xzBa6+47nfUGEcbdSdZaSJcMxweidx2JTet6DAXfRaQ9CLw0enV8XdLvafn3vEiJfGx/LJDOjzHR
rf4pgoDDpwCjyImxmLlXoTPfVxC3k6RHOUeBRrxOnMDVoFn+iJvWpSp+o0xvO90V72QTR/WZmX71
QdVoGxl5d6bkFGTmgxkUiEe/Ym7AlHYHbKDFAQ2vDSptPm3yAkCQDq3id7ZWdyARUha9MY/7b5KX
CIPP8xsh3gbMtkk8eG3wj9g9e+TVvJPlFUWYULG2Kb6fih0R9OlofknktkbB2uvYKT2FAyO0yfxt
z02xRQ5v6/GmOEldoGtSioVtvwtJcanXzJNnvHSGJ2mcHxmGWnTW3hgkzXBsiquTsCls+jZQjPt5
belOcRSAgmEA52dFsjDwFa59EepuYI7b6zYBdoQ3JIzaaI3UmfFm0Hv/qXflFdRWtw1BAYdEHG8c
KDJF7sLUjfwOuALiJYNuZFb3+BHAjX/XDiABqaiYashae0OmQ8I2zxZD8qzzmLST63djDb1IeHxV
YrHVK/UpeCXS3Qhe2n7MehdqqVQbEqbBGPyIC/bpIK2/dp7L21LNXDs6z388SOF/6k+oYrgt38yt
Is3+MkSJNk0c+bU/Vru+v++g4Wng8wjzUE+nIzGM7oP4025NO3y20e/6JLFlN6AY7k3qjeItF79h
Ir82kdmTn2Oy5Fck6HV3VltpunW3AQJRHpheCUrZEV+/g2bHZh14HxnMq3DOc4Q159dQzIyAiMyw
wqqQyRSudK3gv9UL1BtivZZfQyUYUvihLMEXSHBYFmPolYLmca3WoHyylRMIoxT1bwrHEXjsGiRY
zk1j/mpdoOQtQ1lMMApM8hVoD5RU1NoOGwlTlAK/bU9DMRsUAnTWBAD9/DoOU+cMUbaRxKgpHzxT
QEaZUVwskdwN2Bqf0XJXvpCH/L/qNRGYLxaKgNEwNfzg5P6L0LAxPq24MUJzLOdp5PULTxqwqbv8
NA9JUSy8YVARq3Ft37BsAsK8aILypmmU3NBee6DDCtEqWbi2a8qpfJLUPGkOKN8Rhn+DNIXsA7jg
dj1Qc7xZVKzAkPA7fVZY1rQCJZb3vwhtkXYNfiamt6cW1ZX+Z+XBUrFLZzl3qd1BeB/Yhq0NSpWP
Kg1OFOuh/TXOjeNyAi7Fxc+5dRI8oqiznCAd1cmX0yZDCwe6PyqqQcELeJdsdUkcFiJgYgularAO
zZnvnD1tloTcP8GKQI8Rkk+P5YJKUa4mmdaQ+SlFMMD2Ca/PxJbOT3MsdgW7rYplQntB5aRklydH
0bw63yTEXvHXZkKX//pXTscQies9SqbDyoBRerQ/ky29d+PzlUSXUGpZtWQMA6Rs4Xaf0veSxV48
EHI2uJ+DfsiMUHlASl/evwKDvZWOUXzKjB1P14WBpBg4nbaiN9c3jCmussMuL6Agz/9QixSl3wWL
ucY9JO/p3YYQyhyGwHu1XMR+bBG5oe/eav7JhpxIkOiyN02ufBNS5Fxpx4p7XqehfjL3d2iXb7jq
iYIMIO0TvD8foGSKPkPFDedVbpcRI+1xqNCdaDHE1g04URMVkszASkC6NgkSoRk8QWRiLOeHp/pN
6F7ZEdxV0kK+xilVsB3itqUyckW31XNDXm0hv6xXbzUoowAxWskAm0YH4KNRIhW1t3VGmZwlQdmc
6M4kCZmx9wTb4s/WQgLHuFU8i1m58Gazqqwjvc8wp+8BsMhj1NTae34zrF6NN/t2TtGLGgaZe9LO
SWmmjRqoLoitqgf9Dot/D4lEeKrr+UA0cNPL9Y5On9TsKrIPd1mlU4k115E05czHTzmb05kKVvNA
aCCbm1cxUDkY9UIIaPqLB0RG7ZZTwv+mus6ydm4LeZuXCvTNDk9DSS2dZ8N640oRDl3zHAyhYf0N
35gf6BcNukkmNdzCUPtehib2U0c5GYDBxtYgK4UMYPfp+PGrazv7+sp7P1McWqDwq6FDR8GVQHxU
Kb2eEugL0Ze3SDLwpmYdc4jZDgw9kri5tjgDx91mgguy/XF762oUiQq+b4QWJN6DIBQqsb42rb8v
BHD3oh8gDxaiEojVjKk7MflQjOlwkQrPBfgRBeyJplXE9FglBBIh13Kyxy5+HF6Hsko+/DRNCGMA
5xATSjH5Y9CoSmcbE0eukl7jFj9r68VdV39Sz+R+u6V1yiXPCQJOT0I4to1f9WK0TyGGXgL/fufO
xpmQWWBiQ+z+J26QXJJUfbC89VCUhWBJHtn2epLVovcMk33Y1tAjGUU93sVx3lHQI2lLm75VT0aP
1lfHB4nCGQFzfmVeMHfB2KXyynJmnam6jVwNrXgvZ0EwMmm8jquZklFONrJ4BTAL6M0G1mwnCyBZ
a0JwQiV7tjK2+mKqMKuH4FOTthaUB+FXgXXUDk+e06qRx5x0P65Yy7XSxAO6UqVdZSEtYEGFhJVN
gp0JHbZUr1hsxdAg+dtZNphsdKMwFgjxfE5CUUFEu7mMNv+xeykNpA0cYSNoiWuiH8XWn3ns1MRn
gzSGpotv3i+LC15lJWi/wumsjbFg9H+2uAYXbDu82veGx7FO03PFztWhqjFOGbw1Lxd5/K4wj2nG
bijUzDIWuqlKhz4QVCMHFLwEyh/yl6mjoF3D1clksFVr9CQSENue9OxPGfHcUYcGXMn3E5IMUna2
d8gmm9UeuVrZTlXZtiNvSXFWLKfaVH5ts3CPPh0jyiRoJEGkGp87ve8RQBPWyQOsdfIYtcVP4AcU
hu9b/MWapTt2aCrhDt74JjDuRWjf1VzNTsEYD+8OiLNGlkv+JLaVALqOhGBlAKd2JYKdI3q1zXlX
3MjhX02wapDoQsvBl7xygF6dkobyOEWLcrKFXGwEAdS/w6oBhPRMF+BmijWz7dhYPJ1iBbyI1aDt
NSWnUhRFHPlJaHzdra9TKwZ4GY0S9kc94U2YK2rQMiO46iAVN/vxnFIebnys8EGxNUDQ8hHlSv/D
wxTUooupOkcTLh7tGeTSeTxW5g/b8WBFOqho3kRh2VdZFZqY4vWVrwamtjyCsaE1AWg4SbL8W6wT
Do9xDE1VqIWYNReQf9Pqji6w5KGO0PwJrGpL8vg30p2SQCglhZ3KRl09khj1WMH0iUwpaX577+J0
VKwh2nL8/2FT7Qr0YAeyBqYwy/UPrdYzcydmxunkRqpz6ssNYm9Qc8vwhS9xTLrf4+OuZb3MuyQc
yBSR7DdP6IgyKaAzZieCPdj6fizza/hTLYhVTbwmFXVQ3hI/zspfoaIGSf8GDWNJP8kfvyvh5z+S
6+auYvjiNzjMr6VXwBePsGCBEuo6ZlEuFVYW2lPcM243/DW8o3AwUdAPLYtg4TFz93oljw1MUyEu
SEI1uR8GoO0MHkYwohZIWXMKv7DfiATAIoI0uqbkbUDeudlOTaVXrcR5TX++bfHLzmXJLbxbxbw/
b0ot86SE0TmcWmvGM7gEYKwZRjXqVeOgIsGBvp+h8pq1J2LvZOIRNxpPbTW3Vga43u+JA3Y7zvWQ
wv2PFq5tKLVyKJvO7IDYMCn1hZH+cwereZKTlj3gbtnfUu1mAB+VwwSh4fqWWqt0bI/wOJKtS4B0
HS61Pq8GpTpQWy7yuORmq10CqZTJ/ZuyJshidRVx3b/LlAkfKtFtMheJwZ8TJ3mQeE+cqkaT75di
PmIOCp5PQCaJytSSkhL6wNaWQfH4YJ8aUh7B3xjwSqeLT0yd8gSsGB/bB0kn7GzD/HxmB7gIsSt8
RPwxBhPCkLnGrEVsW+ERghLZXTJlhv86/kyAZ1cxM+g5mHR2IR4KxMsfCcTUSH8KuTztxWETQ0mF
phYWsgXH3QrDnubjwFQVNSCV+7X/SjHmqJhfDt8BxHhTBpLYkyXA2Dsr1fh1QYIlT6T5+tDGsftQ
G/elM/+Z4nY+u4qEXeroCzJhaONK4e2qiIyCcPH+fWcD9dX+r43MgvMA46z1kC5ta7VIuz7JAG2i
lVRRUKIiaM2vhpgwtGENDwW3gCRJ95Jznu95fa9QSN5cd5NcFcjcA6m5mSoyB6ImUrPCXZNXk9iS
o2FT8lsIEYvhyBepyCeZZ28v2YVtZpA50qUJKcEJyUS+n4tXFGvfjdVC2p+dzFRK+m7TPd1BEPW5
0mQHBV/LHgvu5VG4cvRduxIx6Dq95/pR3G2+0gfd9AOOs5mpoQVO32SXXpioFd0rOmep1FlKRSxl
4TH6LdCTHf2aKaX3HBHAnC7mSyvjBNz6N2wU06F0lQFsTbr1o8p5D1EBloFr/7V0LTYrBIyecU3k
fELJfWIINlMWyDWOQ+2/653sn9qLd0pXWyH/BxvneVZtB+DitfbPfmD4nFL0LIRdBk5Za2X84R5p
zSonoKBf6tIrf44HHetanfjkI0FXl+hTzFdINNJGcci3TwE0IMWssButo+bpyMk1aJIOOMCVo++o
5tJiUOuN6+5D1lIdottvSyTK98XouyqKIjqKyoJnXq6bXnjZPssPg1xpUlGa+8tCLJoepAgLJr91
V00rVDM+m2wtU3jozyaovEwXZk9PDlbdCskypCQSElV+/GoSbuqa+Ca6WKWsaeAHW8bdy8IXrxFa
O3/92DS4MqqPdktVzJc48xmKW1/58Pdr7b1J1vZXfONjynN9B/l/hYcZFpEw/jfY31G1NtuqUvza
I1D6VOSUBFoPDdNyzQ2l3JqK7GsUnmXIGm55b7tdxYIWATJUmG2KHOzcNxmqiajkOhzHe1qJ2dER
U17ujIZvqBHinr8NbIJNCt7alJwt7ukN59CiURh4dbri6Mv1asOYlGZq7TxLjTEowvn1sIB46Aic
BgFxAVpLchv+2qao3RuO/dkSoG6ReWggaAdRHsBvTpl/0p0fx7sdyzQ8h4G6vn5AaIHwFxOToBnW
z5JZ7bSm/W7RD9gf/sQatjRTWFwrhnYVl0jOK9KsKr6xNhNhvg0EVcu2jw7x3yKiHWNv4IZl8jmp
ToodUY2mW2CTxsigZAZmBtON+TzLRufMEubVsFhlulG7RNFqiX5rMrBT7FCEqfjjymoU3uSMBPqW
jFSCDPy2BsHtXzb8YbAs12ecZ43x644JYGLjn5pJyJca7hKtc9dKsvhHj8sz+Y0a0d0+pmpZSUkS
sL9F5iVLZYHlOZttQMUpG23sDVyFNi0Ju7ZCf/HU5w6A1kGe0Xbr4CZckyqWjdsSOXNqWH50TEqE
yfKXTaWgk+Sys8sQl7vgzFJDRsINUSnrQanRfRwD76zP5DSF+0DKdi5qx0hzeyyQqTSuBtV+yPsc
I/pP9e0+ViuRCWfxxi46YeQqHUMYXhs0o4Y7PnWYBZnSeIw0mJHSdCHiPh1EzmAtCDdhZfTOmIPc
2D1ySqOAzNCRCyPxkeYbL0mK06r05MFetKpc9DD1Eyvp9EvLGC/X7fZvG7OLuA41iH7/yjrzIpzh
yDHtqik5sNVN1XGnpd0vH15VJuI8vYmXH14Ppbvjpm6y1gaMK3e7RKKjrYkLL5dBJ+alB8k4z2Ms
x9KlXjLuKx39wvW9SeJ1u9LqB4kpRYHpUbgug2DtCxrY/3lbaV057U+buXdV83fzJqPhtAdk6197
NyZBB1QtReYccBD3lJ8rKMOWSsApQOQnOMUhxBj+Yfnh+jOP/RXvzWctYQ/PTUkgCaUBHrRsGH16
y5t9gIG5cc1fRvGjq1+WixnfKlk3IwQNkF3eeoFExheCrhegnSdEH2XdPd+KRzvT3XF5DjOdaTfJ
Oeaonem2FdAuNEVFAS7YwpXnmKE/F4Vi4gKp1jNCW2YYAeYoxcreiVyiujAWdrC5ksIjtTlr+TgX
BWmHaXMwrr+05+zodidlJKeTvIYvU+m7ARUqMulVMP5upgAl+O7phhqDw19mtjpo0iVe0HASnblb
lMOTCm+wVxTOLg84itkqzyIJZq7cSZ5NBbUhPnZpIdOEO0IFj/XOl81lOra392D1Pgw5cYpvwkVM
pjYCx7Gmn18zN7MDwTc7LAz7FyKyx/AK+z1k5mB+5NoJn+k1lFVOHEBun7yPQEwIu5P8tp1QLqoD
bdOAy2JQQhRngSFoMuAVwSLuKx9DuUnox6wfn/0VxyBsOLwKW1fi/fJeAmdSS9t7tgXzcP7HFPxF
spXj6oQSbufpDscY4QhGncW85gxEUPjal7+YSOgJgKWGzk1TR75xEFqHtTmUuvo1ZRezAk2r3G1X
Fww+g+QFQWeIXQRDE/0w+dtr5H4hLLPC8Qu7ZQx7ggPjcoTeO+lM2Tty/GoijuL0rFWh9TTHXkRx
BW5W8EDkWG4bUL6EK/UppOiSGQenTEQc0hpS2p9tTNlOCLHahLemdk5DqcE8lrXmhOrs0f8OCqx5
Gtvs6yHPn3flBImKh0JW2wUeHnWwb0KjD048/gyriIh+NeaEh+3G1kbruyIzGspt1zK9i0Ky9j+P
KF74A+1kI2GAFU0asdn5QD8xttPDoy7vuUv8HPL8Cp79yg6joLeTPtM9Bdh4/b+hV20/f/upw8Wp
nHZgsHJWp4qzBaoMpvbMF5fzzU7Qo3SZoLsIBg/QZr5bU6o4P2NvVb6t0u3lzHkYavrN/wRasdIy
RRhjdsQopWhIEMzL3VxUe4wTabMVP5SbIah1jJgj7asXkmKvqu5qOBi09eXiOHkqFTtaXrjSz8so
D//3VmprIDf5ZBLNF/RyN2VdZvNdqG9YYmQ599oHnuVJGLpdkvjJ7vxSKtHLHriRyQ+cvpgOV2J4
ipnf6w3dMevsHFPLKrhlnFmCmNUgIFyylc5WREHtyBMYzZD8tgBh9ciMW1Xr7tQzagnYwJZFObIs
L7Z6Fk0SJne2RzNqqru5FiwiZZnfXCDlx3JT0qkTBBIztKov82J4Da0raA7rhTmY6Vgxy76WoN5L
H/SkzAYbxSunyfj8dD5E/yMq3EjpdODfNKOvSyzEtTqvIO0nyoR5t4VzzIF9P/BM6wqufV58WRO5
wmjrJT4N/+Ez537TDFAfL7QA1ERn26Zy3JPBXDBxyJC04N6VYHdaWSw8oa59F4Fq17iZWPdkRjW5
lwYLqXz/bCO6NNjlrNQAThWe8gTJzMRB/ip0JFhx6HjsDv0RKKPSOQMFIfsQz6ZLhO9WIQW7xukw
+omlOgzJNPXEGMJd6HAfIf7DOPeTHqTR4IRHh/ZYEN5UFhRoIK/4jGmhqlne7I74jOGiS2y8XAZP
HAlpGO1brkOyTgOxDvBveVyaLu1IO0NTUXka2mE5NR1rNQQmyFqTRL2vLf5CkmbibIVWJ+zOIwHk
3j8OjuqtUUgoW7HUyR6VYUkedisiKEttXN32Wh8D++84A2KuPvtSVifq+eY3mnnaUsH/fcWsYULJ
55qOtgY8UpjxaoK31tej4+bzC7iRNJR8x8cCeU1lmpz7lddDOs7uOqEpF/9m6snqCAfVM48+4mVS
R1lvLfjJ7V9LPz2q8EhKx/wxjZS/m5jEo/Tsv9HWcUyzqrTTpY+CAwRlC6hGaL7wC8HjI2ayO8XI
lLQ9K2n8xxSrPcaxpWiex4Nx7aLiUhui3VTTj1/Ej/2z/H0/Yohv+zj6AJ8vnATCCWGIQmFhi4OV
fAsjpJU1hGEtnuolzQSJti/P97/Wbs7v/OVJyW+TDcYRrFVie+aATQMu8yw5iEM44h3gwsCPZhIw
BGXy5N3JHFebEHSinvbjXlbo/SGsgNSSOaBsXnokN0RlirKro7NgieeHYUSDH9fNFM9unJaIg3n8
aYjOCmQR0/aN2eZXPyyN6Zptu6Y7f2qYqEhyTWe058p8SAjxAnHJ/gY6tOzcoJMeVxxnYaJ/G4a8
iMQSON6dcxR4h2CGRgy5LVM5qW0Pq0KAlOMPSm4rRVVA0N9DO/m9rREF3QBVvpmGlT9SJiW1d6vM
AzWA8F+PzWiTvwWEVMZ1sRextV0IGFS4hiE2qtMlzGudEWdI1vvgWUuisg3s/58vSujhWbIM4Y90
euFyDMAnTtTijdDYoOP/h3zboOmKOPwzV4OSudeyDqtoLESZiz/r9zt7IVidwEjUbLL0NVqONbzY
vu8F7P4inuSj+Ihaa1uMBjrpT6uBEdOrzRupu/cP2F2Nn+UvcgGqySO8u/I+OMbh7Yj7cs7na2Fr
7Fg9LAUJH9suacIGZwCwwhH34lUFyyxjuHImgIZ96G8anygUhVeVP27mWh7U1fsYfIdTrRhltsq+
n+gTNLI5pmfHgNxvpIVq7BJDU+B7NLJpJvx87ynN48eKQMekQrDYHOLQy3dLN6eMBe0AfaBFKs69
EOje/H1A/dvFfHKjI8UgsoQILMpajqooQHBYX5TOP5FH7ZN2JHRkEyjf2mowHJM45wxYfIQFsp7a
ouIzi2k6XmEDijK/7dQ/ocBg6Hy908n6RWpzEdzRYbla2SS9o1hqIZ5Zz05b/1xTplznKTHko0sW
jWsSrv3IE56oXcF65SbrJtsbafIiklE0L6e8xV+PATSd90JFT/WHNCDU5uL8UdxyOoAUwZl4NHDW
MS2fMS2/tQNW10GsLaimF/RwiQvqxl39DODwAoioZmDNAvTinWZdCOQ232O00EVcGjs3J/ex369/
64SBoCsXaiQCPRidAg4cEIPJWL/7zPRClcPKdQwmy0ZbxkRK0uJ8azxCSYi/oSH1wWRDIyzr4vFO
KmqIN0vSn3Yg+LYsee0BkoMGG6NSEwcrY9Ep7+qU6LCM/LA8ov8EMyHZKPX3iBOPASXJECOv2/dk
UKTEE2NNE6SOIANgd6qd/RZiLT8gCMyIOITRPabKMUoLw1htgE0GttoQhAj9+k4i4KIDnDCaCbww
jAl4i9TcG6C5cq/krUn6cNbpaghY41HClX1moCPthePw1tt8/mkLsL7qBQMYEx2J6k7lLc/QT4h5
KCeRjiw4NcyEsF7Z3ltBz347zlW5Pf7fPYFAPFEgiumzJLw6WshPN5F8cFtvKGhw40t6cTD7KpgU
h8aKBMajzz5GULWbjrTA1y9BygGTnAxRAArPAofUuz7MoIBEpQ37PP+GDzIjzRhmHrLErbnVNTLq
NptEcpix6bnn6DaB72NsrFBsgNMTETJ9OYSBubBGL3fI2C40k0lZLcpK8bAjPwhrm98HN7izZTEB
FurkKS6WXghj5cq/QUvaEOEGe50YFvm7AKfxHGvMKwzIVk/TvUTPagjqfNH5ArNif17svjnZHvls
8CcQNJ8U/EWkJgUIRQXNtTiBs+kJHsKmKbzJBxwLgu6KdY1aZDeC7LlXpRF4nm70HYZZm9lu6zRZ
kFZfcrwtoVgOmo+RXuOgcd0x8103VykqT6Kh/tH2YHZTlLzThL/t42J7sPcX584zQ+9UJQXWZIq6
AcC1+UGfAw47s/3lO7azdDlw3EGl/AXdteTF/84Dbenoz65Xdgc6BkmMs5tAi/z7U65PISk7DJgD
lOrdAiJBuCrsOcyeELtCSt+V2Am8g1KJF0cFc933vnOc0kiJCHYaCfyZT3JvfLFfqrnOMp7n0Tkj
QOpkZZG+nc7BrM1mXVEIQsJ3sZftj2z/sG84BlA55TB+4wEC1OqHtWsjc7L1HEYDaMqZUY12fO7q
Y+P8oKLO/b/vAiq/nMyEeYKc8hrmp92xMPV5LlGKyCFzaz08vg1WaEGxMYcwRvgQdeySK+MlkrSG
tGS8SzSl9YQzkvnzErnyZkiBNURTtJhUTE4YzhUyqSLW2LqATMiTEc04oOfNpzYHffOlKRv7BXEe
gf5upHWA1haVMCpDv/kx4uin0ptmAmj3te44ALulYIYVAe2Hlc0DEN9RKtBafWJ1EJDEEqAcAP+a
aQjCq2zIEtMWuRAR1+ASheLwrfrCnp7sTFcNw+fP9R5P+GnajvLDIiysuUEB0C9I3Z0cgw5yIBhD
nkPdyU3MUxq1g2mEruq7I4bRsrEGXqQ3+CYuwQ4TUGYFF8VAvao2FFoBSsiJfcl/DGMyX90MB0l3
QLipe4aLhsVkxgDXZ9sF3mw57brJCG8IOnVQCECDFAkZeu6ONKlYt/FN3zXykpaF1J1P6FOej2sr
xWT7yx2666zlCO8GmRTHCVG3QEAQYMsie9TNLBvGA72l3Ve3oF7Got+R3zkRJrBhkPCb9pAkF2v0
IteKMMbsU84FUa0ypQ6so4r4rcf/ZqH6oJGaW1YslFXp0FTyZP/mH4Uxc2y3UshLc2LUdAwM8suA
6rey3hOws7dbMB+2a7lfrquubBexZSDcADD9zuho8M9B/2+ykDZrzg0BYNGCciJiMEC45fGF2mQi
nMZ9aauKux/53cjQY98peUQNyvyezhE/Efsyc2YN16DywxUZ3jKTShgndasLJ+1sBo9vbkXY9o/e
L5uQrkx58v9fiRvrJHxS0ARdlZaXWs+wrBeLkgT5AAnB5aJOlzwoe1QFGvrI53LeInhAtWTIZlc5
GksLZcdtCVkjyBtSb1k9SEAPlYnSVRQ4EOK4TmZfu5gBhCTOhP3+T3d5DQWYEJNMR2nzA0QKpAY/
DNGs8amNaQKrD3wFgOygs3aNr460Dcf7z66JdJ9a4Vy01f4gdc+BFJXxWyginrIzxQgrGhLMm9Q1
DGPZehr2aai09/G0Um2IQDOFNuVYKFzY1EhgwHAvJYpk9O7ZgiCYbnAlWsOrIeKqn3UiHV7e72jL
96520b2QdHKhLPkbG6NLbl+sQ48zBiBfkquOzAwdoCIs/mnrKLYH8NmGGsdKwG+CrzOdEW1qzUkb
XZFB/G+n1Z5a0dVt31ompHypih3IQiRIypewXRSIZ4Yi5q9DemZ1jCSMvK5UMXohFXTHrQfHvKM2
aEswR2ftpJe9tajQXwGQBpZ1hEcA1NLUtpsVO3vmCoNAclM4h9ESimeZ8PhfE5SQ+3GacdHlT9ON
gM+N5zk5CMIrEKmEp4B8yTeJKZTGz0NRxMchF5Avmh3ewDaLXzpOG1NjOC0cqC8/uD93ZgTFVoBe
j5zIm7QmdxiWeIveoRj5faYphvEasZe1hjnqnMvdde8BMOJK4mno0RFxA6Gql1+jr3B6KXeGz6E1
5+Pb2sQBFdSKDTocIlv//8zE7LJjpfU35cq0SVrxjVcAF2OORXxztQqIkmT2PGQgUbvlH3thWum0
DAEuEGmhgEmq5N9M1jYidlk0Z2MW7kZOoCv75w3YF3FeXz4LzVAHQFAwNZsRD0h+Hwe5DMgxZLP6
eo6qW0buIn7jqOizsCbNXZtaDszzooDXOrk5xd6P28Es/n7UrjeZDMy+LZbcsgKorc8DCeS/Q378
t86aWPawMpCYghflZp2s96dm0DnsvjrupbGqZgL/+bPelQNWfu9fYuPmus/IYb5v6gKhAwU+Qi1R
e649g3tUzigDISwEqEhnX9RO2REfasbN7VPP+mRuN+1nuKBoZJVGMDjeDYgX5UA+zIZLKUualDje
h12EkdFaUkaEJ7q6rJG2TcJxqWmywQnn/oxtgnLgtbUeE9LEdyfcukMt9I4oM25XC+MhPcwbxQ1B
LdvwByrcZbISQfXNvkzrQag9ErTk0x9ZL18vlrQYiwMjLCLf+lnit9dSGapmAdWeCwBzA08ppaYq
0/zp0/Bb1gzbTOYYF/l5ng5JAZSNwtPkD51TMBXjswQk1khLdwPMYpjdLkpp6iypso2boCW8qOFy
UhBsZ+pXdHz9suy6qrIHnMzM4iC2Oa3Mgb2Li5yc+o8JacXw2U7S1cjApOuwnANV7aumoRfgitjA
sLdqSH7yTomXKKirYJsZ5S986Xz8NoBt8WGN3reND69kfefXQy61t6EL+8TqjA4dbV8znN0WgjS4
qQroA1oYOf45EN+k/hKrCRKuu4LCatYrm9kNHijobdU18DLSdLUuFTVHKmphbBaLe0L1rkGmBpPr
s7lyK/iU/MLArdlwzzT1+Sv9P4l2vJET2Xjgngb0HloFanOcHs2wAopvSrSKTPrkX/oxcIYlDsKW
2HgS5d/qiNfdFVKMV94P/7njCNTWCqU5MDNoOWhB5qDve5hNOE1OE6fbUSE/SKc80A4Z5aGyfDE1
PilhU/GCqypgbgtcBlye3DN7jb3Q1APpajQW+oCrThLyUC71qVIEmKfhQBE+9uGWFFgxzHdBGSYE
PSRE5WK5yX0h98bttOftgSPRetto+pSrMVgpCWe59VAR4CyP6qxl/Sorjjm1BbyK5oQJdL20tuw7
GInVknM6N3M+GC0kZwaqyWDx7gtzmYTtQuKbRGXp6Y0e6U6bsjv8Xc2YR5gTQ3dCheHddBUkXqq5
NKkXhbVVtRUjDOeh+5UxE+sG0TxoDSs1AVHYLM2wYjfeTsZmJTnX5uInvnhoMgLCcGbiQNYjTeqE
Z4W+0LDyKvJZKp4Skxsm6hyqfo1+/yn421uHWxs1LS8/+QI7gy/AQ1+IYgFIVE0SpOkg6OKjUVmP
kg1riUkoCkat2LuutsO3zsPj6RM0s/EWALDJF6a94FTUOiW5YMxLwrXdwl0AUExBkggHRpO97Ji7
OxPDTxJXjdBi6nYfQs5IhMPlySTE6+0LdGMsjWe3bZUPGIATE5U3hEO6Mlgh7/D8v9IxvRPpAKH5
2tpEdhbbgTY7sG513xxcA70jwUOTJZ9i7WW0Ljicu8rDKGdgf2ySIS74ZoDimIcLPExRzfm+T/h2
OkUgWPUKOfWzIOWSMHWeLFZIpbtXN9d035XGri6S+T2PGkVkiE/TakvnXAo8FGcGm09LAwPabSuv
HGrTOXgPPpKbQzpQhEIrS/k+0YvjkJXs4KgPfVTJMnlZWAFgdtQRcULoXkxLvRw68mWFWu3vNPB1
Vl321feLCcoHjfTmODc5TsCNnFYMwBUuyFZLE2A55+F3PEUtavZ3k1l37ZcknHKLuLozN6kl5FWj
o5eJCcbhC0BhYiqSIm4WQAKCs8GKs5AhWzJ3cM96raDSWXp6S4W5w16vcZkP5ICuq0ZElUL6UsdZ
A/5KmgFspPYTcFetN0A+rWQvNufi8KXsWtNnYHXGHXngaxHrSmRWXo6LJKgFqATN289x63YHJPG/
b3It/P3/fL+uF1jq0ZTQCSJJZgrO/yjlXYL8mJSn4GvfR1+sc1eFQ0iRnP0Ms9WbZRM9UHJo7nq5
zScSqNQ53qoj1TeMGLtdoQq7q+lW+LDCG8gmlKDV/mkqMitO1XLM4x+fKSfi6IL60jpohcmKHcA/
2axW/5P6OyWV6RY57T8vSUFTq6NNjs0Nip97vrTMWlAoBZZpTZZaSNtZ7tJWAd8j+tvLzRnHgc5J
u/Vd/FbEQXufcafsH47ugmvhR+PbeLVdTNlKSTQF0M85Y9plh4ynpLofjef9Tz74VNRPOaRwqEWI
p3lT5nXMzuozstpn2meSw0ODGcQpzr+TIBnBGW5v2/9Nu3Ms9ySQM9IxW2lX4sjSUK6L1dujyniG
X9rCRG3gqhix2TyBgYIGljy9ngrk+fyR2K5x5NefwCfOOx5sbJBJ61m7B7qWTNHFwKTwpM8Ycpt3
ZMcEkSiS8RoHJxV+6kaR9pJYFNZWgevXGlzyZLIbYEXnsis0DNw0gtSyyxnWg5VuMVtqgLr6gkDJ
9GOWCVmY9Ugis78chhUlEHlHLd4ox/x258u2DkcKGpFyI2x4dDKSGjpZk4RM+ewZpfqmI1f9e/TD
dwcouDs5VCA1WLYV/NkY5PUUxsHUWupa1S3y8bwWeArklGlqw1Kzaj4czToJBCfAhm00ujaJfBmk
RWe7ha8DqSsDw6PSdcqxgvr/UyxOgGTPmBYQKFbdVVikTdlpZgYrPUYATSe8J91enXmCIUVs5OXu
YnV54XasMzcXyKJFzmHqS1uaZB8Q+6yYpT4pPpm78jWJt9QpBHdtWRH1aCcHPi4hcJ1UX9LdopVV
wxBb61/aSmfsfjKvTRjEU5Tkg9RV2OM0qMzD2AYMN/8IE/uo69vO75UbrZIsA8+WDn8o/ODGBPIs
n2cnINDvS0KtQHjghLGv75zQJJGBR4j8nOhfU04ZMLlAA+VI9dgUcgxzbzbg85IYAymwPQZnHguT
twrpS6cPLErZhoJvJORAK10g6P6Y5ON4ug+RjuxRRG3C7NA6+i/lAlgsi4mTSj5I+6efWNW0Ud+w
eVwJiJ7uPk75rmwB0IUUfGsfAhcbqMm8MLt6zsqCvdi40s5eAC+o37O+77mNgRwCmt67SYS6bs+B
VRNxFtNQns7rl8hCy16+19UnvhTek+IA+Th8Sz8VVKRAbtmYK05ssOLW5leaQ7GJoh9z1iMVFx+1
R1U98NsoP6fAYEitkhJv8nTxz1qxkoeYKgYTGiQYrG75fRTj3MeyaBsWiTje3Ldv+0Y9EJTj4BpE
OoOSB4pw+mZdXcNsJkOIhxwqJyJZLn9C+2zFKv903juANALzg45MieLKYEReiTUYu/VcpViRsuzE
DbyP2XjFOxbewzNEBFE/e6N/KE988aRPZwkAxu6oedC3tBRdWejn9hc4gWH4j8dxGIxFUCWm0Ml0
hFBi0fio0/yWGI5KU4cIBfY+G1a1ACMxbGG1vcCkUaRyiuPmmiGYmT5m8DibpL0ROHbENDh8rQuJ
HYRUs8wQPwpKIma86kbJo0EwinjRKaAfyEXeJkFzGGJj6YInaF64dpKaNpxgcGoKmbk9Edq+K/VV
pAVf/sg4FZppT54cllUtJsMjL8pEA076FRkouSVBQQ/uUPEmhb7LunD4xlKJfoxrrOY4M63dX1K8
lfe1sUyWX+l8h62e/a5rsuBTKdJHsFBxI3iMeE9s4bvbcYpdAJnMpb/OG9XU19+e6sYQGSJui/Jw
8WxrP9fBO7xuOmqokw7fK8Yz1sHmtV0mFVIoHa4J8MlpLaqOse77jD+rOe0dpWWA2oxcITjH18rL
8qObw912yrIFXnrcZjyDQ8M9bI3d8uDl2QXz4wNbOAya5k2HMgL5gF8TylYoL8l8SmPu6Cnhllya
9Wiy5ahrqhH55J3u8ObW5sJA0lN4usjmauzfyTFD7f3wLAMKIc6kf5rQ7JFJDyZY+62EXRUChNZt
q+92bZbw4gdjmrCbikfCuuTOqjranIGIRAgywR7A1UEbecji3V0W1MEMdL0hF0/3A5ySR1Nks5xY
BD8N18bTR5S9b9HFTrugOR/UmkFDkgFCke1xVY5G11O4+b7fDtXfJgKjsfgXKZ9ILp7XJX071lFb
ZuMbfQEEX54wljJaSQyVbCc7Q4qdfcUbGlyBc/ryoUvTLOOycPIwTl0R1yeFB5+pzxJHCUD0s7o/
WZAptwVoncm+tES6dTj3+FI4p0uHAWb8A+DWnEgWk+ktpMLWPdAX5IGsWTpw+PM882rV1DT/ze/X
qmYwxt0xw1FOJyGDN2Nea0EcRpwFwXRU62gIehB2FYLjOb7guCQba6iBFx1wXIyHEd0f01urRK9o
+oD1YFAOK2ajvrjdMkT7QVfLRF9qQ/rkEatT9xs7PBwv418Iz5JXIgiQcHUAGmoe8rRtLOwvBuSk
Z26qM8EyNHKpOWaJq1bF6w/MT/DpzVMb9xZlOBfJ28QX9eu67e47YQcg1Oap7HUfSZ8M+wdJkimb
Dgb8j1kM8TWIu/4oMJKKyBHvrw6mi1aArPVJQhoFd5cdl4K7KIxa5+mp/xS41raC0LeeCwiT6zwn
0dBlCOaUzaYr/X8gKy9a+fhYPZEbqK8QcHDAMjJqx2WgnPH5Vg64loK5fHP4ffXVfnfSg5IYhr0K
v+XxeZTIYJzcBYkYl/KhSq1mFbUXxnGXJTaJ7DJExNoNIALKlHfpVHURIYpea0XkTlE+NmjFbhdk
V6vqLa+2sPqnZqqJgdkuCdixqHmMvcqjdLiv/QgS8zyWtWXt96VZgy9wTUz/RUni4jSKpN6Z1p5l
wAX21UqpIeNVhNd9e9rKWEIMcLBf5SEvT/YQvQaEj2lE5fLNwtwNQBXMyhnXt5XUbPO1rPri1FMd
Hu0GYzfAybq3KAAjKz1hiLH3ha0nvDyo4Qv21iMBpK0CrNGIm+PLhhXne+lCeoz2mZTMd343jYI/
ZeHCXx+4y42HT6q4Ac9WMGKCTaVPuE+JbHVaApeGxN81ZaE+945bPIJKkrIxZLYWsCHhFMyn27Ci
l74PLPBTagqJpPRpFkrQnDU6KHHPMgnnEKLcwyKNqoKdXXFcFGlr78VtPPK3/zm3hIQEAKxG23ac
bHS/1Z6XHEaemq4pU/NL0DGafmmhNj+roE1E8xvtGQWBL/PfOcXsFTO/hKiH5toW1CsCgPi7nohA
i+aB2SZo0KxjQj6bSi25eB7ubh/lHQT9vW8SiIa3abSqaTwLtr6WoeDI2rv2kzkaJpDGqvsf+h4G
C04ioQO1npY8qy+yMhJgvLftKKlfmr7r92HXKg6EOGddwewAmnE6+YQFqU8rcbgGTy3sfJ4htgbM
d3Rl4M0+aRCb+LQ/W/UJu2ck8ujFG12GYGgK6bT+eSjcjBoEZFtrYfviTlwqBlGo9W8/1+apx6Fv
6I2fMFlJ1MUtnZ38xmfcVS5Z6aBCv7dkFUmOBSLuAXdS9AECBnWq6uV1HU7yMzznkkk+5fkjFBSc
Yf5hKrvb788m2aznIDMox59wvdU9SazVCUS79nwz5a7Jggxg5ggiQZ9+W/wzXFXmKCPDMV8h3p/i
Yy8PKEzSdW7iaB7IxlmLt9UEeC/rwS8us4A2PeSW/L1PDs7m7kXUdLTQ1xv3mYboETA2jYMNID9R
PJep0pLHHqfbwx8wP3xp6zzulNDCRLVpJCf/CXjzc/piI9X7pUJgrh5NqlKaTf6ablF5V2g7vLJe
F2Wt1/6JMHZNyJkplZsyvulsQgkYQG/y6DC5HqmbZnJSSFEoXDlOTZAwr/VjtP4X7YUUONs2eOzo
eVQ9CUXB6hv6x6KWZrL0v+pmn6nqWQYa5zLSZGVJ5EgjJBWtZ0RyjIf2ndVe9fICYUr26XCyi0As
WcW3/u3Hhwu2wVddQoTNdwivekYptNejAkq6IJhFy5paaSpnhbzRaLLX00vY2vZGqQ27drVTLUJW
PqSAugmdyYZCE5UwbL1L5n2/Wm2LqwMyVFPpgyVEvqIBMNmSJfsbLowh/JDhtLto/aB8egFd0jKE
3ROLiU0vNcLszZGGaQYW7s9j+WLlcG0sJZIHLqAgOAxFvSDeGvva+HzYMZMAXnxYETX0iz9UmLe1
DDYrrXdkzIHm6e23u3GEb4XUMrokVLgj+gbypeEOx0skzT9nlRLW0h7UP6HsCBwYW11q3bIEkWAF
0Mz9OquqRu381GQmv5QjpE84b50vOQNX/CJkgBzNeU2A3vkFI6CYXncsyyAQD0nlJvAonbEle8gw
8Vp/C1QHoYStRKg4yjqLjo+TF9yqrZpyC1e/EcbdTh8SfhuC3HU2YNGx5VxWXLWQPsDcmpJ709qK
KwwvuNcsw57VLjhQukJanwupKPFNuMBKU9sXN1ledg8MG4zMTJbJckPnu/3njOKUuVeY6X8XcmAE
U60buZvM2HqbS4xiugiU6WWHWOL8ymYYN4sMR5tKXth9924On9iZAqCT/WDXR5Gdd9xqLBevnVdT
44K7gyhLWGzJpb2H5d9m+shcJKfRddjzaMxw4owjuziUlAKB9xrfVNFzDhC2VLTN35kMX4FyS8Bd
uONwVdnhXmEH+sPFOudWvVX+6Z/BLzR1va8OSaWKs0S4f8Z0/GgIPuPybX746btVsxB1lGELsUvt
UPCx8oajq/pc2tWU0A23CRFt1GR3keMzUvkl7P0ZlZGUbKDyiHiEwx8cO9dZ7VguLHRAh/z6St6g
J8DmoKqOFRZyqyREwxzWhhRjOyiL5WOBajLOUwmzct1m5WvH+caLX6Pv1zmi+KKTcicJBL4uoHQ4
wjuJyWBu58CZYBv4hch7867xza5n0hhyvXog5m3Cwzwp5j7DxiSZELGXKOAVUbF1CGv7Ow6Rch+y
WV7Ab6zGw8eDWsrNkYlAADkK+PtvPG1bVYMERk4/cFGKBg9oUsLXUVfXIJWny4NOCpXSDq1qRZ9b
qrWdsE13GOeEVUyF79tHZLpe7oHAHPQLjaJp3y/nzqG0jixUmXKsn8ieVHGrw/1Rgxw6aSL6apMi
EpbIcUEe6o6w9SK9Tco/CYkeftlg3m9+tj2vUhvfDDXkiwjA0NvMZLgfERStcxZuh1zfAhKgAGIP
us4ftM2u4Fhq0ZIjg1yRK2qw0CDDtJTddjkw1uAmu6G3BqgQWzpS8h3ZNQj0c4lsKkA1vGaKfR+e
ukV1h17xmxzisBtFdNNtRtzu2MfYP0u9iNfkwDsYaFAwYSz49xzrgFpn4mikpahVE2gJwO9+UJcr
lADjry6/hNPzddKZ1gtHc4Ybn87gd62w/dHqpvzHwTWfGndxxq3D+fZiDg4QKNxuzAi4Zfy3sa+D
EM81gjMnHJD3F8ucvf1+9RkVAHfHOLaG+SlOm869dZJEGQG1NKzUFFnEaShXhEUk3Up5VctFgEgM
kdIRar2tX3gOmI3Kok0X4JbLvH2uL2jB+n6SlnhQvgNweWXAW9GejutpPILTVFBdQ0WUWzXKMDVO
pnntgAx0oqKUFHkvCGBab608prL1Y5Mq6IbOklMZVxzSFlZgNv9v9DyuhkO9TbKk+bNowDNXbhUB
c9SHse3LeU1cTq2YsoQBVaSaZZi1mJ7kOFZDPBIcBq6Km49vaf9wlYN+FysD+OROx7rpYvFW5LAM
N8fvG+C8wLgelA7wDQgi2F/EWzFmXQ3Mgah22H0WyBqnpWXz22dQAzqXB9WzV5eEPbMe9VfEN0RA
rkS6OQiEXd3cdtX47KSfQm/TH/kAAD8aEI5ZAy6UcuVM7vwB9b7teBdg8WFUKojgZ45H09Eq0+Pq
Ukn4RFONPcAeOYI+hOKaIx4wSE2mSGBioodlIGAzs/JKE3e4hTsWU/bVuc20j+sS7TmPVvxz4/8z
A+I+373gH6NumLDnJRnU3qlg9Wr/M2m3S5XSNKCHmYOaG9Mgv9mAlCMR6006MkkepIAqNVsOGR8U
ycNtOKWd6FT8IF4S5uC0kuT6newHWglbjC4Oovt/IufYj9upG6aLeyIS63lGxuNCZiuiNUUHIZFI
yxGKIXyWJ9KUIy17EVQqVNrCZ1KsVaMLCkmBXCzTUdQnFhFeNjyiykYn282y5k7mf2BxZzoMRm4l
kaQVLPjVE+00uhj0uJlv5a51IGIUJBQf8Zkd20zYKZhERzh19naqhS5MNQJzphaeqxgCz5h8xcCO
Lf9Wlxe2gkIPZxLhkt1Dd7pvvLZs/WwaqU8LfDfG9beO1aDKrOPcZfaJNUd5kw+SRCI7WOGw0HiR
mzUKtfKwJPMTPTDqqGI36+cBDydOI/+GClsbD/cg7fqQRubQIMC66vPvybOs+WfwjdraXMop/RgA
qt9a2ezv9iyWxYec1JBmW+cOv6bnqsT94xoJQ/jz3kMCBTHRpHKPVuz9nFx0RIcPWfy4RxRWuCUj
xoeo9UEMDtN2s4EdHm8iup0OTgdR6/kEnEHwyX5F/E7VElKQkFLE/Msdn0Bw84QiC0AfWL+DsfG8
O0uohuh7yMBieoZkNUJs+4FgBT0KOC9OzgCfrKPBCQ13dtsnPwbyy+3+kAGXXGF337IIieMQUxUt
yErVVYBCY+Cc4WSjUmYMvk4ZJwqq3Q2h0CjFjecpZy1twGcDGfou65ayRVZSyFZkYZH6zdc8m+eW
xXRD/29oZsstfC6nfXPHlslFhANpzD+NgDMFfhJccw2t9ST5mSeSTFRpjOgSKYl9rT980/pB+Lne
Aoeh9qGp4VE9l6cYJlh2uNLa8VRz+UqfJlcOenQ3J2hqShrk9Xna5yM78xbqeAsVU/6liYQVq5K9
eWUeInuN27U2wepBfv6pWzkAqo+fJcqhpCgOmxv3wMyW8GYqPuOtA3g3bqpgIzhGI734PRF1juK2
TlJeB/ynxd6jCVecJCZUj8cbmsdoPTTAmuinFVsNCkdVx96Bl4Y3qKKF7YpUT7EDch8yIvubL3lh
HJ5nCTuycR+/sljSUsmj7K4dlvQNnd5uZ327loMDZeFszcDhNWizwd3FwLNveLBvRbQPwtk4AsY5
FlpdSLCu7EK3WRg2a+iSjLrmH3UvaNPbcPcpd8kS3TANm6O5vJXhXXpN2Fzlz/vILp1r3R3TXKcy
bhcZRvARkYt74MJYm4EXl28lCbUIeGVycZMd0qbsWcwpyFNnQhLdAtAnddmmOq4wyvPxaX2y7U3r
P1Hf/xcJ23elj5XFv38MfSvoOB1Y1U1Z2MfrsCQfjf1S6co4TzsK7+FRedi85sJYP39SP2lqMk5C
FnkalVJ8vLqWrW2Zzra062vlH8I5puVn2/wi+pAAnURv8pvxC7RYr9ligU8qNSs8BpDcTqaSfw2I
orBP8d+84jUxdS0AWgRmNsRX6k5Yl4DMptPCOzYLJUJa2oFvt4MlbwqET+wz1B5mA1iigsAr+UL7
13UpP3UPW+0+2lYmu7drsX7QOczT/S3GizezIbdhQTr22iqlnHFqOUvuoW80O5yH3suEo8E4R5dd
d4rEG3sT//13CDHxmqUrx34l7HvyAeY197xQR9j14EryqnfbOEu0jPB+uorc6iqfbbJ23Vf0d8Ei
PxPjZtCGApQlloW85indRSMmjq38cRfG2vRmyskLMIC2XehY4EggAFMkhHOcnzpM4hWy/pcztnWB
xmfRWowvPFa5mlSfgwGdtPwQsgjWUAaz9ffmST/IAKEreGx5H27uID4Md47dOlVqJBuxI5F0Wd2x
s98pbG2CWbJT1A1wUh4gNCV7iiRx2MeH3VPzv/ii1tUxEmwTALaHDiHmTmh+tWF/ERGgnt4PAW4R
+01KQ1kayvyJuEsqpXWLM5vxQEqubPq/O+If0SGTxIiQoNjHvU7ZgKVTJXBj27WIiXgFNjGvAXaA
Ieb/cRi4qOrYRHgx19C+0AGVBWKL7caQNLKFYTmG7kNZkf20c0ve/GJOvgFKYW8NVnuWVJRlABmm
VP3WaGbk8PVvZW3WxaBy9RpOFMvjfi3s1n1DS6Jhx2wqqybnN10fQYEJDx1kUPePzk4saewQJFqr
YhmZ9tVCTuYzc6lVH+I8ZnjIohSbz7fqaqeXmv99GH6lAVWz3d3KhxQoLHfFFPZUve9P+oGtsdBm
hYgpXdmCN8jxB6WmWBNQ+P0gAcrsiykC0Bn7lMxuEvmnyLUdSyNaaAQ17WH8EUd5j1qqKnoVszPK
50y+lb5iN/90QOimuCjMKiN7Q8j8lII2jivGGqxzimL/vRGZYrjwBzSkUpgAwrvO/KsmDWFTquOC
AqhJzPifATtJI0I3pY5A0R0CMqM3tTDMHAVNF09hZq49rXO+VpPXPfrKHnS9EnFloYRCc8vvCbaJ
viSkdsnezBdyiPZWzSIYPfYIhf/L93I/eGR50wnJCnKsoAZoMbMPparf1zxs1svD+9NxoAqFRM6x
YdFPKhZQ4e3z7LboFgzmGfxeqbb6PBgdd5cLLWnxVFqpjBWF0/wNUSSlwZoSJb3gjvOeNsz7IQJq
dSKyOEL/D30fKMK1tJBGdcN7mMaTfK3MhXZtpJ1l2A6L5WEbdgfWUT90tV2uRTD1hTE8ob3o8hSE
5vYLTY4am1gcWbARsI7YkSh9R/tN3WVwUymmPh1WW1Ufyos3YaeMjXlH06JEIadocq8d70XGm/YP
RS9B1lfsNvAZQyq8VkBt00FRVJWmlt/kRwX/nOP2UQGvJDAzB+uHHF+T4wBi4iH5dqVNewIjlJ+T
H6viSaKbEXG+TAzIjAaJsQmZ7TG/XT2DPUJWSyRZTiQNCFnWaHnaAq/bNj4a6ly66KDjZrNejGkT
oQ+GRjwS7DMprlNmzXF8xRVCHmFVFHxNxPPtxi4fc9TaYScU9vDi2dZFekgV7W2o3sVipB1om/V9
Z5wNsLyG1tHHervL+ewAkUTnwZMUOjJm5aUUiVEtO4UR8JK/moWTUqGx6MFKhkKamZQTrmxCOcYA
Fz45hn6LmP/ZI/Xq9bHz5YJxn8l9xq3LnAO7KrQs3Jwb42G2zDvnar4ZZOqgFdlIwmqjIEmh3G/d
NuHMbp9MFeJlDRXdpC/C0K1KkOAOu6TpDy2F1Im5LbMvB6Zr/5BKpfUGR+KBqX2SkBGeKxKQxTn7
tE+q4cRUBOVUd3AWyULFCvazbmZwSG8yMTlGnQuahkS7echXGejSRvPxNdnz2skkHjaopPsfBnbJ
6zQX42nqMN0bbHrhRHPMFOuKuBRnpCfilFtyUuBTnTvN/fXgHW5bmNc/U/p54zD4+xiurrTl569s
ZAhbssN03C3i8hDWQQv/v3cnZxIjKZgYzW7oziCLOoDbePjvBfWkUMkkeZe+D/iAusYj8linl1hf
5m0axk4WMxIm4DmgjzBjLgk0tUD7/JbAtOwr/Exj4cb7xpZGt+ryP7so8/siAk2znUWqSu0G9pqm
mqcJOVfZtz4GR1XuRl6yVTueE9ZRAzGFG74CCYeQutukE2ZDqZjtdAeUL17IEDB7oCxKfHhwhK02
oI+jk+cfbJNjr/1G2yBgskjoT6MykxOShVDW47kuvUCr76ky7g+ZcVrK9djhE2AEykJxLsZe4Y5H
kk7aEeJfRKc0DImdpTkr3WBsA+oSg4ApnNqJ/M53Lmp5IAxBq6oncRLsMycr2XdhYD5mDCVGdkQ6
hhQ4SrVU97Q4kp7fU0Xep/z39B8EIbE30FETPKSF4aBXsHB0JPbrK3CiXu7GjhmE8UeFjmPoIAeF
HCjI+QUd6YmT3L3k3EA5sW/WKYnzoXfC3etoFGu2BbSfcpOgVISeiGH9h7g4wZUVBY4a+1uLCmaR
m0OgX8+g8ksOtpN8ssFNfd+AoIcilrotvwFKLSdqk3Z51ehm2RoiY1itX5VG8n14tassejBOYzMt
/HmBX2+TuHQzVJbAw2wVveCpkkT4K3Wc4X52QSl9s88qs9fnEjMkdeA6E4VXQlSUy6IBIn09Xf1M
RrZgwvzjHcJcSCzD+jrvzFvIg+g/vfaFYTyrupSPLQKhuDIKy5NVPczXMF/aBky4LwHpOrzxSz6o
6BBbbvOuvZA88gz8d13hIPTwzdxnre4dJON/3+oVYNvK886zjYXvqBzsQkDeN/9H4XbxbWdbE8zJ
8BUbsI1kveAbmQwkl03p276PgbB6qdjlO5RAo/hwO+4z7acyd7fn41b5Q43K3DVSyDbeO0Ude9av
J3iJsksWIEF8vQ9bdx4BXP3PyEiWsjsBKgZA3s0EX/9t2wmBSdaljKR2r479NoApWgI+1zV8apzH
CCvl6hzAkbAECvYWiQffogwtq9gzBy//IZE3lk7k3OmX1S9sLHxm7s4g1r4gj5P/nXiv3C+R+yp5
N7DDQpsgwteHoCPX8PlCiepnbZYOwiJtAySYnyyEyUF9lGXwNiXP0/3uqk5Mk5PETFO/FQXOXPM1
WfuuwAD10eP/oyiSIUKvuoYhSUsnKZO5oyWOJDkOQA/zcIYNjUm4OpBOJfnYNqFyhQYa58TfgpEc
zpowjRnCh4s5M+79D+xXsAufeYb/hwPN4miQBwpVNf55tXT8X/vflvnUOgt/5TQeYxO6uI6F6EZW
58qn+BsG0slximdi8QvOO9nLYMbednGrtbUGaep9p5rz49Pb3oFn2Y25YmJVRf8bLq0+PbXGUzLW
Qx+Eh4QkqzAuDUD4IDHjFiio4y20OhVRUlgBWzLyPk19W+AhOhPegBQOKwBkMJjFydPSSzov8X09
qXYDPg+uvAagTCJoUytqyU+6khqzuVVDK/LjdnbhaphEehGK7E/IYIxsLxNWrEAcAIILyDqyeow5
iCSw6dnSA7Jm4X6rupSLrXP7HCuRX7rKewFMatNm0gdjzpdPCl9KPiiGiewuC+sBK8jraLY+AwGH
UTgIkzkHzGEdf9Zt6ROSOfoQx8xPYZUnIztZ4lF9KZ3clOuKdQvpxvZIK9VY4ASIkh3gIQbh0rfz
SB3VQH4nrlastTyhXhZYhBe8+8ooDb0m/jiYbukAhA0WI8m0JkPakcdgJnEtOitYrFFAQafG1Ovx
ut1zBy3W+RqT8ohvzCVTdOQE34TIf1fLdQygRvpI79Ivqr60ajPh5K2JU2DEtAZU9HP7kt4UNXP+
SkdfJaONaHK4VXiizIDlxWj/pvL8S/V/bqfK42kmxCdo320Qod6gFAjvUm21f8QPm5Dvc6ZdkUrV
UpLj3lqjI6Glyqi8uYuEVZI9D762xSZGZ79C96enY/G5aMcRZBhdU1EH13JhF7OjYrbr/nQ9Zq17
LkZmf9utuqiuCy34SWddx3B4qNoF0NAb54/jMWtcPlvIH23UszVa0k/M4r+D79OHhSuvwlah5Up4
er4l2z/qozM1QXEgtR5+1fhYwSS7akSz9xW5WpyrLurhmnN8ozAY1o+eeenm0tsgUG8k5+fDCxBy
YEuhEsezurpwnrI/Y0mM5cjBkPPQuFx8uJxHZWfFWqLLnFuOqJEBhSd2Ye04eNseXCiXbBn/xQ6+
syR4IfOhHQ10F1OZlYudLayxk95ztZbynOiexMH7OvPvhhMUA9a8bwicqVj+gmQ2Bep8hDBdVYFa
vqo2xA1IupVW8et6YiN3pWHTIZRUAmySI5+9j5hSttFCvTgwChVe6Fm/alkMBhg3zqv3Gkr6jFvP
vt/GavEtEwG2nuXgOFzGbDjOLCJYPuuKzcwIGwij2MVSjzSLUQ7QRSIgnkjEyvVBT3IjwFw92BpD
FGBNESYFOXRfBVaPZgPVzXswgKX3UqyzsnxgB3Eg2Vod1WO6rmdVQADKeS7fK1HGZghFnDIA4BO9
86hIw00qxR1TUsl02aNzQ5XVaiIz4NMqtwQMfoE2Pkx5yCaXT2+mnwgeBhCHiZmSNkJsf6sTZc8v
xqmccVZIQxRtdZxLwA8xsv4iJU5Ss0EEaewFonEuEj6kukPpJJyElb66mkTUiQKdVlc9Tz9mWHfR
McU7v6Y9xs0L+xtOMkJtDEioxcZdLbN72H9fDl3Xey2acVXmF+qoqJ6Fz88GK9UKqozcl3o1WZb4
hXl1nyITrNJL3jbGgt7NP9dcmUrVLC5tVKBzt586BjidGH5SyI3XViiv6sDzrl6gmpKin3nvtov1
2828zX4ue0Y5wvE5lGj4z33u0MSTPGbBKGYiWpBQLFnmA2tHF+5sy+GwL1mPJ5oz6rtbu7tzUPS8
y5gOp8pLaEgDLCnyroYoLGEs06VISFzGX+S0nz1eC66ELFA6ZggHbPsywXzdoiuTkFQML13pMQDb
HP3sW2SzI3IXb3xHjHq0szZt9lhLMxQZWNM8bLv+ZMEpHAzbTtgyrYCoQJH5RnD0TuWsHdNggaHY
fzelBXK/XIpSY83gcRC/t9FAq2GfXXydbLrqgUL2JbeFUoNFqwTrYfF7MCLKoCUbMHRWOOBvAXCi
csAfLuTi8uy8v8axOOvg3JqKj8gbOZPBjf7dc77XVZIT+WVQA9sYXSuMPCtw9FS9UFjEHvco1GWa
bVG9PbAA1xXq5Gb3HzXlZqNaizyPDpPNdQzHkNVVsUclgAkkwYabjFak0YZZUQSNzg+E3j/fSeam
lpih7R7iSt7T9bIHxL2vWi6W5mdXo8EjOoQ2d4bHI6DkM9zaWGCbP/x4ekOtz5d7xDYLKGmemSRz
9vLuY6nRxuHDbLr8WC1efrmw/+Q6UpYLY/w8DOoalQ1xX7iblf6IKN9rNRA9Wxpy9D/BDh9pfX4R
c1g6GbJPGIpiboZ28YcdJCb8xnk2Y8s+XXjsu9El8JUj/VRNuJax0CJIAmWSI+LejgGXqJyjptuZ
lG2h/gY8Cct6SF66CK4bj8AREKEU0Oh2TL9H7rSPHU5keTuNnTo40n3lbBJOzM14y0p+5fTjF2Hx
A5nvemc4vrpA4TW0pjy9AZgA5V86M42gp5jTTYkf7363sSJ2+ka4zL51p6HraY/gbmAmEZcbucNN
owafSLYiRZ8LpFA9hdZJE5k5ZxuL1WZsv5tCT+LDkpmQniffrBvp3ZCfOOnJsk+Rh3iWsKFOmjyv
/huVGuaiQ4WcvCOn+vbLY0lkcS7Dky9fcePC9CF97roUDY2aq+Git14C7+7VrwsEu4VSFIUUoLSI
Gs7uwaVCt5/dETWXC2sgLoChzmqY0ihskJ1IlhLQIv42ViRv7/9jvk2cgJlvHo+w1NpI+iMy/tG9
RzM2NJAupuxBTZyQ7vuGhubRv3XEp8g8/W6i+kTPBZaqJYasbXtUwMEIkNxrR8GWTFfYyf37N9dx
FvvsyqBN7qEuS8Nuczhr1q+mehXRyRxmmKFignlqMiXACNSDIw7gz178LWYnwC3Je6XAIIyLQ2aN
SHpOIkyYh73a/kcAL0MIMztu1+kJUY+uvgvn1dJVG9xrzx7M0GzD65Ii3vkCi3gXDSOv3uE5mufO
50HlqxOam+oq5lEYz17EwdYxmndRUXd9nQDJQqvjj8gKaP0742LhuufzjUakyrJdYbmNWwkpBUR4
gnd82MgB/CaF8P7jOBIaSBugy/lXLd59tOgtAaqCwYTS53jvSaA5icm8ljm4ebqs7C0XqFG+v8Z3
H1pquAtz52cfHOInDRPKdjrddIh8Eee6aYRg5qWdQsBnVh0wo8dqUU2p1GIEArRgHHu9wKlHNbCA
WO8QrpVS03YY+8PeeXYcqQiNJzKfA7RnVGs7rNicXFHJe2JDZyHQgJQbRzQZd7oL4ODpzcvVTY08
0+TqnexaBDKzZ94QQ8sDZm3zTkllapwkUzic8l3NjIGZuWiayz0VT3nPTgRjpU8aFkNK0rs/Uors
gWHBufjOCNYnW/m0/Q6X2M4XfOA2SeBrH/SEm8So8DD9Bkg0vPwiyMe5z1BYJkm6th03xI/eRxNV
F616QLTNNwEPJHRybCM4XJj7VkWUcWUee7C6jn/o59J+SIcFVaVTwqoXeV48/5yBK2pHjsgTGPJ9
fSaEgi1TXJoBFyupdPvGwvwqY6bQzryjEYUAFut9nVd+nuqdnqGGst2EBpygmiUO0AZg0geQPSCN
5+UXbCuSesJzpDllzhmG7HUtQQRFFSPA3ww+fgIt/AioE6fU5fUz305AFnZutIekdTRZMBH1pUjz
V07TncELMnyduK+JJDxXcr4zejzJGKf8pKrMBwoJ6wbgvTDK82YnPvJEG7Px7V7mkC7JQnGkPbIs
4Qg6VHQK9mNb0Gq35ozuBiLWN5B/qOOiQUIVGa038I/Zpqm2eO0MhyoNj3fyoEVsNOpMiUH+RE9H
BSVK8XqCWjNM/CRP0+NPW/IADkTg5T61Um2huOF4AVeW3n95ALsPCJSARamfe36XY9RZ9Lsiitz3
1AfJ1up4RG3BiC+GjBV1OMEWR9LyxE/BgcK21rcOqjHkNxL9D5T52YovLhHmQJgv1tTIcKIFprmL
+Xcyy171Jhc99GEF/QrLG5FSzMEvTUu4NwZTrzdJONtXZIsCMKSbs1UwLk8s5U/O7mgjkEaZLN7u
neYC7clmZBkfYOTO/JwmtCxvAjzEHGH/teErIQ8cqvZCFzZ2Wdwb49wLliYJz0t2/2CVcLAKXfLp
vScy+9JLx5cRrqzyUwSpj10Kj26aOpTRy62Bif0Rzc+GnJL8zgBtD82ZbbQfcQSZGkN+YO6ZMdo4
LaRnCkDrP3X0k/lWVobgS93vYh7wbtxFFLvX0Gcx7E0jnHyO0mvgKzS7YKUWFFfp9Ui3pZUENYRl
4RxQGqx5JiJ76HRkzoTUXjyB8efb0aN1iMvuhKSM32UURu7qjuu1UQDSLszHnSjWZk1JBIhN3Pio
5GC+FCbb25zX2QnBZKBau9ovppVwYSlC5lpaVr3RvX8lsRB0Me4U+Mhpk1ohKAvXLCi1GRUh+Je9
0NVoAEOOM19/seaB8I1mVsljKBkLKDS8wWs3brGEPWsOaR/b8K0BX5yuIQsPZs5Uj4mNI4QmC6qq
2D6WZHcbtHt+qOlyMhwUHwzx6NIKBl/tIyYf8SqURy6rXaTQuOFB+RQS+RmG4kjzRKtp5iEHhFih
nteKYY8FFpfXnyVcMgL3N8j9nZRVbfZag54hVTA0dAwFNU1LPsiwrAd/CSWchxVSCtZJgYh4EvVz
x/rE3ZXcpX8CiVNZx4x14hW7/q7pJ2AO0Hmz+cOpI/IV5qg737fAVMAZgifyMXjNAikTQkBNNV+N
1H+NWL9o0TW+b0xaTA2fRy5hXjuTqxrgR2b4zbhanu4Y//0pmn0/0MmHOrUmLmY6iAypDPfqQWgg
4NqoTSKL/U0KnW+r7h5HteCB4BRxLOI4UkQYKjwzSMqNN5JRhAJ+BQAnCLDjv6saNYNgLoA5auVy
89gbRbXiO/w8hQM58fjNZn0SkivW+2lcZhVkuHB5C5DlnOzRbqcrcnU/9RU+9dczpQsz0UdILfgs
YLqRQEqpWH17TbV4Vtlg2k5kQeeHnZbS38tdiW50AhPR96VcI6qWmbfLQGntbnohENoeefnY04nA
JrkBRu+UPySk6IM0E+ESt+YUSpI/qK02+lWE/bCkNC1xXF5BBt6WsWcDvTzUgqyxK9Q0/9b5pya3
8gRYJdsnXcgwW9hyWOAqKUF8BFS6GEdq0ItWKQI2zQRsvTmsJTwdznwxVU843Q52U0l/DIJFmw/h
0Mx/DFuk9vbOTzW8nsCBXYOZrBkosfgJXjepOVbVUjaJSMw4DZ80YdHW1OpK4t1MuVDscBUmbm1Z
4Yhq0okE1DAatgK2jIGVWCN1lp+HluprbVMwDtOCkJ4SwouxSJa4NK9qKt0D2gaHFbSdXTZUCoEh
lObX44B6Edc8zQExyuL9ytCLINIQ2y9nXYiWCLQAHZ83ieXqcSq6KC2nzKP8H65DyOiIEIKs/P+C
4UV8dI2kQgYfeqn7H7L28RhP2AguzLCptaSjn6/v/A+1/85FOJuI/hESKMwgEDjQ1w+putRErB02
Rfte4ENVUZDQiDEbUp9W7bGlUq089hMwDWEEsiyxLLF9jx5xb8UW/6OqHJHS92mxbtIMt8Do8Dg+
ri7MEqjKQxS9mtdTIqJbYXqE9F1SIHAHkSyd3WMXQzAnByYdgaJr2TMlp0+gNviBRP0sovVnR/Rz
3D/4uKpZ7xAxF5JIl2dgT8gsd1sdz8v/RE1pdRz2xFIb04lPxdQoPSwpbCEwEjcENIt6Pb0PfTCS
kuQ2aY1sjLstz1XJBqrKhOVgEs8J9PPqQDqHzQdJaR2Pi3xtimv487aMj2FtZH/+7mbLR5l/P8GA
BVFEKkOjLefaAYSdKuvcAuZLEiWgPr0y3pZkwUOQwl7T3De+4YC0ugGz0IVpd0dQTk2aDxxEMv70
NZ1EAi7gw8+u20f4v2OpA5EEP/Mr3LnLzR0fEprjM0bftqT1PIYpLF5aKYCjbZthf98Qy7OX61w2
ODT4WHZR+PjWlu44RuEiEBypwkz2Z/HGrAoqTiu9WwCY/MgG/bf4EIpOAKBMmoV55Il3ZccZ4Dqe
ggpaTqpmE4QwbJdoNtcj04+OFyab5mvz1HqBkG51jouyPuObK9K8AyZFGCCBC3jZIRqt0a2fxHnJ
VbXX/889IsyOHzZPzaBN94Kz36x2G1MLAgy13v9TDfYBoAUpny1pvOxWHwJlT3DQRbO3rZUw2JEi
ekEdov8D9nmTGPu0fnNAlWvfs03xFENnz/smw2kKp4Et1etsA4x6rl8yq+MVYRf8CHDDogpNHf/d
dQVSe8OVxi0gAFGlWU++fRtd9V6PYSC+HMy6c8lRcEJ4QaG/jgRIaNuJW+z9fds9Kqre4VG/Rtc3
wnueT4k3Fc5oVYbLxXKxBUCejEyu7oq/DaXvHN1fGN2ONJSgSdJQJsNZw3CC/aHmUP/CeGrBU+lU
1yxNzcaW9pFklz6LyFisrA3p1I0UXyhsfDDdnkKOV1HJCYLKcrtHDezwPcapL8qlX4xV5TLNETob
TqzZA8+oxeXohDBf8kBiB4gH9d99J88463XuEWguYkUDHUIR1KrQnCozFnQoIjDv3e77KMFJD/nk
zZqqbAN++sSDIlg1RJc95Puljq2mx349VIlrs1sDjvqRzSGmlDsLTS7jRYm2J5W9Tp11a8dP/qRU
wKonbl5yEsnfIZ5XMVgis5tFffogiWkvFmKcJsgIVBsNJnhk/6wocWovy1SGleSpQXsKOhxaiecJ
+jbBwETK49TmqLs+QD38oIQ2d2EV/UVWmxgkR7zXwDa2NNsx7xpvw34Kcvj77rCJjn9cSorGjQQl
6IACuyoLLPLPMi+wD8dWmWlw9yuIv0C59Ql+b7o2WJKWlDQi7n+UfxPISuNS/nt4UsIbX1c6swv3
gzOMbhOgi1ny0PthOlm6c1IjsId68yy+yTk4gZC/s180LsGsEP/DYVU1atfQL7gVzM6d5EasCDwZ
ojvCrtWcrhaVRsHQ3bJ8NvW7KxXUaqlhTvSuA6wEEfgxc/wgfq6DC6MTXUfR3zIeXinnbdKaB4cP
5DITl5Y9FnO6Sk3/VPt/yyoEXikqBRhjBNwt84HGq5zd4DtJaQsSRUaHpy+EE2hbHhQgRK00Nkv9
IpBzj6hKKaldEqvqZzNGTQ1VrCaBb+1h/xBb4GPXVVKmWv2U2mwoQ47LpOwVF2Hiw21wGKvL8Cya
TgRDAM04ZytFpuNw9ulVgxmjnXfyjkNRdxWNVVw3ggSDyitEpEJr/OviS4rzlB7u7wuzni2cA/0K
Bl9rcq1RaTDncjLHegrlj+DM/4y6NR1Irm55+Zn7/gFCUz8e6IpcZtGUne/MGsXfgUztvhP75cnU
xRx79s0IpwoAEYqxSLGpcd49utwVPULHute62ZFlTO3QOLwsGUmBgRBNBKDAldxWqGuYzNLlXO86
xZ0SWq6gejSWeTA0+EH7oBCqOtz+NS816odNNRWnjEu6JpofyrYNyS/vUs7n4G9jSTjVigpK3Smy
y+I698MSDmiEJVdA4CD0jsksFQs1rotM+LIniAjGrODpr1TwFK3BgcE3ryBzRxClfpNOFijKn33v
kTXF7KTYmPqVZN0GxEd2MaGvySBaZbesGcWIY5OZZGMPuzUAsHutV0ex1r4kZJfHwLpdfwh9pUr4
+HqS+84oN8IxS13ZGmaWJOKMNqIkdCYgWmuyW0oxZwmk1OFELtmfifVADD3SZsFOHPTXPVkGlovB
bdhxB+DHrqk3ZrNflU8n2Ds1rBufGJx+/MB7st+k5MvGEUhOm0hqXsJAcwGPmp9HGI5gz2i1CRTD
jEbeHeYxdb9BiHUJUsdscwRqoWz8vKPJ39xGt/0N3Mv8d55y+R6B7JYdbJU2DCbjkSQpc7+AApJc
GQmI54k4hVuYnIAQJmydAM2H0SssYTBgBjJdFdvmelkre8/e1kYKwa3Yi8tSdDBu2XwZgzV9gkxM
TMxr+2AcltBB5mP1PLXnzZZuyLMJDUhq02Hqw/xMDond3YhQaOL1qrQ7emANZb/JYfIo6STpDj3O
RxKO71OQNGC+B9SZ4XPXAN/889wPLvLpC1GfNdgBLvfQmQl+Dm5ufEYxLd4MZXP4JBrnru46fI1+
JGYeYxEOqcGkRFzY1S6iFe01Hf5+QyykV678EiFw0O0q5qdZSgskdCnMUSazuxZyz8pfunlC12eX
ev57jI2Q7W8slSSatnBRQi919iCBz7OlDLxfLPjKP9X71t3FkL4LU+TPlW4ck23PRYA9+gsi/vI8
T8Gs160GXmixxIKmKMgNbwg1LepSgcnuy/ejzB7XrsRzIqDOJV2e33NEAkohSJrlCCiR9lw2OeLW
kJNXl62szFNS2/Aqbpe5VxzXCx/pPRlluhuScBHSugg9S+Grti6LQF1sdx5iHog+FSZziS6zm7Ck
1bciD7tyJlmbiHUTUDHv7toF/jyLyx8EvtadGWBNJngWk216FF8OLPDOFfvvK/tf9zRvp/I6dR2E
7v/+MjBh14CPzoEAScB4T/V5DdfPvsFWf9x3HDMfOcN/sWDHJdAhXjuIuyJgRB2U7uuTpq3FwPhN
wqS5xcFTElqia2+amXNPO8X7ZE8USBB2tOeNCLqIbJmAbsELs5gv3xi2dtt8muP23dY0FpagJ8CZ
8cCDsWKvTLmUFy0zvABCuE20U5V9fj1tr9vcZET2d+UDrrk3zV9w9jcLtgQHT/+gQ1xtH4KIaw6W
sm5C6JHIGnklrsiCaK3Gto/dlxfcy8mIEBM+PE9pQVOsMh0HWIi2yU8CGlV08IlIt1N8WICXF8aG
+FtbPbqad1QWsD/6MAk17sv16UcJUJMdKopW0/4mCBQp6RoDjZxLbwVQSCRbSh6UFK8uzJ2j/K/n
15Yasc6U/rF8vh6tKkccLgDt/dbEAT7ySywPWmxe7WHBJ3Jb2ChqgC1qvHpB9dHoYdkm31KCZ3ae
KxoG95Ab/TDVvbxN4bzVn7R+1OIlhle7oc7dsg1RJtkP63kypYdMaKQ//fBjha6NfzfHVnTjH9fc
h/XrDOnxSblszFQO64I5YwSChiJfG7F+8qFHBiK18BOKOwf0D0qGbyp2l9q+T8GVTLQmt+Qw36sk
fzBizJZEAOlwgydZsjpe2MeRodgbakpcWiRe5A9UPFq7hNoUFvd6CxKquxTdGOqtmJ0swcObmi3B
M961h5bcB4SybT0eitYGGqtzOlSBbJ9+eClJby4IHfMcnFVHhKxNjY/FcOwJhiipj7LJ38W8iU2s
rqniFy5MdATE5kZkQrEnlOUtlJg5NNIbv11wV++/wfcPP5ABw6X5HZ1efoaho3WS4nJF2ur8J09h
gGrmVeGhyr9KUGULMCrQiagF9EbTVXbIwIx/viUmODvPlwILWsoeX7Rt67qXQwIAm5BvHg79uNGs
q1Sf/4L9k8PSitjLATR6aKTMZmIJe6o+Ni/+33YpGPL7UL3jhdY5qaasFQQZQP9/aF6lmUYY5xgp
skEw6RqxModcTqtUgwY6yzLa0bp26l7oi0BpGgw+EpFmymasvnzeZzClqNv+LaEe2mcHReeamQYu
Orcft0WfgWSO4/B6AT9kq1TJxDpLYeXtj3v1WuwzXjH+EhLy+kXvr6OeMMcZYGEHkM3eKkBKXXgT
tsYbNieZSvbR31KZctSBgD+KZXBWx8xvTmCfQ0d4y+7EuX+icqitavkxF9S7Eh3CMrlwcxjdUN1h
miOTIDKJ7pARnOuqeLIqtda/U/2juCCp6A46jKvffzHCGQpIvR0jDMsbSSbY7UyodDH+kvu8otrr
S+4+Zeo+9J79cn/uHFumc6dtuelOnx8z58Zjvv0n8wjhEr4GtX5Fj97Oju12iCOdOqRhR9kzd4cL
Miy+yLr3R3Ka+dFqeeOAaW6tx3ABD1RcLn9wgIXUct4xD/RKY1etiQ11KH/8dC1g/NRGi/iZ4TM5
NulnwSgDuSJqG3q0AimfujJdWO8mysaAXt7KH4fbyPEHWKFGOjC6Q6oFs55NUXcHaqEJJVKCNQS+
fbv+bUvxG0KX0mbOiewXiz1QLcuhGlOzLqgIsBiH/50DYCaLNilFEzFcpNBpoM/UScUpW0MtiHRd
TcdvmaNTbmgqgwDwO2siewMGIgMkS1ApVETocr0d8dae39Ts2KqtLQkSaM2fQj98AQE+W1tUmKDu
vNZNzu+uIm8DBeghxQb2mtyGrLH9OvdLFg4j9DIn3adauTRz1LQWKihKzw/WzpQc5pr3DvTxnnw7
Wke3OdXx/a/++Mi0LfB5fTign6ptG9xKae2ijygladq4BHbZShJ+2kDnzObfvb6iB6zOhXsoswsi
NF2ytOT2bdlLCktWMiYBbdDi2FnnILfsQVBFr81nMhhBJ1BCIc/qdtQo7xgfZM6sJbdUdY30TD5k
gnmvpyJI0dnmvoagEpbmJApWk/t8fNhHXeOeOsbDYe+XaidaI6GQ8XCSF1z9dUEjMfRfQyyKeCPE
vpyAuPnMwX4T2Ijt6gygTF0QrG8OsHb3uydBq8EnWDESPzITgC5ZM7uNPIBs8ruk2IV2EGUw5ZHD
g5Ddr7sUDyAf0vKPmC2N8JGd0WF4ZspcjLRvJ1nQK3TGGRQlmwFG79P3+aTJjWsKt3RlsbTb2fvR
3EsuBQCHeeEmLTN4Il9uluGtnhb++8mYSx5n2tEnMsyTHHKwuBRk9+Y9US0G2PcGJdcQeQ/qRdC8
IT44zxwg7fMIZAGqO7ze1bt5qQLu0nxYBQbE/OjNAqck0OLslOr/JxbYVH4LmnTq8UDTWs4plORo
yXXeidOqm38i6s+idCw7b3s8E9L8nWZDAHjtFXE5QwJM5JfM5fMbgCc6Fa2k+y1MnQi3KdNLb0X7
a0JuiamhW+ByB5kIaPTs3T3uE0gt2yCCUUxK8cEswj4fA4B39+7+mGOSRUKHHOOsdgkO5B02rUQz
D8tM/3FFlvaHvDeLGjLOgjXyt2DnBMtStHV5E7U/sC9dD3i8PTcL3XR1ytlrorggOTwnTWvPIVz9
zHTtaQQ7myDjxz0vW2ixy4Hx8zxKdZfqzoH6qCbqFKqWDDebDBBfWfeZEjboxiLvaAjJUvHZyi4p
ts9cLfY59Mqzzj+1vdkulg+Nn0ZKxtQcWDa8O0N+H6nqon3LtPWYwgVX7Fn2Ac0WIUNeZqsqKwjE
EAntygReDwMKdng33yM1ViIFn9cYAdoE4BWcvebQewp7EoowOCTdJMPAbOlCKbZLjiLb8LUo29o5
IKxSGmlrhKjo3UyZ9LZC80Q+XCafdJ/mBB1ukP1R8NyUNqTpKPm1PDiY/G7/4B4nfWc8Y8ca4IOL
fj5ghjULl6D2WgpODtPbAxGHftj4wEngZGDJutcKf0xWYxI1iR3PGx1hj85G5CJZc/evBYQ8BiyV
p9YiQKzRooA84pIcR/q+nPfVphPd3fXWYVYDcyw1Z1MDBKOgzLBtBKFGaqoQH1JY66vnGyIdrWQD
iV2LvIUESoV96zF3jDVUJP3vLA4q1JsZYaunejz2UwXIWVFbksmyDIpivHTaM6oaxAevebP/eYvV
Rb4j5uIDxevoK4tzyrjtbsYoNY7B7Ih+hOdcZ2AM+XRsHwc5KwpO64SIy7ki04qezyScrdFJ8SSF
jLratJNIAW0QsqMkqR4lpKDlZlfgZ/JTRrTBE1vdgo0ESNsTJ/wnCUo6ulxTs6BBqkZgWmj0oF7g
hkDAOt6JK9DwbPcnggvXaRRtbih29w5W3NsMj1gsHU+JCEuI+OIDz+79gsUR4wJ/isCwxoTRgSLg
FW3Q3Lzn8EhsjXoPEUvk5tdHnEUvPbCxuSjjOIxsljtdItOtpn54HZNeRrzaVUMqd5KEhaz0UhQi
GS+VBqd1TK0m8AEKEDCLn1ziyR1VMElSOrlhk0+UC3pG3ic0P/+MW4Iyi6+lnf6+JcGIFDmcMhhY
uPHcwBCLiA3nZPUjCdY/097Z1eh6r2nfFpzU47LYpyAtKRz0yD60ikj6KGbuSHfpOdgDLGsSbDMb
ZqAqLxhyj0twcDYKLomuJcVs+yxQAXj7q0ZaSsTQ6iujEgSA7I9luY5EOd23o3VVdae18KUKd9pQ
7CfnPKWbg5Y+f6Faw4wNgBBLFcM3SA7/L/v+3wEoQhH1INLYjoorKko+dDqTYlLTiz0cqAXdykZO
m9wZybJkbxDuLuiB3kPDUoOj1Okg5VUdFKfTdEzalxOFy3VQ9URd5a49SEnXRUoGb1QCVnWOQFgW
ckTcRqG3tr2V4W72jhheiTX0HySMtJZ//dfb7hKbL5jy+HAvQDbyURpeLGGv/s1+OfwGw8qP4VpP
eXBdanCd2GUYweqEPqvSuyqRT250nsqQMFlPUzIyMIOGH9A/ZuRo2chTmAGOuBNwyEp/t4YCBXjK
k5C9OtArJeTYo+duy4fJjEqqDBvwiZvX8ZrQpkaB53HbT7Fz9kvexyOhydIZuqSdLcwSQZ/uWQTl
2A87HsemILSCowQsQSMd1rfJZ/tSd7YlsSJJ7RxjOGeRistT7NFWbOCozTlAom3bhlowSbc2K8Qq
VWGS1UlaODIJ4o0RE9ZdTSbFnESvGjU960aiHcpGvjbc0OCgE/kCfQVRRo+ypmczCQENkcFQ+8Xv
SXzlWVthcuFhCcbIk7OkqzVgo0slctApdcS9roNX581N8PKEc+M1JgkL5VYj1PwDmw74Dwji5Roc
eor62SL+pkIi9LAS66ojbaLg0JQxc0E5GsMfXjNxAkfkuaDv3wytrfFZiJkBu3d2RW19Fh3qRnIg
8I5cvfH+nVwaCShJJwc0WEyjjOaF9JXk7zHbOT06gPPZdiBfz2ZMcp+mWyBbMtltfxR1kbF8oLFo
yBNGLF3Egqsv8sRFCLm75ErnN5Abcz0DtbeWPJQo+pMzd7nY1dUrSJNwlFf1JLT+Fe6939EU8SV6
pvYejmzC+Fh80iga/tMFe7M8OLy38Z+JcWiHYKIhS1zZLZCr9bs3PGnObPx6Y9IM/Lwo9b+xvOVk
tMw1cOyhn1kszX9mk1SPbsoWFHOYMt+HB5HqcRseKci7hSxKshVEErZxdHSfyxOyqH6XFVDbTHA8
ccUdXIF+17tuzZadSzlBsb8Qw395LgQidiij7P5TxETfGQ3fS6V0K6jarqQmPNPdTLplRoRnl11S
f9EyZhFITqEPOiok+f/WjXrgODJwgcgtzsD7vj24MOeiaN2NoMltaMOA8ufZwc1RmK+KPZEZhpdw
A2SE8Wv3DO6jX/lnVKsyYPLayAxs+QpswNF0/AfFC6RxFWarYumEHc8OIc9zLL/gCwMVcCv/GrNS
DOkjNsxrBjDSINt8yRqM8GRLHES70TsjraKxSpBtIXycJOCgqX8S1mHtDzFaoud0+MUianBIxsCb
xZpNbcMd3dhjYBZcmjBHFv8nLgci74YX4WZWPk1Uf03MeMewF16XMsrTGsoMd/VeA7XGnC0piW/b
RZlqaR8/aYR1JK7bXpeWO5iLes+mo7q1KBEYXjhsOIDP4XWzh8o35jwOBbBzMxmT3f6l4LfMXMBo
+2coKNictpmvq7Vdyhr6WbnOPClZFX/PKEwjmv5Y+Imzb87DdRL5q7jq6Dp+vwyNzd/9c4QJcAzd
25i33C3WybcrZQPx2+786XQyE2Bq5b5KLiggL3Mou46iqs9OALXXdiEGcqu1DeY3znlbm5X/yoZF
lRb3jmxTdgrqAq8uu8bdOd0gU+opXrGlW0ecw/vKWOYcXS7b6YNdWNhsBXzocXB5hk5AKMtMOrIu
FT5P7a32MYGTVGiBszZZt2c2JQcqcLWfwGf9syuwmJx6393shmEgp3YX0aAjBDB2Ac0cmjsN2nYh
lFncA3ONtHQAlS2R/nN8Be0pv24kKoYuX1MIN5/ZLdmj4ilROSPtnJyaf+5pd2Ak4WmCSfJZsLky
zoNTU97Tja33uPjKa12OpStvJ+DAYGmW4uZSYCQ+JXSQ1fUzGrnpJHyN7fTnX+jmQRjkwEuip5fW
b2bz1JiluvRMNTXI8bC9O8Eca5DoET1su+GWfSW8pGPJB3rOe+yjYW2egczgjkwbpJZ/UEK+W7go
qUSoAT+d94mwo6I21Bcri/XrOeVxvRc58HhjnFogcDeLjZUekKb3X1ETt0PmPe9yi9Pb0zPedpmR
LQgmvVTzCVQWQ6r+73HToQ3XGQxGziqOpHke3mHVPr43sRaQK1tJf0rryssb5X7kMciEZ6hVhPjG
Yqwk+wsiealJXUvX4F0Ew/IesZ8Xee43rl+adWHer6DSS4EtrTNSHfBzhU5iKcLYml3pW6k/sZKa
VOufmv5RVXe5pSCSRoczgvafocm4q6j2KcOT6A/GSC/LIb49tXWTyRh+fxJtRooL64hnA3QXAULh
G9Aj2MIX4jwxMOCyrtzp0tiNwi8nxLekGFLO6W5BaKxOZqYBt4LruXl03sKjjZGSmO6Xboi0+zjh
93CAi8A609Vv5PXxr6CwUE1nzWB7/ms8IIdkaz5sN/siJbdv9E7TlRpQ/dz0HM3tXlK65T6xZcw6
Ii6ksiylPOHriSk9w2je8S79JJqzNAnPjUIVpCIWS9ka3V2vDUuMujRw4lZkSyhfcwWoF1e4QuMi
VlOwnA6iidXcDi+4Ma2DRyQozYQUmGed3r2akF5F3cdGkCvkO3hT6Bp2s9WXmhfZL6bbNIWKXx38
n32e0CQr2RPae1S9eww3EmLRuhRs8cbnLx4RDteJzB9ksN1CBcJKeWia3E5iMRFXpftvikuCWVvU
hDKk1ebg4lzqfi+plzKWIXh52Ds7kSsaQnPqIrqt9Xa2J3F3t72isdjxZXNKRcz5dFAPdpUN5Rkx
GdDdBVHQxQPibBXVJKSM86x5AkW58+VNvqPvyZNBRFtlnoSY2A4NF+4FBfh1CXIElOBjsdnl/o9B
EVb/5Ei+58J/4OTrSU0VBopaxVT9JEn8wD361XEEFGXxU765d0Kj1dxwueJOFUphDy+pUJTI96js
eekP521WUbrPpBNc5vyVExpHerGW0cebh38khfVKr4ijD6S6LS7a/nsypkqwSCJni99amVvtck19
suTuGqhSW0AvZByQdxNt9wNOQ2Ft/jpcI8Z6EbUxEyPtrvceASKl1nQBgPHyOrexAZQy3r3i0l7R
R5AQVoxofiKU1ghH7eKXgFnbnhADjFD3xQu3pYZCBdsnKNK6fbpE1maW2v6ts2Itygb9pAYstyoG
DJYQpeDd8hOs1W1Dist9dIiFw3L8yoQnBRaql4OUWEIfCBK8FYSPpBRi6YVqZLwlXnAzLvjU1BXc
KOzGy0wxNIS32ZwRovq0Uv19z3g3DgbEUf8kSoFiIDd2zhbd+QyK1CWyr0MUFyel1dD0TKi4oPz8
iXlAsdpadKuc+LwDubcVd1xw7sJ1A5WkGpISrxvmsxXQfTaLdB4eXvCjw1B0gEHPHV19IMjFagmk
JLLQh9T3iP0E6uo9xPnsXo2K549xiZU0inmCe7FQ5xlhyA51RxJlCY+Rg/NIsGzpU1l1tlFjlHGC
5D7rPapZxhslQqMItjA6s5BZ4bcjWZ7pYRVzRtGJ+ycTQt58v/WNVnkt0ylXNNXOMdJ8JKZMQZ/G
ADR2sgfHoSYLclHU0zF3bJP8dzPQG2uITo2yiz0zs5JsT2fodT3b0Ulr5WZ3R6rVOw2S8bj45ajy
znfSpJ07rnpgRUetbHFq00o3ZUCev3oEfJJRmmON9iGHDQb8bH7qtMus5bFmAFjkdJOcWbcoPWWn
uqIkJ8n7z9tDMUSpBsMKK3huFix9YahfsIWHUHKGvHacVR4mXTLBYYn7dWuqKg/noL8cJ2e1L7ly
aSdTZ59qgQ1mI4A9IuziTwrjprzvnsx/nyA5qY9xMkE5q/RSKYuJCM4XpLnYnv8uPtVO4ioDJh8Q
FJHqAQ20Nx+8+2Gxzf/3S6dfyhWghv5yldwvp4F42+Hdi3rCj7pz8rC14hEM6Bu9IJIHFhdMFGT4
TVSYErs08YVo5qVLaMlI0Vri6ezKhzf99U4VGdyFk7Jj2Bp+cQLBf90Dvi9y+1jU80nIVBVsmAeI
Rl85IW4xt5JMAwVuqqFgEVWfHDckNHrN8/VuPqaV3X1OOBGp3AjCIRD9etcq8iu4lu6DGjlge4ry
Plij6BueM/w7GmBC6YNH4bGSU0uudNnZYJ6teZWTsrzxQyIH7lP+BidEAMntElZyOeBi86Ddubco
+lFFC5KrOH/Kb8aBioEpadfBqgVCaXg5a5MTPawlNhRDJJQt65Y76UfUBqPlh7aoyU/7Y7HzsRBN
ZzbGHzm6NXX53jqj8IGRDhl3WGI/AqS2GABRlTGy7ynQcsR+9o5M/Or/Jyhd78sI4wqd80ZePQZG
ea3/eK0wX0hO0/wWtAps+/M9YpSNgQzGaQUGZwQX7Egv1JEGH8lWie9jN7OQqdKUfbSDP4Wa+YtH
iVAaKr6CGxhDCbj9hGX9lXzA+l3majyx1TP59Ltpxskr1Ey+Z5UuaW4TS9GQP04/KugtEanAuWkR
jy/tV863zAoIEC7jAvD3hG+CDtJdiRKIpEcSACFtzHkiUXScSZFTvs7Y17cYat/Cp7+uBTCVySCT
TUPLInu/ruync8gwoSj1AtfPUPNr8vkEQeItRhrW13oykcrgCEMjxxF7F+xKaJjTZb3KQdC8NAUz
FFLjeByWy14uW5b71mEdADjmuwSYmPJriMZTpirKXMnh1EE4DX5XIUq8Lael75DiRG/yO0MczLXZ
ioyuXablM9is9+0vTASj3kG0f1C9TUhT5SXgTx1dTLGZPimI3Y8bfINd3FEDrPHsgFlElSpzqpWD
NTOn3MhJkZMYMsECG6+ZuIj8AOonWQh7bx1Tt+Os5NlxYOj/MmOCyj3mLVkQ++9yTzdsoKsaKPGR
2X+YgbYBPeiiaddsIPhwj+r8DbeJ2kQ2J7V9If3IyHEW9Pe+F6UC7uCN921HlJylxr7zQ5mJU9NE
tdE/QGtJesJ1hwxkiG/vSGccqzQAVmFBZq5AWxJG4pi6mGWuHfdbc8sn0G3LVONdkkyFQw4ktTsm
W9KPuzIlHH0xZewPDJS7ScSD7re/c73YzCfodvnxWsFoWczgcz7JDzQ6TAaL0B4O0AuZlVR89oMB
I3NjPPW/tPgTbHGg0DSak2GTWWdu56DLD4KeR/Pjm/42mjTAUS+WbSZnknMR2ylX34VFkFNSMYpf
Pl90hyjd8uS8zMfLlBA4N0Sbp3NC8GlxbNLzhWcz7iNFi2L9l4sv80m7hcReztANe50Er+Id7mbS
DNJuaim+nsZ/2yK69ato3QAT1IclWw4Pht15TqwWcX4YpYoEvBBU+4YAytGwHcKtEmgXjpmwA55x
Gg5nnlOHEe7b7fdCLl5Nn8jEnV5nTbJMIlaBhNOV1/7URx+5C3KPkLUdrGv1axJwrCzNcUqZwfPW
1SYmDue0zqbLYUxb/OvTN6aIcbzzHk87lsWGM+Q8Rq2ow7lQAJL4dnsJfrdqZ0mbqk1sFYwLpXKa
5X2rv/wp8KzCGc+HQNI11aWcFwJQ2lBLmOKEilMxmCXK2cAkcZuXi2fcG6dde6iNGogJpeyrjf4g
ZmJ4To4sCVCXyB/6ngrlpH47JOln3Vz450AcWH9HwggxcVn5R0QXFqhMRZu5S0GRWrwEY36dzui9
RaP1p5h5VjlWkOv53yE0AzEXs5cmARYdi5/FnEyjDzbMxY9yIBkc5BKrc3up+KGYU7CeN4TB92k5
ZNQQZGOE7iw0Of12Q+A6b7d58lPD9JYwsaoOE05DC8OaVE1viyT1VixPsVn4g6WoG0fuNwsi70je
fl+NNb0I+9w1HDaFhFf+0hd61LC/PtsVS88065RRSeJAG9fgf3/AeKI1kwtXYILaST+M+IQ1reeh
z2tiacfgtAG8GW1pMWAYMKBxGAeb3sw9S4s+nkMPu23TXtxdleLQM93t5/66x8FVUj+sskSqGuXi
egtBvvIvqaWEPBaCT7erzkBqB6qb4E/zb9pvQPP7DoCtKxqyUxPud202EQTqL0fExPuTKIva4OpX
x+RzYEwiJ5NdX+UIgshTnGNJtYjcZUupM8lc4xupoJEDpd35qY8qJ3y2E0He3RdPKyzw3X8GtM82
U34fKPIIF8WTVME7udstsPqHRfSTpR+PLAleZBFXFXjn4zfrmevi33yw5A0MTDybIQ8Z8uqD6Zpd
4u9YAhoJmCleqAfVt2Wb4ITP79e13ygYvUWn65kMRdyPwN82QokXLcutzd3nhhHDliLV9vSUL+lp
MbWQFOPKZ+zlxVDQFUyAkBiqXjAxAo3fhywDEw7QYoTkQYVdaQCqb3X6qVoQdQGuuF0TB73/pm2A
mbtfMFvA1sUS1CACvHKnMJhbHaik2+yUysh2ZTgFmWphGZVEveZ3N9KU/3FDGEZ4QrmR8AHT7iIY
IFF5Gv2e7vwq8vTBFT50BWsTzNB2AH1YeJEQy1HTeSntku+8WwEY9MGmHEMTwKAMd4OBVLPGwx7z
sbI51nnrXtL9ORwGeEg6WOUdU9zFtIT5CN5vKJHqva//UQY/JjLBrXQfVefi9+EOoSfaHbmGeTIg
ebw9WN7PTUxR15p+g01pGel3jAL/woAJb3LXPcqCHBKG8kaSTmS5YxqZfKV+OGZmNPeJ0yOazZbp
MoGjVyK/BFf2AEW0COKN3QPr/i3E3y+t7+9cvroPgXEFbyWJlPDrYSBojjeujQiDfkgzi6Ivug2B
Ocw9i3BaM/q5pvENJHprsWtSboFG5C9mMR6laWwp91UPbwuNZAOhQdIHiS5OT7Xa435tiBLvIp6O
z5R0IyCpL8RUwzGkkol8Np10Cdpeo1xOZssYxeVQDU6wttTR1IfuouNowzV4qgfCG9ay2iY2SYCR
gB0zU5N+4Y5wDlJ3/XbWh78cZQwjySC9uS4ZDAFQLEV7AJoJmoiuEE77qDBzlxQ6wmVKWuGO+1KG
RIZ7FsHViMilU16mSYEEFF7FI66GdepDoMpJdXHPaUynyDhdslPsDCTXw6yOoWRe8TUiP+wl6LUU
gE9yx+ekutTabhc8yMsXfLMZwt8CHAUbty/SCvTFIgh8IYIPg2CvNKRvrUbooxRjRDkLEDDAokN2
XDLNT8ZukO6IVamsH97qQEU2DaHj0ByrbXnvqpWyVosoWOsWMOHEatLSH3dhdFsBc7kCv6Ke++tX
2o1T5m019B3q/iODuhEycg45C4FxR0TZG1yoBNND6aszBLOhFu7x4HpD1KTxOiGbwvrMj/8rUGgU
vyT1N8uXWJKvzVFb9vGEl5dNsvjgE7tnj9xNMeRM9bnbwlLNHd+y3k77Z55CXxqNEPRQ/1cRNp8S
ZPrbhuiL/Cg52XUS3ha3FBKNCKwqLl3LGxcrk2OT4gjH3U602bjVjquEhntK5FU8E98KdWIaIZpg
6il29SkOODXuuLlQjzlQBwO+YKTBLGhSYA1/+XQi1OimqLkZ71l1sPXYU6uDbBJpdDrBsGoj2Az3
9z3ymfMZ9fMYK0iBlUV8/339POvany772AFo8LoPHW0657XhrGr1UrQ5GI7jWgjQQiBvL5DrWMNO
Nb22w5Z20y1XgV7035kzM/Jt9eMbU+ZDLF8fw/LJaSI3KYjYXYnXVPNPCQDxD4bGOBvxhv8RhwsH
eyceqF/R6llROjw9f6RrciDoGxc+UyL59Ns/EhIkq41exRcIx+zlBORiatw80ofwtYl3c63Jny6t
C8bctL6tCL0rUKQvh6X5oyVIYPYV/WvKbbsnpIQusZcU5fw7Toxl9c4DQVZZmpHNrOo23w1aDRKU
U9LpKreomWtUQdvpQANnL6FQJZhI3eCJcZKCdJ8fifSgpuo5kPOGYaTH6zhukyrs3Qu9lnWZkK1x
QZrxYKUAGZOtfwJYv73UOihPz+RwXPkY4mWm/8pD+Md57wCCPIJY30+pjROKCq/xaphXNCv5HGNJ
gs1XqegUxUPWzNDxuaCRMYagrglG8TBRyY3KhF4qs+bkLO51f4+TbFRVxFxiiYXxnmwDb5tdJSnc
UBbGtffwwRFVFkDW1rFsprMOs0tplNIfJSGthQBjbqha0vSQxNElM7npvhEHq3rKdCjgbw8MLwAQ
kZmSaVwZEvwgs/CjKUUSydkzSHgEGBT5mwCpHpeKIWC9ev+qn63Dp1K0tUntKST9N3VCtm5RHBx+
UHeeoL3AO+pEAjWqeJkiUd5usf9SrjXDZbKpWBH1ilHWWxsbVVih8C5/Hx1Pv9wJynvIPVE49Hp9
oknmI4syx0oIsMCnQtRJ/qxPZ61GAdti2wK3QDircRN0mChIdhDRgHFlgJPSkMuHbTVsCLvOY6ha
k/zwmBkm7wW02KN1hPWOGhofkvLYWFAu5EG3aqv2v8vD7NOP7ak7sbdvJKEONg/3d7Xfsj6qxCZy
oAdGey2grHni/RNnoqbBxKTT24Otr3Bpaz2q5UOuJp1uYxz/Uaxuhr7Qrlf8xzOMXDSQnm20ttbm
d5t//hDuzUQZVpe4QFTUw7wFPwXtwASXMM4cw/sdafd4A1RPrgPn3TGC9Mxdprif5HLRn9fXsoLe
Eu8VtqQZBB4dk4XEb8j8qTVi8IUeL5Oz7/EeOb5U4rq1b7P2p5YWBChwNoNm71KdMS3UgiZ/WuSy
/7DuFMc+NUs4KZfvfPJpPSC4k6WOat6TNNL/CKyJybVLIcWGtTP66LwaaYF2CRM4z3nCCF3JrH3R
l0q4T/lJ64BhpJVemxmOHPzfNH75ShRppIomd3Y+/GaFVQowmDg7S38TNLpu2HWtzrWnbDahzToT
7pjOM1dxNe/Q4iLvUd2oum33IVLR/t/5xIAERX74bpwT+R/vxpm1vYXqudGNqFyCUHL59inlI0zC
jPKZDdv04r+gRSRFKtkHrYM9NmJD1CvsFQFu3lG0hx5SDpZu9o50WZHTj+Lkykn93uI1EGXyxTDO
h22gNPKWReyG+47/2tsH2K+DkAYhoJBrJqvzN+9tsQtIaciXcRapTq+7hj3DJ56StxQfqS690pL+
yyozA1O6j/G7V4sP7fyvsQLyEKbi4UJAviReJZMK6pUFBCUigXHvlhArilAHelWhCBpcjhuplTG6
nnjCUMM3ZfT8jjaRCm8uSr18czpPBbymHWZGg6yuKzCNgHzsT3VOkmDBv195jdgzgvPAni2ddfm8
rbfQmljxLnjdveTWKDkUeZUQWvs4kL6AGLGj5iim1Lc/0xyoAv++vJ1zNtGAs8tWrONIo1StnbkC
q1qNZh5HgIDDvoSOQgMP1MvYq82sBEkB5aUcEj/Czzc9qVWkWyVgClpqQHuYkl9VkOqV1/zUSq9n
AprS5uE7rP7xr6i2QBy4utMUcCyPJI4P3gbGNkETElWg4aZdFYpbiYXQFSFtQBx2jn1fK+GlzpNd
AtzLF0sStmP7hD9B2C78TaKuS3wnYnrFRiIKMb7BHNLa561VChRUCQy6ts8BUwHzsDgndvUZ55Nx
ig2d16TSNwTTu4lzCNwLKp8vQ5r1CcrfsO6vIe6mTdB14Ban//aBXLS45RJ0zUx2+yIdkZz1sQ/w
rjTkVlXkC7NWTUUOA6l++v3NxtR42oAArTQjN9s/5YoCpYOl5GNLk221pe0lADi06OieMd1HHAXS
LT0i3MWs5gsGWYGGWbfCCbJKHpRlNOr38uWdEVLrU4KbFjhyPNukRFZVZr90zsEgICZlg442Di4B
OUTvreLg/YeCAJZCp2Wi1YL2DbotUL+zmdxL8VhSUplDjkzxTqmilHGtei2bXSC0PcX/pHBXEhXN
GQMXB5z4qMuV7a09d7F8eDWDoIqQPZYc3uQQttKiPOGYcwqWfDJqI+4HSl3Ay/qy0x9ra9kL+sv5
NOoZvgOlLwfXhE7o0vuH0BBXiiijmPYt/Yd8se9JGYH7XFK/i1difSau/4iVSloRzVVm67B08C3y
u+NJmYslKZR5qcOtF0oZQKM9YhIkr02tb5mAOA6BuwkrFtbojgo+d0R8bC6Pfdk+i62ltCvL3gOU
BgBYhTS6cFO7i5MKNX7h4czLIbjFJ5/FyZlKtYjawHoqpPlPje5N6wnkIWvNoISU6+LyM2dXPL76
EltIU3ju+cevtkLBxDdpe1TJAt9U2a+sypcIvA0fBCkwNZIiaHI1aoNs6HroKwYcbY9ahyPuoc9N
pYeME9C/zw44pmew7hBHonwlnfByFMbJbZSvx25DZnFfrZrVQ3etRh7Uw9jocA0MM9n3Qkdm0VHS
/Nf9UDwDaZA9esfUtwyF5bn0UqZ6niYn06DwKOHvgsgPFECSNjFpjVmg1Nx2m4o1pU5ZbsrnDrVF
UR1jpyzvhEgYTpwSkjZkRoWkpsrkNIF2Vbb6wF9gOge/t7ovoLhKLMxm7VOObFCYHvmpDN7zbHLO
/jFYNawfNXT7Dj6Okm27ghuGDLHUNIyNipBOupF2Oh5T1udX5hsWmpE3tH2/0dKduXv8ZvexoKhP
i//0NQlQDLS+Ajps/dSkAbDDcwrDSJSk6PEV7W9D/n43fmmaLBJ8iEISBg0xVNdIxxGPzFxMPK4Y
eRpRKMxriA5j6Ygk7w10I2qi9/GkI8ZMxG1g+9txO4aaY79CTmzB8+IChPw/Lhm4MwwaXjoOSY43
JIsqg0fgXss1jRUKWRfe1GQ+Xt3pDLHGIxgItd2cJ/ZAij/GDUsu0ri+OXBU6dwiUcBIWecd0MHC
lf4OUT9xwXHOsmRmOSIx3Brt0/s/qEb56bK82iujn35R9COlTjYerkjLakgmY1aj1VBhLbT3xkec
C3H0TgQDBfZPhSSo0rss2LMuvSSzNXUYcmAH1Q3J0GWUWW5Z478KNoTxkU0cvgNEFT0/hA2W6HM2
/lCG4yHFRHPqF68/W6COVg3IUsCfeXXwcMXXDE4usDU4KfIsCTEbh11VNeMXtGfNwMKP4k2pF++A
1bZ/wVnw1x0D+IWEyWLAiEFMuDN2hRKsYvsi6+1Cpz6wcDWMxVhV6Qffjuacn1qBp5TZTaTpZp7G
Htlexl5tAnb3zBJbhgh58GLndbBWKR1gJywwWwt4mNtu7nFqfqq7W1Z85uPP/yVwR9FrA7PWdfgM
FPnPGIePwxqkD9BXSlhlLzD2jXoC4BtrdmahqZfSZCY5yEGwLlqH5/ITnCh364EHVBW1lbzlOeLY
9b+jwGqTeSun1IGknWE/lV+bjkvzNgTDPCZ1S3hsPelRNm7NeSwMI+v/yovGIJ2GiNfDMDTUQvOd
nMHrs5+V3Le7GUw7D9rWLbwAsVUbsz4EErdqFy/FeB2sd+8BkQooiv63SC+CyideaCrIeeO6vMBC
VS1Ikv2MfbjoASw6cO12nOTGFVek4ZqQBHc7tnmR7lLUz2JJg+/y++q9QeL9JXB4rVsf5gszrtBS
/RW8L6ylBTyClbDb8eoowUWQPJ4RNuBxTkevL7Drbhig5nKDfiW0U/18eDos9Ub68N7VT00A+JrN
VHt6VCy3TqErehsnd1Y6YS46JYiz5111/IBZ7q2pjkEG9Qn6Jw0EeWQWs887iDu2MZ3uVzz3Cbbp
UZ7nZgG4hxokUyMsna4c6C9RCXR+Z+i6p1gGMY3BHWbrqrZuSHBfe1LO+7nIF9IPTm25oLBOKamm
gKlPwX0VHBwBXbGnPcYUmHQKzlJXNNwWwO20ftlDN5cpGTL0sPkagGoh1S7tMHTj4ttHaNmXwlF7
Z0DDUTqDkJK4fR8uZOwRnN/MitUQ/hZ6p0FGb4Y5Bq1IwMlVif9n+pXIyPZxkNoSuyIvp+fs8tdV
DRQRKW1kvLCoOavvH5OCaq3tXSvA99D7fG8lBDTlaTGs+whAE3TdaoI+ISdZaMRLllEnpjc5W9Pk
M02rZD8tPF799NLB5ONOeS+erMyrcJQuRhH2fbi/hJjjTR3av/vo5+RL4tdT0OLdbsGN/+xrL1zt
uyQsz0xbRY/cSlyKmkTtbdrk83hqah2mgbWrkqAo6nVp/ao+XBozPdqkQgyhwerhISXq0altu197
SFBfscBB3TiEkaZY3pYsR9UJeI7bORiqoMFB7j0dE5P+kpRuZGQ7Hgs45FFgXlbNcUWs5RqF2OM0
R06dufxp4gzMns6bM2tKeLHONQ9Bh0tc7/Sr/XQ/eWEcS5kCvXmMhnZ1gGWHbUKd+pC92QP25W1J
KIsBq9FD1drdqlWsfyJ+KXBW3mo+jQmDaPOjuAm1dH+tVGHiPvcKYt0lADFFm+nAkmiOakRYccOA
XVKsBwazO9aItVV9HFSz+gOvw3E45UfL2WTwtg0gd5EL9K5PoiXpAVPvG0LnFtxfbIoQHrD7KGI7
5moHfbxgvm3OpftGRVWPvsZwYEYri8Kyj19zVLFN4Hj0lhCkA/691kIM/XuVnYJ0pKHWl0ougJWm
WfSsspfDtamV8i90UBwcU9CFxL+XKg43k8XWSWn4ZwmKA4cksSoWQcKy5OJKZAXty88HEAtIDXJt
aW56+6u9Nait8bJnVrcdOyr3avq1uhe5ZzTbRFMa3R9eUNlaQ0OMBGYS/jQBRHjrL7P6EUGoxyv7
hfm/vkauVt/ZzFybUA+tKs29TIR2tgeML1gtCoBMInnYidOCfzJTvUHKe5SSROXg7ucBe+wenhf3
lbqNkm9pHJpjJgYG4IhPg4N5+dxIPsQefKftnTq0Ayiqjh15bGoyDNjw+y1247UUszGzIhpO/72A
UwcvUTCanI4LflXTm5G1tXwHZJ6VvNguI/KIM3AsLMYaDtsSPQtTJbnhC7oLpXuPTHKEiowzPXRL
PqRs0kvcG/ISZJQrusItYqQyDl0E2LzimLfMJjG9uuz7h8Xv4kROXcizPF4kyQm/31ym/oQ6wJV0
bY7w9tVCeGAGEP7X2QYYQ6hFz7zNTNH7x7onACXTmMMjsSs3FNm/zKxVDh3S4qknwiD+waiZdfoh
8/vQx+TdYBtjI0Ja0H3fWDTxExu0GZyGXenSUqilQNCic9Sf8T6Iv//TWdHxmP0w/yA183AkjEMT
GsFs4YsE6m/y8ZwsUemiLVADpSlmiBwce5LSmgEVCXFDIqLwNyk9+QKmtHncebDVqaYwKhSwLZBd
O/RMD29qDmykeOGtkciu1onePAbhWsCMT6uLE0pP6QtWSK7ymXYLHU/xPBLRWuo3cI1FSa6Mzqfp
Ia3zfCfp2WdEq6esT+v+kZMw9CpwJ4p2dTyRxafoaOJrDTU44ovmroHGIzkh9+7He7ZGaGikgQ6A
nUDTYuEHI07Yga+Rq/gc9ATrW7MOCHFEbajVP7mwkHxkb4lEYh4tJ+xeIEbJLrh3CD2NKrs+ryZZ
/T7SAINBO5wxRu/t63MZ7QrV++MtXQkqrfuTLaCcWp9ATs1f4vW5EnFWRwXgfuC6LG7JtC1Opotd
jlU0nnwv1dQH1oaYHynuujUnck/OBJHJmWfl4xt2H08YOzIspkpzRLumnReUMeJc2WxHOdVB54QP
8ITMVK9Jc5euorPB+4m2J1GAkFLOEBuSvhsS4hsd3N+n1z1milWlZLZjHrhdGhmqrlt3b9sNPsHy
HvtODzvst7LOpJ+VCzrP1JRAdy5wGOUoK/Rqfq/rTeiaQqSOGvYWqSww6o9xNztWKyN9c8lXHQGD
PZqsoaTUe32Tm0/hPpJN0v46N2diH4G0W5V21VP6xdF9Z7dNwIMaHEG4gVAezYPkPGCJv32knncm
zM+VlHdovmc74n5xlVOcJ6Gk86j2n8IOS4O8kAWopSEdq0T+ygXn7vELm4ZOIDU3XBn9VOg1GXDH
DmbeqSKmfzN6xDkQqJguHPAVrRR8oYokE1TEmj8RDa+HCM0g6/jngdq5ewpmppqT1J6Ujk+fGilt
m7iEieUyL4gY8a3hw9RKwT+Qcg1pmUBM269h9NS1S+15KLSukxj+iAqBHZYdYbjK0tMvjThaRBmT
TN8Ypi4C4Ka5ZRI2+T4uk2dBYyUAgBAKxTP75WAn6Z8LAFrpNvkpRbAgMIepiD9VvxDmdwebSsic
HunADCogfIs6nt3Jiw2VBlzVCwlomist/JKG7zTzxCb08zq/4xfrJTewKPlCTe9hfseG2hbdHpFn
qGOZhOj/KGjE8ZowkpJn4cwXGI9s0KRK1UUIozVcp+NXwPt92nQOcT0ktte16LCFnsJVtw5FXwU9
K3eXgkWZc6ZkJExnsLJPfA2QRmX0i5fCFnmWO5WqN0e3uFWVBROQsCUF19cxFqI8rPzZQzrhcE4R
iJhejhEOOlo8Twn2EVW0diQlRDY28O7+BhbrvODZtGWKv2Ib74uQpJh52ufT++0LEvWFr6dAD5VW
MXHtWbwmLIPTIxrTWAhuDr7+rznbBBPZtDVqIA5vdXrNrvdfnaBvT+0zo0JQOE4A/Qaiwn+9Z7WH
+vXkaWQlx6tv0CsNilR1opXBL0xGpG+C6ZYfzDJPXBO7lpgNDsBtkZRDVKrKZjYgcj+DdKR/r1MU
ftnmFbtHdEmtlEHyfBU/TgYxerV4sx3M/fsjCURIIO0gRUmF1i6o2ueXCL45SHHPS5aElNAeysf3
kG+pmoR8UC/eUdbXuUYM7olInF+MsC0Rq1EGsh5QmX9LCHrOCioHh+PMwBz3E9MoBkPpvysND4nc
tL+k5dAE3zAOODA8MlMurMuxm1rXSAsp84IerjrYCufFm6aN5m/DrblPZjI80B+E1gJo9lfgSQRk
xnoJbZjRtx6DyfUk7XHlRYBlf2KrfNev0r0iXK9RB9nxvzjzGEk/IVrDepLAMZH+40CpB/h/zWML
fwxq09rvEBChw1GKv/UuC4B956TMIaExap9z4SSsk+DVPGwytshoadouoD+otfIIRbM1Ya5cXT/c
mFVgqn9P/XOsN6LnrR/GIjk5DHMuSWvmEoW8FouK9pCFS/ZXyic6NDy/LbbG1aR8KQCzSfy3uK0R
FzG3BhXAu0En+wnhYQsqzhgZZkVqQ3pG26x6SD4J5dQ6mRRZUzXkoSzddKSVP+8+oCbMvhx8nffe
66DM9Nbcn1CuXf13vagFLg5vpEjS+6+/bZR2iNTs58mwk5ZDPNlHUkd7nKjJMvjO2RbR2Dcty7y0
T0A19WyLowUtsSnd3F3lVv6t/58Iq4F9tAyI3ASQDX57OvWVDleea8jAx1A8wAx23kjvqUmYtgAP
28w0QMRqvmRMAyuiHErsWcwlrnTmu7jCs7BsEhbgsjNSNJMj4C5ycFvmSf1VPXZNj+hhTEXRYQyE
2xRROHEpB95i/ZEkqUayCepvTSFy2hzDiq/XL0Ppx5oPr7lNqk4LXzr3s+RSPapWRSZk7ft8a4zD
00QdWTulOq7RNe2q2grtf76AZ4IL4/Qy6INPpp3cEPX17S0+48hGW/VNICbfjOK+aTW7Rw91LIHu
QQGH00GJPP14nGNTl9+qbToUdKE/70yR3EK9VDGPgsB4f6aRGe65kOflZ5Kjrgti1EtOLqp+YmfY
owZ/z+C1gLjrTqdNGpRCVX7luNvPgBgwn19SmY3ECp4QwZDZTRuV3K5lnJs0JaW4ih2Ux2/49vI9
xbXL1CQGkjTi1WHhtKBiGrVDHyuj9+9znBOucO4rKYI0phaf8xZHvjEHqv3cfX+llVIp1UkjBk0h
kT7JdFKpN8ZcyaWBlyd903CDjJ/C1yxtpXzwEILo3ihpdgvxURwRbPjpolCuX66ts7gha8eiQfDg
TqEIMYq7bFaaWl3RzxDk3cWKJXwsU65F79+CK8w5bJ/vXVeJdh19RzQLbHwdLL07OH7YdnPyQDkk
TG27JWXOPmsCRVsejaEwcjbXslJYJ0s2uFy+1Ubeb2GBu0gR5ksr4FzXsw/QeZiH5M/RGPP9lUdo
xNiYxT+YCZnyuA45fZYZATt+3dqTLzWZGA8+BsSmZ5NUqKs02unLKWThR5JBYYbiB9uGbeUrWFJ1
hIcEs6IngiLXOkJjK+Lb8KGUEax22iM/ytpl5tumvWOkrZOKnhw0VRbrxp2KvCgruTI9HuQ5uMgZ
7k4XyUZi7KMq+Jxq0ZisiWqIFOv5uIRjGZigM2dEPvzheP7eNwcyOuP5uzrLCNLFrOxKdz7wLmEN
Wd994d1q91m6j6DWU3oQKzu/nDa3V0p7io0ml0WT49Di9k5tfBRQ120NS7C2TulKoYLgM6/FGcFD
50ccRQJKHPzYRHeuknnReNJp/5KfHV+e9vGylrqa0yV4mK7tSVo9wBvXveK4abuW3ZZasuswxWji
5cMWDuWVweTtKoKF1eg378t9qZLJzHJSf0z/dQdwsnIrOGNQ9fK4aKwdVW/BAhvm9KtY6SlCBc2a
5Ytk6k4eQP/fbRw4ZXAUr8M1Ve1THmy999kopCnM23eAS6ret67XFvqif7dMNFMA/YfWA4Jflekh
0+RZ40IPKyAUG9EUGUfQF7MNEKO7yyVT62qjCoHPZQohTCSisr6A59MUQnalOceF9nBplWo30ziz
6Aiy4TKnKtNjkYcDLZcQ9SCe46HGuVv5XCtVuEz7wSmwcZi+x0Cmm20mljnzY8eUw4lZx2QjyEIz
BkpbiQZK/CiuVWP+zcLLSh/ZJrqpUU9rk3vW76qJUhPMAWAbVWsBs6407z28tftq4QlLxkhEYS5I
Utm3jD4vV9wWaZddC+sTH2dOJhfQqHtNSXy4LxWQGS4w8p62vcF0hxlOHFuOstIUUBkz/45fgGAY
ZTZJ2shy4gUVMyGt3fGtvGRx+OTFLDq07Ny1l0esEoHK8U/madthzCcYIzSLupVqv6k3j/w9thH3
eYjfcOqYIkeG/S8St0WnaUPHDjymRYFSipFcG8NYksG/xa6+BSutF/qyB7wu21pdGwztRRyP/sYU
IWFg1R/luDwLliqqAnd4vFd9E9iMHpKx13Op/TE79qC2yjukZkbc//BzRVo201LWxhlg+vcsljyo
K6X0+1f0Khsnik2RYFq5imhxgvgPC7sAnWocCYds+9IRg6keJ7UQrcvdF6FbEovt2N8uxHYvC3sU
/+ZkxXsuoPne/IH5oBxq+x5wL14kf38+RzwnhP9If/wN7dvviq7uirIm6GkB/PPcDwTArbuOZ+cR
vyFn3OeOeBKcJA0mzd2nFoHLoBY8t4lECmMZC9XlrqUiCkwaX/tIubyt/gB1ots+W8mp32rbszue
icOsFDVEq8fNZBMiCudY+jTGGPVpm1iUHjVNJp4BNwb6BYqibkv3xgNOCq8anaOa7rWsk5YZ42XV
D4nE0idAzM0QRkW2ZXySgv2fSugLng7KA7EruEAWOAsC8HkWc0bKESp5KqVOyVGnW2osrRxCfMO+
7bZ97KxYwj8lhsmZVLk1TqEHwwHcyvmMSnU0CoC10nJMjgXe5EkNL7NAi1e/cAi1bCM+TipMEi85
VIjv1kXEg6opUaYbNeMO8xMcLlCM1ApbOqIvALmb1eRgdS5N6nIGbhCVs4zIxRaV+EQiiqzKOoy5
oUrdjKZSvyytlY3fhOwWhI4Nk4psFeyHe3Ltki4zI3MAq6nZvNKcfJXOug3PcebAr4RtfqaJvcUW
IA/73VDR8qSnc2s4NRizOuEpaXNsbhbqBxN4QKd5IXqqESuI3PKhDKVaOCRmzM9fS6+SNd/FgUne
/NkH4jqEFlnzyotDQMgFOrOpia9P5IRCieWfrIKAmNinW6afkQs4H7yh6uBr9k50VaakAbwgfqkg
YKvd7dG68zYey+FQLZSW13VM+WOTl8eO+J0m2gDlD78hdKyss7MA30ztGBetQ+tsx46cmKBrT/0J
64aNUNiJaelukWFGZ7nFbQ9UI7lkAgUZ2RwtJyLGHWIK7wYGkpiiur6KSTfu/X44MICy3tmO6jFK
RdP56s2FWqfdElQ/iThaMQbjwKhwrFxpYoDRyKt0x2nIURjN/AX4rvKPENlq1lhwn/GuzuNGnQlb
+ZcBjzC+ojqUCL0qjH9uS19jOzVXZclhbrRkTvlUSGjltYl/MOTh2FwsSQ3eMrkfUlLPb5SYTZd/
Jr1tco1vxxqNylaHBoivV6BZUiDrkgUInF5oRJCM/OUcwacsySQS7wxf2Ig2VR4I23T4dqd591ZX
iBTGFa/BlzQQ9SnilllVBNPn2rcNXJuSDGAHWlFoTVb9OPMz51w02h2YSamVUcCga9jpzFT6ETl7
ewePuIeN+GX6HVeUg0ndnW+3+nT9XoZTT8dcNDGyRImPW26KgdZpajADyfzfwIfY+dAe+vLN+YiE
FZ2GZXb+J6O63jMbMOJpM1FNwcaXbw4/6CNeO2UVKOw9KRnqF7puBn8w6Ht/lJxvnMvNORHREqaI
arVAIfdvavNxQ8TifE8jrJxgnk/bjJ9zUm+RkQVvo3x1pieyaynaf1bsrRJZbQx/CC73HCLuGJA8
DONH4rkEtG2KpX9qr5WlQKHpttqm8cVJh5m9ThmlOztFWWqtOc9PZxlRhYk1KpC9OuQtmRV9Sq/Y
eME96S/Ovb5ffjVqf9VrCERPkA+HQPWm70Ffc3itUPBij0zbzfR3EXGijZtWXQYlYVsEfMVUe2hg
PbhW03JmP2dX8aly23o/niFSQqKm0sEsacCLshW7FZ0IWM4TdUy4PVGxSBDHWGJt2bhsRKKDfkaD
jz6loh7+6xGRAIfPriSYXeyyYeMlTORvHIzmVI1Gu/0MMygD+tUTNQ/NkEf2bv4OmSoirPwW/95f
2hfGo6s9CbpyMLZwqvikhGs0rbfELCKy2HWlKWRrY93mWY9f0jlcHxrclopIOUy8sfS6PmH0UwuH
J+NEx+lPzsVIgEegCQB2J7JyXsHMwly79U/SGAgzM1PP5LHjEz411bOqPJqPbuNHqVQuCmPzbGLl
qgnWQrCQ5nmK6QpfXKcV4+SBpFL37ViFR4IbweGD9KC35tMbbZFYVFy/QO/TMX3RzujB/d64cmV4
wvJYN/QscxTv6834qXp8Nkz107Nz9HWI4kZ6ZSg/JEWChHmiZ3XAxbOraVG/YDc0EVkMLyGKMerz
ce6OTQVhi114afX6fzSuusOxEmCtIh5Onk2uYbsq2ZxvxTYo9UGCyQRMxMvkw+CYFIcPtVKllEVc
6Mgzq95HmeAv61NB+Dxi4yz2GL6wrL4CTINppICr6FGoadBQM37+ZpunyskzWAlGGb8aWHyvMC+l
HTT2vwsar48jbQ1vF3vzqJf054Xw722fKRPmIxlfmTalRSB4Rqmp6AdKfDdXI1qlce47uw4dfnPi
cEyE+l1bKzgjb9icuo3aL+ZD0yjvT1ODCIHwoxnPZC8XqWpw7TP4+INW0tJgVqJMd5seaSqbVBUQ
UwwUzfWu+BF817pBcRzD3oSrjmEl//FasPakBMdRApg3mNCIcJZPY+yI4QCtrJZ+q5O7h4AN4T+q
AW92B2MF1WJBFnT/WE6McwQSFNQDq5q0uiPM9XYMxB88rRIaarrQPnMqDA/kPPfAxWI+3epDfO6Q
gf3uzf8Ek/QnFvFoo408pJkWaCeu6Pglw1sE3bjKhLOYgVWhlrTYYtjvpCL6U6g8cefd/wHyrWkc
XG/u+p7dFcocyOiQm3x/D4qE6HclO4tctdTRogf564ErUG8z7rvjq5R9vc3JS+v0dCrt4hPwqPc2
RkOYKjTkGZhtwNOltPIVn5N+DtUM0c9LtZTy8+sREQA1SYfIIV7yvzNtv652wHRaujAtFyVxwhnn
Msh/ZXuDCIoAGBG4G26WtdH1fqkzGJcyFYXrvG1RpPHkxwhbcaxHyGBJqx1VFaLr75b+z7GP1xq0
DrqknGSsozpBDxKTrEVhMGPQ06uITmBoCghvVdeAPY+iay+4FTGTWPMiYcq2xZqhdr4VL03w+5Wp
n08OntZ0nE/TbiGmWZgsTjpPC/DCqwaXKRSxIldshzP4hKUC/Npj1L8tyzN3+zql4Ov7LlO1kM7i
zkvJd9Ku1M6sl+nEzeTslNgCbOpSv9axNdNzsunjd9g9rowoBrzb7WGs3RDy9QqEoxapCYL1U5BU
73w6NUfrnthJRDYHTZCPUYu0b44Z3+gHiPRZIBvR+6wpO5bTMnp70Cx57vwZSWJWfTzV/RoQEfaD
i3M7ngN0AfYnwy0U0VY6uMgyMgnVF/3q4DiaSW4tHX6nMEOsyYiYb02+fcuK2V2XgBVWzyyqyYBU
YJvRM22lJTtnYek1ARF3lyfPH85LN44OKwgmH54z8utSFoeLX0B7PMqvbl8IeZJh3CihZGDmShjz
HN1yuQLzcHqrIT3Ml6mjDGp7CSMA80ROr52yAtY60rz3qY36r6X/Ua7XTRpzwpOOMjO7Ln6HeVOF
Pnw+Reuz/u7/syDk+Vjmk4FNGn9nhBbxGc1egVFw18c/ZuS1rYpN8CftWZ3UGGiFzEnmn+CjbpmD
mkB0hg0VzmMx9e847Y01dnaGBp5q8mWW3mbnV8TP91Xzebk9jhQEJGm7letdKGgQAwDeJDDv3oci
4wv+RY3u6FvOTcXkcubAHTbsWo6V+fL9/ee/La9zPAlW0gt7MgsUKqDJRx8htkkRmEH4kyNTdbWs
gv7QRGQy4VXvS9WIQUk57eGlwSxR8Jb0nzWqRR1E4rErtKhXiVQdwJDQ4hJexvxuDQcl8LW6G651
uh0k3GfXzGb+JvedFAj18HQDB0dtGMHfGWpj1ZKGLZk1dIVdXs0ccyoPt6k5agybcQpSLoC0DGgz
pnSKwzYQ2qFGMqwQ/SeJzPKEU+lXqrZwEKELVkMydmWsbvbw9+162pgrXpV5Xxb+QkwGOPetTMlC
Dl4lUi5tOxdXvOcs6x/c/AHf2IU60uA73bpPO3gt5wyJ+kW2IPZsDBOSYWoqDntitJxK4pAMu3Qz
fnkyJGpLCn/FZq1X3JhwuHd15wKC2g2LgGhAda9eya2T0e6Om+5APIgQ6yCArlPJfwq9j1ZQmHGO
kc79Q2MTiOODUHmBLuWMfhrsoB1p5b6tzYTmwoy8UnbidnXYz7dtcCupYChVxYbxBPGSFKleIOp7
oO+wB8DzX/sDMYoA1T5RsaksyjCjIy54QYPpU+8vQ71lf9cs9d7snAsrRuY9TNdtQjetOgUPYkaX
oXvePzeZ38jr3tYD0+RdbKB5dkySSPR0ohfbxjSEupcf8zCV9GAt0aXv0kYj/vitEoWHuIxT83Eq
+5V4Rmx2U8iFedYsDb/rGVVuuwbkrEADz1vVT4O+i7rkivNUz3qddvJnpLsVuyQhWUw64rsvFb9a
9GZWcp0RIei1SizORcxb+lNSuJugh4UTC99elJoLKAyrmmzL05lZ1zRbNmkFNFfeCbv48N9BlbIx
/ObUP59bv3zhSUQk+s5xXJt51+cE1o7GJtGSc0I62R+02EB7R9ktrT7Jn9a9e6v8fbAT/4rXiVLh
5RZznX3/XU68tjyezi3EtFYmVEV9xSQ+3H7DwOI8krMSJQQlwfKeZLw3qE6bOzXlNPSpqUl9A8F8
w9hz2ATidgbRKZsA1/gmB1KfNy+QvOgBNcsM7JkCjVsrZZRtaqFHnbaQ7egU2Py7T+qxhx1Pxzz1
cQ103c1qrQD5Tqq1XV+ELa3nAmXydNlp8otDCgqQ+ajUNi9T1/6+aJOKOUrd32Wnt5TUEeMNdEZC
z2nQTOzNeEfmOfaVUf5NiSBiCW5N7lYwmE1pAFarA5NRU1TNtp+VrXpgHnG48pmyK/0loPK7XwPG
hCB06QdPqWFzs63gi9vvL+i6I6TFZujwDgd7mta4kaVFllmrbi1dgQJxQerUTw66Ci2I1dfnZEe5
ZDdXvuYF4epV41b3gD9VRh8Mxy6lq+boHIyX2aooSb8GOu4C62M9+F2s0VOOC9ifk5CXGWj2aa1e
nL8VgDWUCRXke+fj6+wOeS7YsFq1lSy1wx/x5x+zMJdhSqrEHIWCCrjgFHy38g0AtVxXdY1sicFg
7dePKA+0FAwahNxnwuFaddWtIZ15XTazOiQBZu4Q5w2JbkXGo4RvjLL4ZGRcC9t0InCzN1c76no3
zGcZRfVT2NWNf7iteEMlDTtOIjIHHgcDT0t2RSMaMFiUv9tvAh7IFJDIYbeewCPcZkqs28kXiqNt
TGjFtezzeF99uaHsfWqyKTLsFeFNoolYrWBpJG8tDTGpOJzT2JtKjRAqoztKXXuG8yWeF4Dq/c5V
4GcLD1KwxWkm3MDqjI4gjHLGvRoVyexNgm5oDGkxiQeEjKahGkvJ1W9UuULaURBhJoldl01vEapf
Ip5wlo6/yA7enAe4E2wwKOq9zdfpbXy8hFD+sypJ9UUUzloESm8Yi5k+04nsUtCihJkprT87vMlA
XL3HNWE3sDQPt7Y49FyZ/xkNPMuM9CJc2tZy2J2l5hvP35knAA1TiXHLZna6RYPgwspLWR2EmVs6
W5cjSZ4owwUB2WwUPH3s9oqvQ87RcH9oh/cBAy+WzMjwz4B8taiXJ9qER/RLRRNImPYwu+ApC1Ud
OjC8gJoQnGeWY+Xtg0KuJtzcfR6FURjsUMGtalOdFlymuDVSn/Vg4X8BmJehNR4JRUh3MLu5PLJd
IAsb5uwLbOxlg7MSsW3bA9NcuCm8y3IzO2JajoGDFZSC7y6CMqA77PavTZkD0C/wM11djrwRAEgR
v/V6h6ulSWDY6FZUjX6G4cBy/88njtppq/RXgYBw8ZidkQqqXBtgD566uTpl+ZdTR6UYRnPz6mE0
eGwLU0Mtz50RkL6VWMFpDSmHnezTXmR4f4bSlQwmwi7roGkHffi1uBXqJjw773SS0vY62FjXFp8t
z/3eNg+cmllHSJDPK78tPetTCpShtkwvTkvyalXrdhB01qc9uIvulJTtNy1scFyEK+Rcb+OS/avi
AJpEcViaNMSVc87BUAp9JVGgGOLVzGahbmDi0Tis3O+mtl9L7u/sY6CajlG86yMG49BB1rYF4g5L
ZNFTyROuH7i4b82Mc1EPXSj2h1FkZGZ9h0t97cRAcfl1NkHvysuiib6WkZWgOWc0IGiuLCzs8Ru3
GhEjGHrrXl7f8hWGVDEcdaueq/EI8xHMo1xA4kXHKnGkBHeJjRt98no5AJus0NObI1OW1OKoOxFD
ykUT5lVSp0XeBo1NYUPWaDwMFVhqgjsBtWt3ooTYbGB/1P379Aek/tZ8+n+9hXLbfXSrtgzLhEDO
D41ufVGpBkVFHlbLa/z1nWRJKwCCRhX4CJykpPuxVUCL1uTF3xMyP1H9s4O4HBzpqmQVE6RbPvZt
8kGCD3AfrIXCYwfesHbSs6R4EL5j4faL8xZ956yuitUeU8QnLuZtp78ejhOZkLN+WMgZOY5LvOXD
ZDkfa2p4YpeIPPwqAJn/DATGQIJ8kjzcVkFHCibAvYlFHpdkvzAhzcSU4Wzax/4dtZ49wlXLzNyW
SZHTDw7oL5cx2E0r6WphUgYfsf2gJU/+VQ0sjZ4vwW1aSGDEFmbvj2dDhnXUx50s+J8Qn3rIdc1q
HeOtGuO4TglGcEQTWCvfdMAGY53TaQcEBDQ+xMUGtEEXyFm77qSG7gxcedtX0a9e+fyDBbdmGB9M
fsX6dufPAR1drCwjJ3OryFgbMcIsH4NHeb8vJY3i9lp/ZWqDqbBFakI4FBGzpPCQddnDq99cBA7M
gshacVq8wKjpzBIf61c3fWWSqYfx4GYZuQFe0EjNK2JyD3fBdml2QrMYSvtsKnq/o5TwCny4aHci
hjdeKmoSp+7sHWl9dU3PmtFWBpbkC1EnIIiDNlPagFn5vUJSvTa51B2hwHp9pDzb4T0XfBBA4sKx
0vYXsLA3REfUDSlIld5lKgtD2Fww9XLdtmGSrSIMVAYu0F4K+woy8DwcQJDJBPMYJgYBVCS9Bo3+
V0x8wyucGd+zaNM0uHpBENCNMDTTiuHLsypBvVCa10n26Gak6pnMriEvMCCUVOdNO+g1Hl7s1Xo2
6dnIZfXxaJLGMiOeOtBfjx6Hx3Kddtayl75fRPNN9NbuvuUGDpff1CO4xr1Ymbt3cDxhfIB+7e5d
5UJ/PM/b4ruY8vOL4WV5gLRFWQT6C2aQqDsB0Zyew5be1uxCmm7InVgkrnuHYhRAsrBowvgRnDC+
6Jf29yDOEpM3zTgACUwVZXUwW3NWgpeALHIq8RzjPAH+iryrihVWO+SWBHYY4pLurFpRiP+cCCxu
AAyhE/k4KrTA8qWlIZuV3qZqLIo+URnqudUWuTGn5RiWZviKpes2ZTdi6mfj+e8mZT9KFnLGvTne
ymc5yngiBZvp6e26BhkZnuQgIVJTMGrGHNin8vaSXcwT5XVZ4WPnIRFA7ffoNfelVwIkUfXdO9FO
cvi8WU0stCvgwXzWrNra3czmLE2EdaXm+TkM6FNjLScOzQoNbsf4TpP8oMyBkkoTbhUu2WS+rRFY
E4pgjp6WX3Yk3iimQhMayUpvraVGySYg36gkABnrCUIiEn/BXkCSBzKSKRWkPHwtjR1JMz23gokj
6EiTFeiWW+NoL9OimG3aSMA/K6hf2qxmK6N9vf0haTE99h3enHx83krIhXnXWW27j67XRa4I6yNE
wwRPxrdQU0hqAyp7NhTJVCKlMNFvWYEjmSH4ksBE6Ho1YyKiR0rjEQHBuXiRks4XOdh9H1KD77b7
e0M2N91+wYxWwFm4pG+lTjgYeIXIfw5G+4baJ34zxChfFdtuBmhnrZNk2KzJgEkLpPf38jQlNG8p
piUCUdHloMnWHrWusxX4XSpytRF6soszYRajUm/AKS9fzD7NX5ZcdDdqx9ZPepZQIMhvEfaxe1jP
h3rcDUfnhivt7rvia1sOjRS3s4LY8/UKKz9sh2HvIJgXWEQYr4koaoieyehaUIc01QzfhI1Fq13U
zyx8lb+yMhg3M79yQFYLAueGIMoEekwc+eZl99AtGaBatJ360dd/6mqCpOhmsyrHgKNfRaZkb3PQ
4aMFFYuxHyv1/hrMNRVrcHPQg+tVXYOkL3oKMv/P2zusA0wIvyVIKblB2nxAAJMBrwJarAIgJgqv
StnD3E6E4LNL5ZVRb1AUVPgxwNz3jAfBY6uenM0F0v9kIXMgLNelxA/45PwOP33TQSCppKX2lw6T
azz1LqILj9tbU8t44fnVTfmt2xfjLyPFE+TBqKCLijA3YumgxSSm6O+jOcIknwINvOQ9EWu+L9CQ
6IQP0DoiIGICdhYJxrsmOcGCOhiJAn6hIhkFLc7636b9SMufSCw+ZPQ7CLf4EsXZvew4I397TZLe
kutU2nNKng/qxIxjcdLps71d0/YrT5AhsbDSTBsryMiJqIo6+VtrC9rk/+2qBWKhj7nVHtVzkc0X
HIBtWhhJCWaNtXrLOWbES9IVojMHTVUnyjvGCHJWWYaOA3xKoxtTfZZHQ0J2+uYmkfIS+N9Ez4SC
AS1ioBmwg0b5YTHAxPuGSiH1nTb8zGXwxTD28Ra/oBeoISUpoMg/Tdh2uJ76fYMnmjQ7yX0id8MD
SigAdylvVUSs6mOmAM9vTQL4z0O92tQf6j6tlHyYqLkL0f3ulLXsvk+/wGku0aQUenwyPDj3+Cb5
Qz9TGMgxqlVFTAVaHBNPmdtpKEi18o9QA/gEdKqDFVt8CheXRKKFOZ5lE1elsjCoJERP0jsY5eZL
+pa76+jzRZ56xl66Z5tTrqV19YHhQuFExqQhoPcNajnFpknC8ZZ3zagVogXDfS/7Etb4OLyfoKDc
kond9mzHH91jTnnHimdGgwCfXuxgXTwEjYC70fevEXOHKH/PP5+A/I28SFfq5Tt264bD8Mjw7Dbz
/neaI0l1MoMaqGB5uOILNXLOrlCFl/gXcQ+T4jkQXjwrE70TTlLzIzbMs3fd373GSIbdW3wCLmwJ
bBmhn5OOC2X9WYbhgFf5EUjq9r70b38OsHwaM2fvf2zLhodyymc3TV59vFSRdOFz28DcV6nIGUJY
bd95yGsc8+nqdqQF4LNHqkmigPTE18fQbjjYyyVT3hXIYsfoXNGz6nGd2MCAohZQuHbDq4zuRXqg
zdOqG4CXnYzth5Y7Nkay710X+iPgOgZqXp+3FyitjMGaaZEDUBzlGpCJQRODj1IG756xywuG0uQ3
STnDteHOsFtoyfCpembkL3Fx/wKzfC89pGjl1xiNc9wB3RtOTMb4ruCpRhn73/hyhm8seyYcx1on
1bXpMoo/dnFNAmPP/nmIswgobWmYFgRI+ld3MY+sxpbsk8l2vkXbnIpSOqKtH1QnDHrqlrpNzTJJ
3IdpfeGOD3HyCJzQG57P5nz0n8PgE1SsWSwf3W8vI9Y5lZeyJTW6IpErGp6eMKRzWnYZncWVyAaQ
t+kpKzJoHMITeALc9dq6CMBGCBHP+84ZPcmDCMOXd7fpsJSzkUwJH3A6T9zlALzopxdty48iD+qN
IW4yRUBJe5IpJvTR+sGTn5B7YR/OIuKf7xiRie5dimRKMbLMPI5wBIlivQRmxlxCZoHfAIeAorHB
HA2zNkPUIOxPvr2LtSgBnJiKcZzkMwXCLkfbAiU5DyWVNxcYMF7i7SR4o64dlNjdTsCO9g3a85CJ
CRUu14gWHUy+vr8JyOH4lOCDePPrme1/ebODpgFSsIpbzx17csIoclXGE5azZeZTUl3e6h5gRyq1
9YOaJDLKdMgwbsCgfK0ARGW9/adaGybwCWMfsSQzlHQ8ghd/mqWsvdSU/MFNFuFBlej7DtirhpDp
CF97LQPiqeu9XFPwBWU/QypHW6I4QYhoXJIHz+wxptwdQNWXxw6I66Rs3ArXABfK3dbYSZU2GXuC
nHRhhpteSPegw33P5ruM8hkxBL3uI3FTS5JrLksXmZaIyi2JlSwH7YADZVj1anU8jZyHyDSJdxfA
7tKPumx3K7Zh9fH57yQxd81OFzNxTkdFcPLEgb/6nx8gzgZhS8FEvDfCAqimjMbkiGqILyhqkniF
7utxxmMLia//G1ID2dUbc0bG5b6X99C2mUscUKk//VCmL/vMBDRZtmkYxYWQXn8d/JizAEOYSJUO
diK9KEey3BZFFlpmfbLPmOt3OhgJQu24lL6oM1aq0Ffy/w4EY0An3k7NaO0CUvDmAzTJU5uqlKw7
RqZUvaIxHJIx9pPWlDsHC/bAnrMUtA481P2Ipi0ChubM4NQTP8eihjZAYfRfMblBU1vxe304i5FV
+Y0kxtDzBvJioAm/oQybrRNpqEZZd3GfkGXjLngXwiPtHp1p4wrdB21u843vpLREj7/NtVcuW4Sw
VbRm/l1nuCBSuvstCMP+b7O/5y8aCs0b0dEimDT0OR2naenh4QeVTwQ7uy08VhXmx9b3769YXHmv
K/wsYdT9rcvcgcdf6ddHNI0BIZbXOSkS66aM7Ny0nEv3WS2hRBvMBufdhXl+cB+E0cGXy50caAYM
XnWuxN9er9dWp84WTdjraIv3TtdwI1PHaHpe07Pvxg7T0cJfeIOvldu+24LYIp4BA8LOiHlRC+kL
y5i7rydEEd2fX/vxjQPUgpIvaMqWMGacE3r/S3OjjRCs2ua/JXaTcMPD84tEjUaDhhhEJtq6sgtx
ipUl3jSQAMZWzjwgt//xYZlQYizuUEGf7uuevNYFxnCkWqZ4snItIm+qwkFXgYe6uB9P302cSk//
ORIOY0YESZi2hxsNCCfNwHl2Ras3zaUUH9CUgK0k8jciz6ERCnASW5RZhxaYnxUMtvCwihznUy0a
zIS1IcHldMOb90Ad0BrKeAscUjgM/4cblEWmjio6xcwRboITGYlxLBLSPSRHh5KpGcSHg7Sxwdzc
ZyxBZ3C2WeJa8FAAC4fV1Edg69XC+Mjjt8leqCYYoRar1dRX82oM0NcCdzAk6A9IGx0HeJ0cdidT
EEoNyFOXxLnO0gtS6joBWaLszyJAVAb19XIUr5is0oefZ3tEcPEnOx8EI5eOrVWnkBBBEIFKvKUX
cPw4HoF7/hT5tIDbuzEBlppoGJEN21uJ3eEzGo43TKAJF0c49lRzYA0o4JIJu62snpsP21Xti43J
tYwHNXqcSN0AH3Aaxxhi+wXTC5WcEEOn7/yMCeUgsTgoogrXTMC9PH0YOJoi9UiubdW7brCtndzf
uG6d+S5mkEZFMQWx1UKiYrLqNzHnTwgnLRqn2NHthxLOCVI/fw6HJBRc852Xbjjio6453zir1b3s
LZrIgnic5LWM3MqMy6yS80Gl2KwEnkhLAi4/xKJqDXw+57m9DYabdJAgHvqxaAMcbcIK2I70M6Ir
jpQb6ZeW+LqG+FgqsK4OEwuT6xkN9UGy5PP4SFycYq9bRhqhZJTt5+l/HqHmpetysP3Y2BzYgOc5
SsVRM5zPH2ZhGza/b2BnzTdroGODIQTNY/ALCg05xKnCMLCctXiDjDu2s36ntA7FOdOYaP0mxBBg
VmUSsLVXwYALk9sWZJieDsa31klnTJE7d0S9GNchibcz3cemLw9Sc6Ser8VhYpU2K5iPW3OP6Vzq
By2b/MjQsQagf3OcDjbEgcVdZJ586O3UtLEoHk/MpdejKB0Ad9kIfgPwd8xkK9jumLy/7+Nnq1Ax
nuI90PI77nDWPXDzV5vHjY0nVv1CAVn/xT2b+2hmng82X6tAyFX1MNyHqABnBPTaWmeWz2E+9JWs
kLuDXupssjihFNSDszQwEEzWAZRDBbZFHienyTVWVAQgInJYI/2MWhodNodg5LITZ+kFviP4jxL4
Movr30AawK2ShTCPo3Baq0as8t6M7mZd9pE7BTep2ETt47tLj+2yT89ePVW+BqyViMWiUXabkHIb
5ecnDkiz322jGiwVwDBupR2UdmUjlZgVPbHaXeCpIGFZ27EyBrSi1ePI0hEhh3g73LuNv9vrkHPn
Rf9EwdrnMzZprAJ4SLOjKyUb+iEt4b1uY6AzYyG5f86l7ZxtT5jXrPsBzLe1iXidiirRNQivucG6
Ae/HIpjQLT4SpuAUZ1BujNVjfpOBqq7RcuDvozee9bq8d+ne26EH/YVexl+eGq1OgG4g6LUZlu5Q
as5kCUDXwK+rhMqPXphuUv56+ZYLpieIeczau1q2Vr09bw2Mebfqy/VZdw7F24D2FGIjaCAr8POL
idNWvWVDuXdexjJOLKFUF3Plc/d0q3INFZ3g9rRE+NcQlCvZNGlrox3b6W+CD1BKIMsQtXGKlHB3
YZxTK/SIt/jPcD0eAoD2JI18HMsPNrDb/4BAu3iwVQy1XmG9lmlEqMxz6oazrpfjPhc05X5D6Hff
iY07AvAFzMDA+stVMr50sNCAv5a8s0DaHc658QREH8tRfY6ahdaUzTSk0InfGIFT5iVGyrUqHUo3
6vtwfU8nginfmcpVoTzxOsyvfyiPs7xfeTZcZOovcQ7QmOpYKetex6Q+MT5dqTmuqf40NULtB+qu
IiF0bVp6IZypWqlFkx0L1Zpb7u90sKV0ewHHIeRanj/QmgcsbD1FxKbQ8HoV1F4XRgnKVzd2PzEz
PlrQ+CawRpuTDBPyyt5l9AkTQAPj2VmrhDGDk/5fF+JO9kLzQKWJ6RnvUa/JiihXROfQgP36au6Q
vh4ELLtaMN7Z8ykMxuWWSRuR8Uuo4TUUJLjGWSKgF6x2hg9exms2DRKyL6ujG4aEv0y8Yt02YZ+S
C402YPibP140j2+x1UBacvGLZGvi9lrbrjW8Aq97pG8PSMqVtqj8831djddHwHy48jfGogsv8sKz
TzLAhKD0Q23OBSUJb+r+LtCqjJK4uPpICltm4v+AVL2LMI76SniyXcc72rXQewxSugeaOARmKdub
xbnChWbOjWwNhdLSwpIM5wuMDoy//3m6d1SpQTQZHgVsGuT7XVSMuopK4GJV6VOQl/uUBIwFOOLz
odNv9V/biGuYReqsMqTVCLyX/2FaaCog8a5MjmXsU9qyylyUQJ+u3G9aN617dH6wkXB4rcknBwUY
FV7JM2K+KP0mXN3rlnBZwBH6MlzQ8u5i6cQfsNRE1gCgzIr5PaGtbWtEKsro564QZPDOYwTsCIPu
CJsM2hb2Vh5vyvVYUEn5brregGWFmCSwwrW3Dp6z7xDF01wmf7N/jG9d4cfnkEjez6WwpA0cQdq7
YrGUmAsluSnTkqXBFaohEUfMnVIffGfELKS40dwvrxwODIXW1G3PaaHb+Dz4LRxEB/JAOShsEWrD
tlVH5IvAjWVYqB/RLRjt3k86ANy0yi6pQMir3iqNb46/duADZRenqUVWiFiAYPwoEb8bDR+zoNht
Obcnzl7/47u2D8IulG8pElYNAQubCSA3E47uZOnhI/HiQ2c7Gd/ZzXXCy+w/tyGTDGBaOZpjjpwg
tKqvY0PaIaWR7r1mXHH+ORE0nqjaaggah02Lz0rvjktekwAjip/96dwq6nEWJyyaYhOoCxWCkwlA
KhDFEPjY1iahFaho4ZfJtzCEZY+GwqZqhjJVPYnBOU0M+TfX4JdT155K8IuYfvYRTNYmsQLsb0nZ
2iM95v/T+/m0wnUEcjSRe+BIpOMT+DZoAbU3iNPUq5Th7w95O02yAsmRhVJGbh8HXcEGhl0Cc0N8
injsKZNxPbliQD3Msi6bskS1N+RwsvSJp/9nreD44LbZhbCJXw0fV+YK3LsztkEfEXRvrsmdMqPC
I+ji3+iT6UN7ITxtdBEZQ8FEQr8kom97jyJ7cHX6O9dRPq6cES6fZKWW7lrbh+CLjttT54Pi2+rW
lgkbfhYA2Y7zg+aRCGpDeGqnJBkTU2gHM4GKDbpkoQSkH+g69Y3s7jkYief6D0fvHfaF7uDqNbCO
oPzb1C9QoC6S93MrIQX4PM9Dzpbjj98Ev7lkWSpRyNFj0rpl8ARmyoT/NoaNgMagYz1znedS8z7D
MesBHuAl4PeTHc/gYW8MJ2yQVFiGXpP+QEK3xiV+IgHB5bK5uHopSoaLRP65chPZvLvGPgYQ5gag
Nn8b2aYYdpmBw2lMAhr52IV9hI6OwErCkQaq72FyktXpSCv8y9D8YH1AHBRsjDuvvGWJ9eZ1sbla
vG3HhjEpKF56djUaAm5Y/L9pqTRA7OdmE2sc0tYo0WHotSZbtu3kj8P65P3sKfe2NxtYggvMc1be
oTjncfLl738S5iaaxe9TVhsXjWyr8CFbVZJpgcPT2ZmTQYg8zFbDXCFBIJ2YUgUoajh018/nNwBL
p7170xNF63qgqI7oqaKi4yTOuavEoV1nqkPhAWObUGrUS+B9kavrERNtTaGtjbVpo2FFrf8qvoyZ
jtWOQhr+kwslLu/a5Y9Gcdi5xwBnWg4gaX7bG67vA+oySMP6O0TMk+WiluOpHFFw1y8NNPr3XE8F
KPUcctCXHI1VROaDGh3bvd/o7H4W2JBT8wcy//KDxPZrKU1VJa+v8kD2tE8zX1V4qEBwz43uEHdk
vMi18MvcZKUTkU0ziiTJdJjyEJBK36oqc2WjDbNiUrtLcJF1j8ZpMVeLjEEnR8FHPArBVi7BStF8
+xsQFWkCFf+CloagBdkgzvKbxLe0Jma2cpEiqY3KENkrP+gpCgunZGieFhE33dAlP1ReaHgSuX9/
ShZVuYDgzxPW7o8sKxbGgy9zvmUB0pnxpVHV4eOsvzRXGsp78DqtylplLg14xqOtlMKSVLLadjsN
pT0/BCw/eoyz4+agxfjIJpoyHICAbHoHn2ldyB4fbZDmE2W04uqpZQEUov+FB7cfPb4akbeYUdhX
or3Dql7Y84aIKIieP+/he7/ZLvQCLoacBo39ksS/bCxpGLUGZW6OSP3t8li9k/VL6xwfjRytJ/Za
yAS9RS5ZFMrW9O9ajEEvysciPz2O0MvDgtvEI1vUHtCnfr8iLMksqlpP/5RK4Gd458YI++q24+Ch
3FAnaFCZycd1UNbD2ektJ7tkhlqdH6Vlaj46Ay50DO1ck6Jak9U2KS2Q5hhHTsjDLVIxwjKyNdju
sVz7rX+3aMQiV2X23s75rZtYmavuRfw6RXmX1tw3+fFqlI4+X479cc58D5pGdjYlMzXCajQ2SA4B
7NNBnsC4MdPQzVpTVEEiVSDOqbV9dVZGZwoHtCTH29xZ3g+YwxrwtzKslOQF7k4o6asA9Z141lZy
/8nW8gZYGTdF79yukOC2uNfJDzHM8QbEJ7IvfjiglpaYOeYqxyZiERv6D2JFAa8qzBbI8olpc7lN
U8c05u+1tlRzPhxTjCbPb9WI3sh+sPLht6aOJosRkpw7gyR05sFsXEEFirT1OxzmD7LfY+3TOuD3
U5JNHAJldaWvAg5fJNjjZiCkiAJhn5+XZgyPdNVaNCk5a9TTsyeUgeLr5sQLa6yq3kjx7fh+qEQ1
8/fa5N+bRp/F9puxMXZbjeODQixTgBiGPTKfI/PIgBvwKpa1r3iY3dhqIPN7/0VrJHM/yfCZnaSs
owt2HLuDCmVzjJilHYHHF+BzeTvyqp9hnD1PP8bAax5zAiNhFJmycbmCqMCR+A07qCxv7xrCezIC
D+Frh2KvQ/VBevfcmjfby2S/AdPAVC/WdJzw/Pav5R4gy/6x3GIH6zFRMvTNoBbkYk5PJENrbtp4
UUukDuWPEDBVlkTcC6eJ+obuQKhjw13kk4EoAwLc7ERDKtGnAoVsYssTAoIaWf5WcWxRH6eeHGeR
Gs7DrNzlTb3pLhv8ezgGAYM4TmzJqOgVukNQ/TLJ/L7yVFJ7hng7TO0v78pm4kpa8v2+gziJ9p8t
0jVyu7Hh++CFIFUjjriGAuoo8MxynIxB/qDv2+X/r4QK4Dtu7SQU8jgr6jkuTxZMpDkWHHYyDAJp
78t1kUnz6u+xCCos6wxqmZj4Pu0AKemcrsYkyczvnot8n0zq/CQHiRW3OGcIrRdEvG7FPVh8YHVb
vJYkf4wN/pAe4xdGer+6Z1C5IH/26bqknx+c6tCgd2L2NCRsdBw9xG51EHQ/f+udfgRT0q4iOYG1
AhfVQv5CQVKAkbm7Ou5Z5vFyhSpFymUuvCIoVnd/oB0X/e34ViQuMV708xT5k54BqwpijFOn9BAd
zayZieYBWzs14e/nfAu6ObjOwaj49X0IdfhYoknL7x4/yBDNVk62lWjW8LQ3/RuUtHNENbQaCoWn
xpGDlj2l5cV+UOFgznYyPBjR+uTT9/fWpOZUlffkA/DrvCgdOndbR6SzyBGGSiwV+kDdoVA8yGZy
C0AgZFTPaFb509XPF6zGXdFRBHNCBNtvjuSd52Afw7hC+yOOm528vWV4Am+cGlUIo1E5HOeUl9Xe
+dl4o71eMP1UlB1bDO+IkN40eurI+bYz3yHS3WIzCKZNP0RYw1rTIwvxCO1UTOm7aFRBtadDJw4p
L/usgkgtz2mEG52+Z8tgHQrvM3ZXExdS93R7AEWxvO8gv6tD7gsnUve97pJL895RdxKUuLbFZWUF
2bpMGNvpj5z/4vW58bhOyQlleTUNhub4WNDXpm0q82AMPuMbcFn2jHCr1RVJEKRyejoO5rW9Qdkc
z6pBwT5lmh+kUQLsiFPQ0djaexKHd1AgTvjJQKx7EttFeg/k/5q/5/nVQWc50CcUVZ7D8dLV4ZqX
jmbltRpYt+IuOGq4QfpidN+KxT1dQjkldfxc3HXiqiwfBifERT4Df4sqdzqCfwqo7o1/OipFf7cE
x/ij5ywyNDKFWaFy3mvN6sfOREIQ3JTaF8+l9OxXFbcGmtkwk57LosLNNS/9N1MqiDkHGI5XPQlE
cOBuL6FD7TJND8q1TNxThuWOvVwbB7s7+hYXPAeCCXwzC2yl44uFcK3qKes1H2x5ac2Ve+RKYq7q
26SMuDMEKBIOxICSa3jAYjHggt2GGmqU5TOkqrzfMlO4MORBUdoxSP2Wcox8Yb9lsqlsuF7TdeNW
5oXFkJLVP2CRZ3RF4Ja6ezZ/JcraZrdRKgiHYiYO0jlhhmGDTfwvp1sBna3JvIhEPEA+65DJqU4i
34btVBok0VRCvg+hWzWzT/Bo/WsZZlQDenF+0715a8ysLi7elKdOXwCVYrDLcrZNol8zJ4sxTfwL
6noLJ+e10kUKC82TE96W1r928Kmcn+qMM45aigZkVf7d6XnYAdaaMGgAxiXwRrMSW3rdmBeszgxk
uk209DljcOyJSxX1Y9tWOovOQUkUWgRRasNgafC9jGWjIfKDyxjThiMiIs8SFLltC0mecWtsT3OY
CQO2SPQs/VxABPA3Q1vjAVVsMqS4Z25aE6dROpkPD1GFGU4oYCIQvrj9yO5gNY7HkagxeMl14zoM
gmL8ECgPimUNZBMmsV6I+4mZZr2mzjuHZ0Q7ikVB056QoAgGBExfKHa1/ic3Ib2VtKEUf+TnSs35
ku6xcm8g86cNtopy7F4pBeYHZ6jQTvqWLp51C6pZHeY7zx4+t5CBj5WZpHSK0y0vch7QAHXt0UwO
lBRn3nTYq73qxOaqEm0JMcEHFtdl8Gu+DUL7xVwQNUjSIvTDBz+Z0d1cYe/ow10TKhnmDWZQP3UW
TnFva9RB86vYNjEi8SQJrPsf8WnwdWwBjl27YBFWzKMIywCYo+hsMv+aBnnR+oQoSLHuDaJdVYGQ
5Of9IaAVm1MUxfVMhh6/HyS6k+FZ3x7/3iw3cemQB8SFNdM1gZ6+8VRKTyP2Xx9ZtWbtwjwlZ4E3
n+ju35xc7yT84zSOBvm4SySOyCYo+NDKIznwjwFiF/HAXwxsV0g+Rhs06oBB9XkIW8c0AHmW4P0w
a0/rw4rYaZXt/EI9A49sK3TZea85OHTqn2Ipx9BX/MmfbjABKtaTeUKcuJpaeUZ2n6Nsl69mlW36
ha1Pb8FD2bDZZreJsWUKz+PEVDD/OOZmGj/+XybxrZjOikF3Oylbk8evm7fC4NBbVOO5WDT8O3eq
v7pz2/z2PDC+zoy0vV76RachqjetNLC6stWDVUmScO6ne5aTEDqUIHJ8SQSXbHiju7kfFvd7UIAj
w6VKJX5JXLN5xKg+McfQKdxtU/2DpgHsA6x5VAwdtlksrHetozluSHm8NxbRcnHflmCYHlvOJcWn
wYMR+IeVJHs+X+av+VmHuXRBNwKFnZLPGcwUyTNKzXoH2McFvFz8zSNwB6xytkQtoWeaqiNKRZqo
c8Ch85hVkPpPV4AKl0cY1+X0NU3CEt4RhqIh8UZAv5JO1lgD95oQsWFmaJBzDfw7v00GNLF56QXu
7oxbbIEYsNO6ObHitPx8o9Y/nhZII8N3cEa9ec6I+0cmwMTyZKNy3V0ZhSLbM1uSyspSqjDYcxWr
RAsOmaRb0sqT2K4HQhyQLYRvHQxFeC5rCscnHLtHy8wDW0k3Bw76R/yDzeF2eCIdoAu/sWs/LkXF
gt9OoODbq49w/bD8k2t2KcUsjbHsUb0b+/O8pBkXg8NRnKObFw3JWHQH9Sg0OW0kD9pNmaTm3hyV
wZ1m9RVO7hCn59WxSw2Iyz8PSNUgeD6Y14Qy7Mer4xKzS9V0yVFFWkwICJbJdVwg05BG9IfBEOvV
hCxMKJqqwxuw9aUEsAv6jjtIUlCP15UH5/N1WZt59Bvjsej3xptk/+zBSsK9NU+UncfrQCHLvBUO
9Ls8uJBg1C3H97EA/NvYe9bNx74JFbR4crr6CM/G9bNbHXQcvIFZU1j6OFzi9VZirWRstgCFec9c
E0acnb7OHx98RhfurtBgZsGhU64RVDDS7va7Vn70+pww2sqm3UlvClNpUITlELIhz/RVf2Wldg4l
BXwtLoBico0leF+rpEmxrNyczP+zNbNTspXcGnewHAYj9eQJUyixLDVMSWZM35M64MZb2ic7MFGk
X0cawzgkr/uNb0kPdA8qGkjwyxxJDvnzS+ZnGVfFafWwCiqjnntgEJZZeU+aCTwqwQ7p2H8s/SWe
oPlB550ObKqDD7xW7mGabVYOV7NCKEZBYGXRqDVkqHA47IjzCXfapfEZmQkSYANk8TMKM1wkY66H
67iRGOvQZhhFoMixKsNaFiXrwFrHL6ceAWnC43qL1rGthIvEl5EefxfMZ4+WiDno6MXTR+ga5riw
UyjxEC/enDkxCttb/oWWqklK1ADw7A5471KW6JnlFKo3gmpiccTh0r2yQjZYq9V2jPX7Z8dYdk5h
aV6TcfhqofPyebc1IbeJ5/xzx/HuvHUfMQurkdF7fuh1ygZrcj6s59O9gxxwD9GQiBv30bF2fk+d
dCH0vO4aU6KqGKibJ1fnUHZm3yUO7XD4/E3SGYOinkFKjSuBSsPApswLp1QSWOGlZvXRb5a0ekuZ
STz6MyQgZuNCFaObmCA/c180FwAzsay7hdqHoT0odOgoUcixy9uPR8tpta+ZjqP9Ax0e3GYDUqhH
i7sJIonTc0GeBFBLl3IDj0bx7FPV/rCpOuBqQNJLOprK03mztO153CogRLfBP80yP2VZP7tanLpt
9ngcYyGUyBOA92x/4ieAeiAvafVLpO5sJzQqA6clYPMfkW4KatU4SVsyPrkf9GEp1jf5JVbHcrIH
2Cp2atrYWYVDoT6JBnjaTrnbPZrnLNdPv8Lw4d9AW4sZ4BSjaAY1ze+Gw/nUcBv4Fij/9T5c937d
aIoC7PfwtI4aQm/2Wx6P0PivIvOezJ2DnxFtQnt6YyQ5wYfBpngoBC9OmVjWb2uv2m+b+chphKAD
sy23tv31H7Ogv/vcnoyJB4DnbcBz1Th3Kpi5O53OITG27qV06wSJ2wLXyVs1UN20Sdui0YMvGEMU
ngpUD9HBQy6ju7NNOt/8SDG/V6tjs/1zmpdjVuhn/i2MWDAjeznAlEUJgS5nq5kUWYC765y1GOw9
4ML5h2AjKtq2Kc6kKZh9oAinQ49TI0ShkqPgixuisGhJj/bo64pM8aGygqejhhDHL+6RUWIQxWo5
HNgH/l/SF9sQMpGnx1CknpVmIL/zSuN93gJBoF+EUh6EGineqKfFvg6E77DY8uRnNCTNcxsgS1vw
++QIbA1hJBrFVE7vPtpzWzC6n6ieVbhSfA5hRwpKTqPIRLla2ISahjwbYO8qaW9ZbDqAASGN1zQH
n44BzxFf1MdgJkCKfDwn+peTbwUmo1OvKrXW2KpfEVmuw7qzDbDuP4BNJlbjRfpU8W57IRb7YsPK
eMu/6qCL2zJZL2cb+DwJmlaHhKHbrA1lzl+UY7bsmMg/Hc8SXBqAuixj8k9XDGK3tL8lKu3Ff3jt
WyqfY1misPyeAc+RaDD1xHCTvu5NgWL81IcgKMqD2Qj3DRGhxLu64jUiub8x33m5fSk4WZ4h8iwB
vJ11QCgjA4xK2lNSwTUtO22QcWz5DiKJSUKMWTv7FvpLSsVidLPGlOixwvhqaqNQ2HJH+wsk5fMZ
FQMmdYcPZia6Ju2Lb/9dlixxkh0XdNG7lgzW6DpoPrmoSrTFljGkaQdzu9/xOQoSmHOzu08daZar
SbSe8QzVr0RUNmn/5PwixEGVVIAWsbmvepqpFvC8ufuEz919r+rVeq7nprTrfwIyWZVO53NUfv/d
rG3g+z92jw0PYESdZnPjUWxUSzdLXhxqDwYn3wfrEWYxsq3zeToemWiW9+kj/7/ronyjmj65IqlF
GHYU0nvXvNkvvAVMb1rBHmjjVStS8IAXwyRyd+Q1/FZsuNIpQKWpBot0v1c8D9FBnRbpysDjZtc5
F9yTHGqT4ZU6+ILBwKpvRLsuVrA1nxMzItU11kEHp64zxQIZfP9G6MeD1paQeH1KAigz3JdxQPoQ
/O2BmiT6spIssAG7MskWSKTlB2U0f58+R3dKepFZ8A6Kz2Oz/tW7hEcZedIYuoSszpJvoBXs6zLg
8siGpe5OjoGyuL2/VOdtPEkKji+5OcD79yaktECGqzJrvUtd3DaZCNJhoTJhhnmqeBwR6Fd4gvQB
dp5sH71s7z/yokeVFDTirhhCins5jD1CPhKdy5rbt9TrUx1IJE8bhHCp+9oNuGkawvsgus0am5Ib
L9pvwXpOar/R0+Fjy/DAIpzJUVmnSilz3YXBtyV6eJxLDJVIWo5MrASGIr60aRenYq2qdPBChsR6
WJZ5IIMa/SsubRW82n7awMCtLAJtbyKzYmfbuPxWrjS5ixn7fq/WQ0u2QQ4vuAdK7+SXtJMktq4/
hxspOEFtQtXNJF82o/u39xr1C3ZO14odEQlAdI3+elkm0POMMGjhQOFkPSmJqbjahSe8NmlJjTek
z2YNe2pQ8WdwEAlXBzz2PEDvhAAFDu7z+r6OwneOqFu8wH7KcbBWHs6rbxIiYfAW80RZXFzQpFoN
FUc3ySxx9N0rzFqurLvc2TueNnGADyFXFIsOwd/AwhRjrONPK5UV8fsGH5H4lGKwjbRcyYz985ap
1144uUvmeShxN/3Z25e3FN9HDI9qnUIj+K5zgj3fBLt2yATqvLpkx6aoi1ILLP8b+1QRRcGOyi+Y
u3umvFri5c22+huaiy7p4834ZLFm5ieVSGuWAZ0PSa/jriZq3B32Y8ZBEVrso8bErwwDWA19cjSz
95S1a83btGLGjz57q35fMToEpd9RBAjlTfILtYkDdDH7tIl6f/+7tkpONQuD33ePc0olWh9YwtN7
q2nWjy52N4A1vN0sLQyAeLhXP8HgTwyx6XAjST88FkgNH/EVZnv85vc/yLeAHuu0zn471NYIRyH9
g+CwsVxZtMVEmBXYhZYUYdEvLnPkrZYiejSCZMFAD49pQf6NkDIDZoAm38eL6xGQodyTlUYxQ8rr
riGdWMMWqpqUBR2OrnTG+YvII15DmQKpnKmcu+OumHFTGGdpo8iQGl7CIXwf5xhIVgq9b26HGS6x
AY/v+Uz/7rCzFhvo2mcqMQqQJkTIb4eIlFBN785oGRQpoQiiSn6FdXhabSlrs57rsgcw4FqOAVkU
AP0EElLYVU0hZOds6mUi+32cqTbK2Zt2x/zW76hROTsbXdnOFhGGLY8BLC1o+henqQOb2wQjRIPc
cUxKF4srxT9tSgytqg4Vr4GZMpXpXLqpZsX/NhIYr07O9+n3p+EHslKQ7QUod74gtUrNhyUeirqX
CIXC3IxcdEuY9YZjIPkw17ViHPLK+TsZa+5cSICbAXPukmu/GPbQC/GiDq2HLgUnXkbww8S7zyBg
vHDgpBdhk/b+0sHc789Pc9wcunWNyETvgQCSQZuLfTOekvxeSwFhri76fUE7Qav4gdyMJNwOjMgu
Khg379DEF/aNhbuZHK+/+8sTPFZiqP7VL6e0NML7SJi09n23cQyVT91W5EfrEHIkfA2BJLSt9ezp
BeA5w7jdeiYjXOlsm+4xgfdFVfS33AjQfi/qbOZSQr8y/3/MF02iga6SiaioKEYSbwS65wYOXdt8
VQX30DxSr8f0Ja4FiNE7LcnAeOXdMh2gYzpB1Vow2b9XES8QLyFMVf6ACSbNzKNQAcxgaWb369H1
w60FSYy4TOcbCoWuNAq4hvwkznBn8zjjdCvkY4L+Un6/+6EjFtxRWMp8e5MfFWmson0WnJLT0a9J
PFPoxxhsFhe+oMB6h9sVlQCIpTFL2uaIpEy5SJxKvlicQCC10ZAxp024KMFhw3ySPVts118eWSXq
0AItPLFG0rMx07zavWK7PHlscqD617fnb6N8o0NKUk+gdw7I89BTNKFp0j9JClW/KXN3G84y52z3
HUmtFOk2CPJHxwr+n+GohhCfi1sNLPUDVHCPl8asnatCD6ybb2unYepNeGLIETMVjHX0rZxd/xw0
VV04x5H07HFa+3KBXX7PWuF6kCCYMmRAFrqAVQwznXVUZTX+XSzBQGawwPGwlO8/QVBOpEogi9Xj
n//17ADdYckWV3IfE4vMmLuKTGhF9mw7R2ChPVccIESOW5JuTMZIlvHDq6rI0QLbXy+E112AHKO6
eowr8uRs9jwsAAUtAMFMG1SNagjO+XZdNuoVp2rUCoudhiR44Wyh73H9p86ZqWR3xZXqdhx9WQ5u
sFZem01tJRa+eoY0054NdGJsDfNh+qSoz2/756zodWyd9izR1CAxDbTDDUM09By1layb6t2fo2pA
P+c9MqCholnXl1bgbJGuLNZhXXbwKNn8e24LfzDLM5tFgbNazrbsRvv3EJlJBO88r2OEEy//eHfo
z0b8SkX4iI/WAwi2TsANOQuKNjRakMSPBWOknZEJpP4nEP25Py9+0yewQOjVB219LtyGEc1aGOaC
KDX1UIBbn4enPigr/DEmIBpMNXJi29JITJWoR4kc2UdzpkkOcs4nX6IwjyFSX28DRZeHvP3xBqMs
g4PsIhzRXWB7hPTVkjnBLX0U5sYkmT/J+1fFxDZjjYsEmHdH9sPGTSVX5wwj9bOcbsbzeQ/7yIOa
x/oBhzc2XNFcv2oIXOKMpodCYXEIu/vddS4c3aceaPHL9rbyql5nVO6taplmWxmMwkbOstqS5JXa
AupmLiUjip/QQdTZfzj2RERM3itIX8dx+UWqZbNRv682rl6A8xeGWOKdHwCgwjhEMxyanACxYeA+
x2wzy08UgVuM5YJYh19CGahHI/CbzkQ+JSPaGkOPhcPICHIlJmn0FTckj/qOdbr1uEhRalq054oP
SuoA6xLfEB9oCy5wQGHACZH1VXzkJ1KWewEYnl2Gmn2FJ9eLjCyFSxKcB29V3lHr9tZqJEI5bdYr
MEVFRyR/5kkUQtTfBDzKx5MMsGabfBrWhY+A3RZtV+hPPAZ1XzsVv6ZOMSF9IkRxFZJSNlSRJEqe
KfKe0jNlHxDD1VVgNnzCW6/h6vaMEVMoUPXa/sayqMkeht1INln7N598hbVHbZgilKsp1ZHNnOIr
4WFDjZTfWPHqh8um6j7jjDgf1nVcp/QQ7bAKeidxrLKvHrksiwmAcNlj6Mml7LJY5Z3wkONbmO2p
SMN71IbNw6oVZj57BPrjodlK2JKFDUbdDn1xdeLAjN6KUXzq+Bbslumwil2w7kGI/rMJNhzRrLuF
kAGK0tXY9t4wtgEMD+l8SaMu+FR/A7LBa+Y5P03ymgQJeud4V/tLymmY2vRMUREneHlJbhbXOHuH
5Qb2cLb3R5zZZ6xGWH0o1/cXdRjt+0wV40Dgh3Yy50Eq5z7CKgxkDldhB0gp07SJFVqZjXTqRsis
KmhRf87AoKPNYQikCxo4tZKylNf2ogZXAEh32JGO/5N6C4o0utKulw5wQVbseWIbxNn7w/fUcvZY
oh64IfGwivqpwSazsjHW3KO6NfXQjXPrwONmMEljve5YOnOsl0Kf+jiyajXr/ceaxdU5XQUTD2xo
ZtpVP1i+XAt3CWgYhHR4K+ih1nWiIkSV/maqslbQsNFnXUNp2l5s5QhtC5ADFN2AeJHN0mD8WC28
2FKLaa2DLvCZJUfFf406AcW7WwTL/vHcDmindiDNaqkbdu8dYqYvYdWy3NBjwjN8Fp+HzCgeXbV4
20HhcX6RolXCytWuJ9xTWv8V2sJ46so6wPTshqRENXzoyUj6Gz4AGkeUJqsw8e275TFF0LJOErmH
jsdha+yZJQiLG3PsNDfkpDuRkqCLBUjiPMIlz7vQwnDL+ktRaVkH7Qop6qL0kdaEy9mKedwHqX5Y
gr/7ZnmItuuSzZlJcgENN1/i5ulvGLU3wvLPU8Xnbyf2ZIOQRWSKAQCgJlTM879iA7xMrn25pJAI
m5KF+pVF2J3uLcQRAl3M0xRFP73n0Z/3f4ojq8Jaqpe71A7reUbIoAyAjLIdlhfhzmiVUyEmrIpR
hWWZo+oaMd68jCZziCGMVodiVNkkq0beVySe02LeTMG5mh6MIEcdNr7cIQLfPanlNaprpJUPJcbv
Lt53SZi/YkLdmthGtFVgyR4iUAuXML8/atxzwMD/shL606PFuVBbydwuH1dYZ9ClgFQrxeRy6i92
wM/pW4AcYvpX4IfZoJFfBlNcBWlpzgcdsus0ooCdyqMMTAyl62uhu+PCQZqhSLuKYV1fg2nCooMC
BN54QsDw/8fU/puFMaeuClQaWnGKHy6vAgE/EdUz+8W/Dcr2+ICrdZZFWGmvZahOPt0ZDYljqS4J
4XzJVPxqljRk5t6Qe3Gc3RhxuM4fmfd56CnB8tzZ43SmMcvA1PoQ4XngwEZd28moAkr8F1EnveTG
ehfu5dCEhhu4KvTO86MoSI8L+hi0F8inf1/OSCIUUAoVj6/eRLFESNZ0lkL+DNwvUf1B9s4WsFid
9nvb+QsQm93iNNW9Jstp5SpttN+mdB00AahmxJXkTRCAGjFTAeI2km/mYOKhblf8Ohce17nmPBkI
g9Nr+RcfgPL/giIZ/5kMVpYqHIieT9i6p+9eccpKx+nQbixZdj0k678BAuU16yz7BxrEFERn65Nz
H0wsZ66Q0Av+/FTY0mubfTFYXlWvDPcF2ev1EQGy389XgZx1anUer3Vqqx8EXLmTRY3Vt0bRYf0l
+G48jCLo+HlWWO/jc50oSiCKRXqJYCgaVVJ+rdOJNNKdFhOW1gYMV2BNoWljHPtEuVx7i7IUD0jD
NKidkfOfzCC7Mx9JH0XmSVG86/f30dHnuvL/1HrwUDPNpzwNN9pjmXQHkI2f/kzCe6uzk8X3M3c+
jV0XmyGOL06Sv6N/zc/DcUJj1yG0qKsrCkz4NVaqVO9BsEeu5Wqy8DsUBw9Z98ot39i/tsrkkGHR
X0FxxyHBZGoOZhxf3iU26nUDaUmYOj1pMQ9mR4U1b4hxuiZO30scqGJrrJ+tt00ZLqbbJxn1ctj4
9AQp8fMaeCuvCkSVICW1kKhsSYU0+EkKm0EKRwOx3SLDCsxYfbZGQmCRfLFqhSn9xzFT9SneMb27
csc9mxtvtcrvjyolVuIe8/zisddJVSo5Y3MBrgd+02VTnHysEnfQxb5AuX681io3pdAG/7tloBGm
wzQBD0E32SVWra7KUQJqIf64IU/h0Ez+Kwip0ABirMaf2fGBBJnyeORbCJUT1lhQzW2IHA8k3mhL
LTLQGm2Pk+kuc9qkIErGiaKhYy87VkoJZHsk3sPh0tMSyVVm9t7jRDBzdSmsac0QccMAK2Gw9jnM
t5WnSGkGFcanYZwr5iRHJlBq/2NZwOHqVT7379TtQXxrJvwEc3n5VGe0UgeaqP6AgbowNKN+qqfG
uf9rYF0lu9sfMBH+LDcTAxpeS+IZ8wItos8/Td2ndRYsHzpzOWiWJo+BYP66FSX89TkRospMwW1h
5lht4JFNmihNdpwSU/1jdbdgTjOxK/pkbjLjgTFVPqwG1BW5Hgye23pRk927fXs+85uwbssnHe+9
BE3HqTow2bHJvbph7OlmaMX9votP8SQeEf4cBNEuN6rI+Wcq5hezTVlsuQZ1jIqvVlrTF/36cy/3
1BJ4HeTnY/+ui1lYV6hLFvtjBDLT3Iwse4CAaqeoUKsWFzY+0nNzeSft9CPEGcGjXju58v9APLs7
QU8ApHXYRoF0e6mzggiuabVDwF9rN0Z5XlnTE4ciyiFmqJxAzTchpKAPqkxWHbaEmSdJ+S28fQsR
rmAFmHf+YeHkxQl39NAaL4uRR/RYzNLaGNIvzQD3Dxgjyr4PTTFrA1vzGX1oxgWbE8oa2ICzB9TE
VOrtR+C76dhUJ1g5vsQRGukyZkxsDHr+Q5kh+kBmVxZxVW99ANOSxaKkPtqc9HHdSNCzI81bZjTv
nqADFRRqCBPLYbnmaVePwVHK0n/Dp0Qkz5ZrUEQ7W5593CX8vXla5Ors+0WY+xHWnNo+k6suJ8Af
Y9Z948cbalBHJ16vXBLk8g2iaARBoFIE1uz+hyVzwxPRsvzx6mWxzL5c+diZhQ3ZXvgqbXjUYqim
TxRqkTmonZNtf8SEbFl1ndi3GQQY5SxZ90DXwRRZLtbtGT8zuLx+2Rcic5dt6XWiSEJJYDgoHvZH
AAN0m8WQwaQHoaadgLtNK9za5aHxotJeJPsla1z76CQmliClR+um/dym7Dsm5PKkVsWLafFnUDYm
iDpY9S//RDmE077BYrsgfO+JyQC0fBpIj8Hex8OQ8KiZwEQMSsgVEz56kXV1RNMNNkpSdnM2Wo4a
/mDeWrScuh5BNYyMnz0zhDlxqVuF8GmM/8ei2Zu3JQj1mAWSaCuUV7FWjsBXrjPnV6OJnthUMqYA
XXzdzpj1/o93dJ04Jiycn/Y7UIj7y6cvaaTY8eqhGJSHvM1lz9IbCNMrYNQdpIu1QaNf2ZUp7CIm
R5yyC/sG7s3WmAfnUjpMNjl/KFybYTlyIzlkzD/vJKITLDEC2kj1ZEy2WNjTrb+n2SSuFawHB26s
Fr9ayCnrkl0wvUzDmVHOXtEx+Pn9kUfLj0LFB3T2sLTp3Ia8C43hYSNRdEe3A5f+UzY73riEY0Vo
21LuSVvUB8bUfs3hZ8hkzr4PHWZh23GEnpinoXPWkAOlg/B0mJJmM1eqAL21vPifQ4aK94LXTztb
TtpKu41vNu7ahv2PvLuf4Hpxk2c3DXOfk5bV4oS+EyrLsFJdawizbdqZjCxcEZPxtgoWzEGAFLrv
3w5traQ7nt3t4vGsIXtDdew4e4yXiU2j8HRAzmLCG/jNA1FFbitio0ahSdpj16QC+oqcaLPXcDZe
x6WSS9ryYt820aapRQB+z95TlislH1yshNer7/G8YfgmbeTbqodF7pCwW/qoIDiTDwSSfdu5jxY3
Qw71mssDXbSxRdrhRNk+eWO5cF4lX76GH35T9uiIt068riKXMLwMcuceSWrjPbsjn6LRnSpvKpby
T8DSNSgfGzEazPPI3Xfrg7LlKvXaekF+i2M+KqqDmVhq85d5/1LI+dsjp4sM9VFUe9ne7kQvW5+i
Jlbyv0TwNVGPMXIQWKd1Hfn43lxI57pu4tjUNjcYfs0l4ZCKB082jDvpUPbsI47uedL25lqQCEni
Hh1bTyTwEkbPrit+/0pufPkDu2J4AG3tw4RCUEz5Yk7nHiLcgwyjsscb79qJEehvLEObm/lstWEa
63YZw1Gy/XouDY/xs4Zx3T4NFM0bryjtHoMdAiaLodBX+65qJMv4/rZoIoi8o1RLfahKDrU00zAz
DoCP5RC8Gdkttrj5XkezX0bZ7f7Ues7fiujjc262aTBW9uychTMyvUlxtjc70akgGToSiNh+oaFF
F1DwuAKzTci84LDshVH9N/CNRlIDzea6DRPCEFyXU6dmeZeKxSrkLUVbdHfRjWP9dAAdM3WWP7bE
LxDrl1q6mbFg3642Wgjr3bYZ2YEwYppHfXvKfaLhRFatCv2DIS5htZHR8ltXmi4u7sI66dGFJvvA
C1yyBahzEpf28hVmDvXeXVdHqi1zBtl4xDHb547Szl/z+kJxBKyTi8KfWwp9jz8b5a7gtm9S2n8f
/Fp2lmhb2PxSmDawRLvkMy0EC5DtXlgoVk7h6MS0qBafmIvdXM8J+8XgvDkbVZ8JXh0mbyDrqqRw
1giiw7ZGPWMOB3lzXiqgUp9eBrIyVsxHa7+eRIHkNwJX2FEIW0KNtRGtayHRcbThMl/FV0Y10Hns
8S+xzvA6wAKkuqLnEnDOwjWURl3wPPWiQBr2kkBqjvxyMFNsM+vyQNbwtiNxSiFQQDbq4fd2val7
Coc4i3sXflGESMe10xVXqqEipiNEd7IsdhXW6889XnQLmocgAo2kdJk5ApX7dT8yh7UtUMj1oUIs
bFb5D6eDMDshw+tsZkaX9i5UOV6+LSz8cWFttSMhx/7Yr504aAbxoKTUko3yccO12yjzIREM2BQC
y2fg+pb+or3q4r4NQZvEdq/jAJG1vkVD8T8ohntPADNZmshyNEIVCyLrkLDyS3KqeHW7awDF0BcO
S37RM0W2mjvtR5hQ+zGfRh86m3G8iJZBQCFznkoDPy/HfDEtCH/3iI52m0fQlo/jAWYciglA5g2x
A6xIDAurcBR6HTfduNAIddqGKwdeI0m0ujiOFUR0GxM8DPltduFW0mxEedrvS+gk/N/OQ8ArBJId
legL3otv73/F0RMPoONwlTvVxp6fqaOVhQg4oV6nlFHias8FfzW9uIRU67SvDkPGHQivd87plw5r
u4RJrdnDPbxeAdz6pLF5/kn85pqIPxKfTtx5G5N/bNnT6XAM0HcSg8z0kl65hb7WqQvg7olOW5b4
+MBmV9yZX8V1GBnm0f+JQ16ThQc9LLukBsBJXoDn73tuQn0f2o2qYueIgYzrEI1YYoNwf9D5o/PZ
m7rcVr78NZqjqarFx1vO/1JP+3DzCTLqgRJO2FU+2mtNkcfDmcN39ckSqGb6P+VwGayWK/DHbrnC
HOIo5loGpM4bx/EfrbEZj90bwSZtNJ28NAqVNT/57RL9+KHo6OPLVs12mMFf8kkNXe/uGln3TNA8
Q+goFUIfqf1N4la2X6ht2pDPL9dLgcCcFQqBR5m9+I1tfTvrGALeZPkK3ioS2WH9+sL32cK/R51Z
ccf7wkJufSPegYGqqzObp4sG8TL6eW3U7Xw1hoviUbrYbGl2Mk/La8Qq03Q5g1T8tKEdDXDg0wWA
sn9inmntFEQrXfmikOO3peA4Q23xs+DlY03yjxJrkBVOEc522d3QZRymVGtzV2yInFjg9Q4J390P
DdIBxaju8tv0I4JHcYFKCCv0ywfDAx4FDgTN/DS8nA3Q1JHuJWiJ0xOiam23LagcR6/rSbews6pw
FDpZBUmqJMiEJPpIYDbzjUCflsJyNvtOWmBFLd6XsXgxEjdiqa0YIqPEQGypecDTqnr9tqq0sPc9
scDQHWMYfc/YNSebwKea3zbBxWx5EI0Hl5qGSvRdqlohv5LCZh38sBOe8YzvL3HMv5Absf6scw6y
zgEANq1Wl4Xl+Qc+D9OmIVyyvbyveely00hnjQpEXzuDuNaJTsrYLMHYQjAZeE6nGk47PxHU57xA
g0Cbh0Ihi1Gu0Rt4JKiVK8UNhOhg+uoDArZHg5qYhwZSVHwn3tip7IBxuy7QK7xWxZddMZNbJdU9
9JDDo0ZOHsIB1rJdsO9DlG5s8pbsGBwErbogzN5DcPxa6xspzM7jmjW4dpb1uSlCPNg7//Bj2QYp
casbIuaCK4hT6oboXlftxKbHsgsAedtWjugkjkGl2oWIS1m3h8nDZbj98R1GD/2ggzXi22gfFRU+
TVmLGNkm/JIOvYA2x0QkpZSlffYHHdqQJfeNYFLC1ufIWykCx9K0jkYHdTvABZ22GT2zzM0z8g33
oieLgdouI4sKuTHOKQhP32Ym/Nyr5XeKc0W41y2WCHrbPjvvrR8YoLBqaiZ+5KpcXOtp+ZB39oBC
EF0SHOCIiw7ctQqEcXbBr6Bv6SOpcLuVLWJc9S0su2B/rJKEvdDoqWDO7cem4e9HmWGxlv8KDp+B
sD92UFUZIzVmcKoHY/g++LyJdd+y37XSShUEepZzJVfYcW+2YxILD2spQ0iQqUXpE1jYz/y7aP5r
Jne6sGgtf/s/lbNygYMghvQ5iAM49zPJ9gFx9JF2WXXRBm9fDKmdxKTt/6Kn4DtmSs0J+W3nVJvc
ieG8xpN3GbIp9KwH/FJq2d+THbz7vpPj9ccGQb/QUgCJF6L+sbYPrNPMhbmplFjQIYS3C8NCB3HF
3RmbBORFXaCpzxjb2DedBfjJ6DDVL8onb7J6uczPXOGvSn9lgwYcHj+e91PFW4tPWOShSfAbXj4N
pf3PuojhxJdwAHKHKUBb7LJMx/W+rOzDvBBZLEvxZNJPIe59fGPbLv0b2rpeIGmbgxr72mBqT9Hw
Ope/yLElXb3lNssQwvolEGVFQ/9rcCGWhwavEZYsHj4U2A0Y5E5gM2Ghvb5hGwIaLhbqMvbLclgq
Lp5KUdp9Tb414neOLdCbW7cbr7Zb7NyYM2tn7bRlA9TMvhM5mLyPiRuoCjPJm9Irl80Ld8PcPKSP
6JB+6gL+ZIu31rfhwVj9AjoJpUdVK/g/s6IluBvCQusw0U07QmrX2ClPYR/iSe+brtXOOEzTTKqv
YGzoNbt+ThAO4qHcZS7H8GT6bs1y8JiifZED0WXQzUJU0/A8eU5/YSwfjyxqq+G5YTJ7KxrEGwjT
9YiweQVERwf3EOhAHSrAB8jBMf6jR5JruKdcGO0nbgoVkGG4wSSYhBLgIkqrtw3F9xcrWba3Ab3C
klrVxygjuIpKoiSxCaMalWB1ax6Wr2zLT91XQ5U9Hq4ZuWgTuQJqCSr+iJhNyPBzQzvJdwrucj2P
NTpZL6Xzd5NVFDjqusZC8BEvFto3dZCttxdMD61X7Gm4UkL3ZsTJp+ZXrAycIaIUFe/QxurJpdp7
KIQl2fRKb6TJ6fuRnlh7rwtpWS985tMbzSoXcwRkQcIkEkhDU/hZug0gTYDXitUX5q0xg5q6bBpF
AINWXUnTFW5zs98AEk7zcuJvkpkn4xd9dmTK0QwFIPV7i4kEA5INVX245q/y3l+CpgCnMbcdwEtq
x3ZZp2y+wGvClDzNOkee7dHFnUOnX2ho/4i7G9c3lwPonSIIYdkBOWyozUvv2IgpFQ4hXkA+kqtf
vaLJR3d8aWLWvqTIpWZjTxw/p0DUchLli1a2HgwIH7xb4Rm9PAhKFpmqU0DmzGvwt5AlKdNOXopt
Zd8EJtlG/euj3Ee/AkmqL+/UFuvYnRx4mFzqcYIZ4bopcDvlcMHX3BmjiJu9LWLwx5VwoA/SO96m
JL+t4CvVNGJO+zQS/qvIqOfM+mnZwipnyUsSbDxuRJdGsmOhiVgRa9p9h9qWjysJIp270jO0zCBn
bAlzayxjooHVG1YPitUrYtKnP11GvvLQ6Vqd2K1dgAmMRgnU7/ROyVscWv+DmlhVJFqv3fbN5KTM
dBjPI104ZIeAvGTTjBsL1DLLhKgticjUNBq5bPoHJLIJXs2n3gStjnHNyQe0VnYaQO+n5vxrkwQC
xj8aY3s9dSNy4ojsl/4cpCNhvXZWBiCMDqHvLxnUL03HSSD8SAspy8sq0gqX0KfrhUPy30Ovmpt7
Q2yzJ6wGFMU68/+bTMo8tJHkqdgrNAo6G8XxXRa7SjDLnUJbgdWvzzXijXEjgVYgXJtdrwB9UK81
ZgzTWRjWu6CNQ4eG15WDUEe6vf5XjC2uwn+mWkBe5+u2snhp4xxYiBIhvgJpPRPjIDgv6aDxHwPH
iWrAOM3dVNNh7hXuzUWkbnhhKo0je1/FuZ/G4jtOViSoWFyvsUkRRhTCuyDd3D3A4dTw+vfzzKDz
Udas4njq8J6aSNifRVKE5ALTDHTGSJSRjH0nZ6i39rZ28zdqmPm15VHl3vbWDayzgRyece6ySRIH
qhOxN3+1Oqkat20MVuSvT8eGgQ+cL27UTyMAKXqYHZogPOTpr6rnl5ffNp8AQfkloQGYK9tR2bzj
Hb53Plu2Ixq2UCATSiiMwSKWx9s3gEFFjpML3i58sFyyHVb0p2SV73fB9v0o2D4CzdZUx7pvGmrf
/YgFb3y+QYazgdDzbgy4iWBdfWHR3F0Mi2qJaV6b66SYCey1qubL4x15KZSDRQYCJZa4ug0NjvFt
BpxWtVcaTgT2HMWn0RwnoCaeeYk0G9wPEa0k1FbrxcYVMBTFNwxVZHzatgBek49o8l2kX8971LKO
B/4l8uXbB0llL9mgnFQHFt+KDjogRVaZ7nxZ5YB+IjFk1EJINzC3P7Tw0Sfryw7TAirvOCTwI588
wlXybXpFGMYwD6D/Cs/IF8iCeh3sjv5JwRjldBLgbdZHBKHKNnRtih7BFvu/JcX5epr/MhDM/wU8
XNxH6xiXBz7MAhvq+QDSdperiN1cD3+ipQ7MCLzPp0RNNZNdEWPJR7Y3X/TznY3a0k2VreMWxEOz
s9mnJJ7rCgWhUXlrFqt79Pj+M0hpFiiKiIFKWMhxq8fWz06Xp6Fb4c6CKl9pG5wvHxgS50/xAgXi
xmPMpHtz5xHEIIy53zRcnpjF6xRWRpOswzclvW3S76TrdPeHLIkLHbUlX/jBjOsk3iFlit9RS5fV
ei97L6ESF4t6fM5CU7Zax8Zh/YSTm/SL7sjscVKarqgN7CEGBVBS+fKrb+m8tedGhEaRgmIJ1YEE
1ygoT/tqPUtZRCrmZgwhg+O8n6XqyYZMZ9rs8JkQW207J99SjOL60gb2Ap4ID49638m/NYK2m0ts
umy67SB45ybb0CqEEExJyZS3mV6WbITLXSUUG8CfvcwXddkfym8UXOHg5btcV4YTWSLjeGhbIbCb
O8qvNk63PwOg6gjKbcnNInrKiCPhZnY3+iq07Zt+3MDMRxUDLfE6NKMHpi/pD4HDI3DKFlyVl2GE
zVOUGUCoaOkYicDJhMtGqfHGwFq7XbY/BeuWKnpyy/9np7bY2zuG1GNTqdzGskb1qeTaDySQGmw4
+xnbOlUrORx4ZnpCOdeHXQu90lZqCbbeVKV6hAHio7rFZWhxk/6hY3olONCBquWKGcZlJqGUzL1F
Vh0EF5/nx9usNv93bQ2CWizB+0oP40k7SzW1tmrbDYZgBX5tAh8iVC2cSsc6PVvALoaMyfm2t4t1
1/c5gZZPbnZfTV8VdNa9cZFw2elUJ8e9638Qv8E6HhvvuI+4sb86/I8g3llNqKHb1nYTjnpS3Z3Q
FD/0HUEpaequ2sKEiiaHbgw2vjNHQDX+GdvAExrOBXMUwxFN5SfKnVB6yicB13Rzh5fS+2Ug5LOW
mvQiF0jGNvDVKTAca/6IhCkcDUJ9nGQK1Ly8uwqIckezv/x0t1XNNWUwbR22HhYEw41GhhkNTwnX
lhI1vvXWxM6t+wuqMRqqjNLwNWUnd/Ypos0e6nrALN6l85kDfJKKiFv0D212/66iOBad02P3sR8h
k0sk0Fi9GaYVNuQ42SumB98EtP56+KEErW3dVd4SXSiOHI26fKTPyXPZsYy8DYzEFMq35+/4nyoE
XQPvDoGgmY4J+ohvzMrffgoixmBG+ti5kBZsKdbIp6thzGY9BPv0pybAfq/gLtCjIn81MY2RdSBH
ohP5hIvOJZjQ2D3ZCd0ad10IC6gW/4kloXpVWMzzOpFG2ZNne8BcCEu19r1GvjGj09QLbgWC22la
eRxHJgHQ1tbUg3aYJUK+xRSh2ZxyHOvQcngqVZ1rsOmC1nHhj3YrGQ157GAH1mwTrgeFp4IGxRre
9yJVnT96F/pg8MVQRp8TUpjDmkPJDfghGzmVqgPGq48B2oqoHUfUe8O0Abyr/F99dxUGQa4jGrpP
yY8vQfviUsj9yySawJ/NjM5X4Dx7h7lbecxtvNwAnagS96gumzyptegTFr9v42LtNrO1olpR/vWY
Ay1DAsFBUs8sb53NtX4P0IeW+msA9FSYviHft6OrpOFirCqA2AkLXreg7mLYlRTfTwhjjv7LVWzV
+iBueGhHcVPJVwrlbuxtYabLWh+pFyGSitEPsIns+IfQer7To5E8XqFfUpkN+5uotxsVm2rCvfW3
d3icSAZlu5GP5XII7p6GCxeVL3MAXFJax1nD0IfkG9UBUJIbpbMJLv0tTxXxGAyysNXCsjeacL2b
p+vDdngTV8O1ct2eKL9Bq2uXCLBfGPD80j69pbcTQOoGOJZ5u8YdC5QM7lIFu6wci7TL6hnjykzR
pndsu0oaRP66uTlRp7lWW7UdCo/HboZn7c11FhWtZQzIa97CPD+/wuzLtZEo70jNtL/iPmSo2fWM
Lm6NVjyEAfzFH+t8cq8x2kv3DUKthPXYJfqoYRZTBaNoTQoIgDbtnR1cfrn/O9GLgNZTFZS4mSjY
/8uXgymErgJu9AQ6hFLQnCPY4IL/nH8Tp7Ahpt9/g6wdcQFa4Jm0LBJGODB+mR/5gSnbFMoEjMbp
SrQCe63dAJXeivJO82U1ZJEzZgKEdW3llDdNKI+2XOwjUo3pNT/DL8p3aBjpYtdPYyDNc3oLOiFK
OxJvLTPUH8750cvoy+SX9OdyTpeAza+NV0nsAoZoCTgbvKNjBT4hNMiCD/gY16iXj5kuk/8RaNoP
S6hEWUiejxcy1KyYTP85kz8kj5B+CS0cR9IA8TBAq/T5iw8Uzhgp6iYW9IZVdE8STsVmQx5fxkQw
YPvXuKpLPRC6WbB4S4mXLPQAba0vCG3IG7l3nmmnGCmMm78V7fwvf+LqhLp1sgmtADqeYqT+ZmMd
hMrsUR19DGnWapKB9G4ucGUBVC2TAdJ1E1wt6AsMBObWXl8SzzGB9soDAzNfJwSf4SGN9HXC2Q0E
Ku5pKMmJ+2GBW/5tLxSg8F30Fve9yNFJfiz/njrz+9b68eapAOSpFOd7mCihCJXhDBZ2HQjhBEIp
D6I1zzvzYYU7N4z7uZuonZ1arPIJSsOREI7nwbjL/ZTq+K5BBfHvhiDSV3TlpkRUg1KnipYNIaCV
k44r4BScBnJRZtNXuNLCYE6ohHpN6SJEJNpi9DTFkQFXg/4VoeHKJ167+kshQS29Dym1FVaZGFdG
tkkzjpqGdhQLCbB2ky1bZhqQZCuTTRdbNEiqn1i+0ML6+nIvJfJGsELsEPpVlV8ANNAOM7z03dgU
0ThlYBz+gVK4R+6mleJaO3OzR8w00x/ocGY5pXOPsCtfsdPzF/d6oveDGVjjj2f/SBjL6NPcdnVj
ZewI3HBIHFYtwwdie8q8If1yAPenDHuxfNJXZpulHI7HnrdRS7mBLq+Ycpro0QzsIcRtMxuPS0pv
sPbT7hiulJisg2Cu52NcSXdQXusLZv7pdPl7LlImW217+oQUJJlmEwTR2js8bYifDvd+0sKDn0Nn
awbz1QqXaPkkzRak/Zx+RUNiZ+OFMaE+iTr4TpKvIAnVYkdPAqmb5SJSZS4Cj5AkdvD7Ytbgne0E
yoFzbL5wAvy/tlL7DfeIfrtTwbJMtIUTb97EuYxXgIWM7CtK0buNkK3CDDmHuldjLaOeekWYOeOj
Eq3vmUytomvo+D4ZrYE7X9Afe38Fwts2gYvydFB1Plf1qo+gPCtKZ/I29f0DYEPP74B0YbgVejKo
z91vhe55TGWtdk4FdifU4chtgommeJvhhTyZCs9xAZk0/q7m1Ti56dB2t9Id5HS8jXv6BCrk4mSs
9Z8ZkLAyVG0kvEyVpmGNkGVZ1rDYQee5nfXLObWyr2fSUqy/O6TGfI57h87U4Pb5RqSdUTH0KkKP
cSd1UbyCn0PrMpu8uSBV2K2z0eAOTGobwl5InxGn9qOabV7Yj4PB/T2FEHbzelN1Zx4FBlprMwZL
ERNuLTlTBguyv8+VLY/QmcCQm4prmR/6cE93wkFgTl432gFkssdI7UMaMpUdq6U62NKBN+MGeWsV
TZgTooE5aHypgr4OER6EIaoug0JluONQQnzXVsHyCVRRIwDWiX6YhqINaf5V9tz2ob3ZB4Pdjtly
Dmwtyyj2Vg74Flx4Wgz7s9gb/0FainnPdGTTiaom8iZ4/oNmY/4HssG3sbVkEWj/0vY+gNoImo59
kYXv+Wj5oWtb+3CamvOPNCfyneQebXA37oi/5UXOJpY8pKb2gt1Sg6+8T+nJudbwqoVmvwYQhUo5
n9YqIqnYuZ3riyc1jvkYnq5gpxBGxTLf3/YuPNegaEAUOgDu+yP1bRYDPsvRlxe7nTxaFh+coLkW
x93tR3h9eobKFeJO+13jWwXtnxOaJcAwpp1N9Bdeg79wOPJoBrJUyHgOzmhAwg89UWIyR5gY7kh6
uIOfri5DcH6benxgc1J2s+vOzjdOxisXxoflNYR+5Gv+h5MQezZ+Oq0S2DWg7RIzbxPUH6ITDfBR
9aW6ON/KPJqBKrdWqhX10f0c1DU5u5SrmU8xd8R5nDci2GE1582x+uJ5wGp+pG9OsvliSnoJHzTE
83rUaGQzas/qplVC66/wkr+ZxxOkQ2tL9A59GXlAow2CcYo/2iELJw1xiMcRcdr+0Jv/1rIF4ZVQ
O4AqDH0MAPNH4jAzdj4R6ljSHz6/pA/rqoHhthpQI4+/2SaaWmeKHmafpJwbaiLyLGkamlNdSQHs
nPDw6zPNx9sa0JIX4QcwGsAEbozmVMfx/lKcRkNx/A/vR0Qqxv7wdohUO9vL4TNf/BlGt7bvDy7a
tXylxy0MVVVpCbgwq9rqP7pODH61Q46jWqe1XMkq648tlpKhsTeOwsAOgBswQ7gBeXtWQoCsZau2
4l914mdYUDlpuDqp+Of8Qzo/LtW6gxbW7beMn9NuSCoIn0ss1wF/ZZZCdU43qpzc06C9S0GDIj7z
9QaLyTz7bGH922DuCGlM6vIDrYgOMM2p/m4yVOachJjajEJvagCBTeMOZ39FNQh2PSa/AMdOnpkE
sni0CMQZtI5CG9vJK92W44AdCISc4MmpOJaX1FVI1Y2rr1bEzqSSsq49n05EGIeb4yPZxYyrCG+5
NSjo8b1bOP+3mPqhbaxFG20KA5D9TaavfbEvvgpJlBsjbRYkTHynEcij2WejzY3eLKS9Qi8ji5ZE
2gUclHHPAAX+lIMH+p2FkvepfLUKPVRWm2111yJhexefG6xBv/UwDmB1IWxO+pq9/MBWX/5Bu35b
pYIGHz4SH+HcOz0vvYqQeuErsRJNB/RLQHS5Hq1mHFVrbbjj0Nfd08tTwK84CSWKQu4V2FWptPhX
wu8JzKpKGhj3Bxp1AZVKsVG2kHPSWyqgVR5kzGLywUC+zFrWvWlmDzQVBmcNDX56CkXPg9TBawvZ
33L3n2MB4KXom2RlcTAeEUfytRMfJl7XPXT/v67toJi4xki/OHQTBFkPJSwNYKDQsfCS+iEKTxZ8
/1JZkr+heVuSpBOxdGrsrpek8IS5+Wyp/PVE2H1VzMeSEcRULuxR6Gbrj9dRAwpdhdJDIQ5aofKB
Tal0YogHh3omr1mP5LzJwULq1spvN7QhIAVWzVasEJNXMvDBszJsl/tzkFQNLK0gembcW3o8KxY3
bqW2lxcT5AwBMCUxK8xQpe2G0hsCJbxCT2KzxmHgSep1pTHnCAlPDnVSBoV2qWEHUPKG1Z/01reU
cXcfIfTv00N6Ku5wHQQkge5Fyoqx6kFOcHDgY0VOqEBz68vHRu9gwph36UVzulB6JmHsvv7BOe1M
UK7+GHEvB8DrgKk/R6BtKFmwweRabgW8QePcp2dnTExbFShlrQQjm+LzLXKVXqmboHHQO26og7SZ
lmOoGeQKh3qROAtIL6ZLbewaa540MDIu4cYftZ1WKspkgT535QxIBFVrmEY0xxlZOQq/gfDL1lCp
PIN46VRgkfnkaHeg3JgYXDpApDVxH9+/dTAVne0ngnoeI00vJmVNnnUC+Vg1M+/gfs9sKU4AnsZY
T75e2otaJBv7Rt0K/w/9K0qWZfNYhbNQaoZAe7MeSOaWJiDcQbTAKk1ZylcE+y7v7L65BLU6MJ3f
I9RN3JM7rZN/hzpYKkfG5Kkaz2dMm0NncqubMIOmBLoo9Ien/SYjbYz3nj4SEfy1RBjy85nAAJ2s
Cbpz6NGTCsa5818dcARJsh1xzjcXBjRuew5FBjLoWuqBmQ3I8wXiZrhS7W2E4emoxC3yXhjTIdBx
BFSg/YvDr90/fN2Z2mfp8LWtqaowftnn4pS4yxIBfGPtmiQBKol60nynlg3zNkrXbffKtHtugKHF
TatOjEZxHwehID7edCBotYPikQcAvfDupbJ5XrwW0EHTLuId1BrxbKupWmH3VnYlxNN9JkKDdy6N
RYT3A0/2cvLsaKxP/HRvGuEo65qyp3B3fzhS+849f4AJMUPlLToUs/nXGNpK4PpYxTODTufgROeb
sMmlgSgZeIpvScNogTrUHM16mdsIwdxEtDOcbhNpmgrSefXkeVeTjtiYEuY489t9YjKLQb9R8d4V
KWREbFENLaTqD9wM+or1bkQMXOy1FiMQN8VF/mC7g22dlL0DILRBYCMXmSNc5m7V4G4r0M1hrZBn
DqIDzJlxki3XO3UCAJk0nbyjUZU64faVZXVNPXLvaBUrmobVW+lUj09hwuU4HnAvHSlCTeeZnhzm
q+zTEyR4AHmKhGyNa5m3Cae/A0r5kelL1i3gzPNWE4U/eAHbpuKVPgJYF63nrDau0yREf6U9TcUJ
Jlv1BH5F1BGlwJYHkS3H5WK1xIsgfBqbAMTMKCamhLAkZGcBg2k1cgHYGJOK/ZGsJBjvDixofjAO
m6vBOZXew8GfHEurkMIscSj99ngk3TQ2XAM3oxF52P9SxZ4KJob54/deH1gR3YSnj6+1gzp4ZP/m
bHDpPe6fV5sKt3SEcP/I3blrV+aQhaUa0TAXgQe4sRzIYRSqXE2CEj4wi2oeWW2q8rl7f47cQYQ0
+UhOE5ikhLMO87cHODpqBNvv24IkUDzZOH3ouPUlSsTrKnwHXfd6VRDSo5SGrp4cvsUli74ELD7s
vJ3DCzbar2NMzlO3lYkuCYdJVV1VaoSGYra1Lewvs82a0NliNGdYjV8Hmyn3GxhjymrEh273Q+eb
dowpxFWYxqInbQ1zOzOhkmna7l+aZ2h3aRPFpPMGBfJzD4OKYuGeWi8M2KwnMyvFedG/P5BSQkiZ
lkaRDTcj8egZ0gEwvc46QKPJhrMqev+1/Ucmq2YufMGepo/bs7wi4Uvq5OhgOrjwTIch1WCgnz8A
iTP9xQzqdHbtOZiZaSB9+PZXdpyyEn8HGLI+g4FETWGk3gVMg6jzpWxDQSHDfiHkbVMBk+cSSxwF
w1sbaWeQfFeLIvndRMugW/ATirA6WWVZu+UKgJb2eoyQupkLnHFUVURvy7W2FaCgjHCljVz1XHcU
f/P9VEe2pnYHVcxKumUJiGNDmXtcrA8wJTlqjGDhy7lr8cP/ByJUL+Emlaq8WgKgQKDjC4M3+M06
k+d8omThGD1Fuf1tKJ38yMjhgfnMUyfrR96LNoNs+QOumc3Z5DThGRjelE0fneZpWtnD/3Ckf/pm
hNyO1INNri2qyCGVTSeWRL4zdq40e7OLpcsJ1mzAcNoh6zW1G5HUjkq1cGwqYsm69n1zO1K7xgtf
8vM38bZELnJNUbL1Q8pNORs0nbayeo81kTjnCUf8CWmUBRV7BMAzwsAe5N4rHiRaMyOPn7niLTKp
dAk40Mdm64ud+jmc5Ko5A7a/uHyfxyK5ShpygLxXs86X8t1q/o60srxkrc8ou7XSHqSB6D54rRKY
MOI4iVDzeMmopz7qgw2JE2E8TGWUK/mxKLHcO07U/BK4VA8Q9fSQ5l22PmFqBqFpNRddXJRkjhvq
Y4eNy5Tx6OdXDC4ZmvqKPLwBVHZ2txe5EtmnIOowWg4OFYoGLPG6KLaSxN3VVOevz3GNMFFH+bRV
eU1mYYH2odyd+3uKGAGltDsbsVpmjcYJsxvmKQwk6COdCaszGR2nhzzspJInVtMTu1ltZuq/5HpC
ZPZBvH/8GhWvXAQOz4DtHtLzV398q7FrmWoap2zQ5oNfWYgCxIcITjMl2E0pUk+mTtBER0adN8s+
viIwRKIv81jY8k+b7Qr3esbEuO4si8b6e+nZMBXZkjxADQkqMYJpEfO9t3tQ5uHh0IxHQ+vbFf9L
1DmZov7NMsQhr42YYFVm3UhkqaPYQuiAqXYl56JIQNBHfWSwdZJoUHm1r2bahFnLdm322QTkjeQx
BRxXNFE0B+Xkj1V6/A7UOLMrLJZyXKeDiuXrk3BvOCe1KzIEWaShlkIvzU3O8vSt5/hV/80F5JEG
7G6LajWPmWYivLLXULHrb/mfDOlHhWHkmYepos6JaQz9RfUotvhVGaBL4twaUHhuuYBkWuQ5gnQ5
hCRpQtYvul9Yf+5hFjmGDfDW6LI93BwN+B6jkSQVJ5C/i/9/NkK8NvFXhBLghH2jtXM9QZpJbMCD
QiQBfN0JJ+bddjKlvwIlx7gCroS40UjsgKR85TUhAHOrGv4pUpVMutmPpzIJkjyLUGeA0Vj/Kej+
JIZAGvp9XM7dYVDqTv/KqCS+kWfmK94GcJdeCRI/3QfjvDYzZtMtskgHq5h075W9FzRmNI0A404O
s/cnFavrCklT/jRlT0XiCCQKUM/ku/q8xqw7DfqX5Splsfoh5ZPXRLwUVCXAmZMGbbxhQklibPbS
GTaVSmff9dWYiBQt976V7KXopn8jkdBdiOuGFCBuZhpUQGoAyRylIBckQ/qW0BG+tUdbwM7Rzopv
GQQeX7/vn8QS8l8h28mQ8ByTLgx62wz7X/r2FBbM0otHsb6iJFrNlboBVhIlF0NU9fTIhaj6iD4H
CHOciEc1zCpi+OPP61UWkNyGY04R0jPN7S4yU5ZyYNRzsv9NxDBwPKxeNY/aqMvt43NAuuqh7YJT
ObdCkM+QWBIbR2MgAx6TohsbdORxmy0eC+X4pw/AKLEKtV2AQAsELpJMnYX4mybp4jpaFuCUN5PQ
BXvUN3IvSGSQl3p2jz1MFy2IcpdmJ77ccJ64F03H1eMYkIjBzthMpwYypG01xfcjlQBjbKfJS0sP
pxpxmYZtpfm/lbOwfewkypiEbl8xjXg5EM4HN4E2My2xM3qarm92ScEsk53GNwLC5q/dI+3yJlXC
7DCboaKDN9BHoDmlz0WwQ1SDe034RimCz8w2qYeL0uNhTGo8IP8SamY1Qte9D708dSgv4+jabzb1
QO3Ow0r2aPEztkYRQW4tZ55/sNC7dHqD5fYYO454PD/QZT87M4gX8TBkYII9Bp0nVzoi2/8Y3seS
1+HUp1URPUu7a/TPXZG9VQwXypI08ZF9G1mOTnMtEUQ4zNdN6hVciGPmNFPZtGlmiowimguiInfW
9b+VhF1fbBfytij6Plvp28wHjr0nwmowJvomT8FNum2QThboi9Vm/wxTe7ixJds+4qtT+JaKLRLJ
/3Duuy99jz2yWJf6S6kycESOnjLdtLi9g8M1Iiw1EFM8nUJGZlk9DSjQOvoswwJhDogf78kwoULX
tRUutEiUh1MRRE38KISztxbkNQuGxQ0Wq+UsuKFvYRmZnb0EDx4f6FncG9QnvKCt8RwHyIN3RAOJ
us6RQYh8LOZSOJEsbPojsZ/Ok5z6L6MvPGclAiWDFuFu+zMaDC+qpfEIwlcKlnD6dA07biaTT5lR
Y05p/tAapSXZfpzsBUhhEiZzwBIcpSBCpjZ1wH1LgD6Ox6VA9iFq/ZOqTMptT682K88D3NVWXAQ7
S7+13QiuO5Bo0vX2y32gfn4TFY1A7NJFgq2Wr4qEHim+7s0yPfCTTQ7e6J8xUyBQJBqQqJG80/tB
wJ0k/WWmZrqjMDKRQpz4xxyrc0kVZulqs+LyEjWc5H2/bvzzxD8v2/XHsUQBXgADAeRJEZ4sf+Ji
uxv9UfZ50H+Ga+uosBNCileXQgaToGsEi0/VHmZ3/H9w7m93NvZZ5Qe85wf8UApPSLn46zkGLtq1
UEwY5O/EyMjtHsPSVpzhx/IxuU0mJDYXQAnbEi9zE5RceaUt8x8ZXWRfumiitX1V4lGd5gIm9oY5
ppJA2aGId8nnmXKcbKfjf/NQiVlAM63w2D7Dq/Z70n1XuOLLJSxvUTotE//6aLTH0pT0HthQTdVH
tcBZlJGLcFOWZzUQpGw6guIq+ZKfUwTmhVa2kmYKN4ovTXkzu0Sca2A5cxqrNW57bs2u4iiKQNX7
ENYspfJ1VzobumQemWQvXQVvI0m2mrItL1jH7GUpm3VqH2qoYT7Vjl9id7luXDB7Wa5QgoIbd+Gt
xr0Zr0h1+SQ/8vm3WlJDzBCQGLzAJsvVaW+qbbDaOnGwPdwKtRLAKEqwAtWXCebbQfvd6bgwoFOx
9sjGihyQVUSsrs73ZfdI7bLD2FjBjWf7dbXZZy/AnCuwrG20qqdRLfaRYzM+t5vUjcfgk+lRc7Tx
NyBCHKtlVPg3+qUktnyoYFRkxxGb/fbPjhoKTP9Gz++CDAaGL7aj9aAcYj9rqGivtYryAC05oTR5
YqAZXN4PDZ3rO1ovQDPJaV0AXGdwcv8zwNOe8J33JItx2h4FiNB5IQy+H2bKbBg66Y6Fq7dvkBYf
x6+Az1Z7UqT6b8DpCRcmQPjEIXemwe8H/h2Dg5SoCqHjiPo7NzqLINABtrc+rRi+OZyy0rRf3qh+
mJEVHyVOYJhM0gbDBneJhKg+xHakVSXrMWT8ujDKX6tSDbN6m2/n65U7CrkkYwLGEND/GTfDni+d
EIBkXAkPlX1+v6AF5Kw9P9FO/1ggSPS0IpANaShCS1eZRe/PoTJ8JasSk2wGy/0VcS4sfVuuCBrp
3HaTvJbSd77V5Qcc97MIrs15sDBinjNMb6wyTuhl+R4sBwHkOEwoc7/u2JSz/ayXyLJdE+8skmd2
QOoEuBhPfgJ9y44eWrnSuhiJ5FvPbGkwkQwACiKxfVxmEYhVS33KSMVoY2G3zief4dOw657KQeL+
z1kqrguAY4wtmZRWH3dLtYpGipEbYti+crqHRMVzDKmRKA0jg9okQK0tgc95MabgIZwPh7ordDDK
gZZ1E9po4PeepikoQ0SUY6p2/Mvjc7UUjA5qyQ67xrGi+GC4UKFlR4+uyjgeHz18VrlpDwTwtHPW
bnXW44+t8LTDaAvuPJAD2qlVW7QC6OfqVmbyKqcsMhXbAgQg1NHgq6bvSX2jA8+V2y6pSObHppTR
PbfYNOFihkyA5uj75x2gQA/KKtRPBh1g2iLJvzCPOw9BCOBTm9WML7SNaWow1rzrXreCKCeigZrK
bx5Lw1GlDWfnEh0tdnMc3TwBDJfrt1IZdMOogH1Xb4ZBivI2HsCy4tlhC1MXvz/YKvs27QzUpVn9
JhElbmzzh+S3LJ6XBm1ADr/bSTejf8hqYD6pBxcKGAhvWmCdwNH6P9kuYHCH1+xL8rMPxfQhqV2M
076snOqAf2l3u2ExQfjvaxP4KqeJ+W70o2U7y0FSdUI5R9UuxhoHLEr6qucQ2rdFfSiZIDRYvWJF
0J0SuYtPtDoZOUYjDtCjxHGfJsmaDMfEtiK3XXonhNQ8+hfMsyR6jR7/O/Y3SWHYQNEBXkx1/4vX
kPoG/u8LU2++utHCVnQIc35GPJ/61sMXvWiWQViZ3aWvaq9shcEr9/R9KCy1LpuMsq4ZRY2r8a55
dH+uSdUpaKLs3n3R4E19PuwHS52Va7SvvLB0pTcIOFkSU7JNtnVl2I1RY9dhVodJL9j5CbjNc/+5
eUilP623YCAAOjKgTSQ1owkjvR/eV8CxS1/qgAGRPtzqXL8cjFAPp6mUeBvHFeHx1iP4iKJhz9Qe
Kkut0RgR2QusRsRvWn1ldKbrqWllw2nAzl0oRvOjDrI+9rZ5Enh/aEupD7IkNjOtt/DzgcJ2c5Bm
pZMvqmL6cOwktaBzQoQVLwE8Tsiq5Y1z4BqQYvE8222ibjdM9wH9OcgYKpvH+SbqumXGzWnpIIO2
ZJqzKiUgIwWwbTeG9ullM57ZlkumVn5ck3T3pbKLWfLBXJvK3fAv9JY8QOjrCUHQ6VvhJirMaDVl
wRtAEkBB8zmcjH+nBfwMm6MlPLFNZqLeDtn4CDTJX/fy5lxFI05neugSuC7zy2vp12poIr61iq7x
4mamwMX5Lg1pscpQEMHCxDcUg7COqvcFlfvzxjzIuKWJ/s8g9GEtPQbG+P8dj4W0niN9zB+35LVb
tjteypn/6rzKS/5i+cepkQTLBsGkbZYjdwR95acVtBrhFcLYgY+eS2klhb6vKIYSSMxBMFHtTmq0
1Pq5mtfPVp7fGC6FBxXooAsdNmYxQcJXGheFzAZeWCkLhK+f60hzHzP1zDhybiviakFInSqgFKhh
zvWeiu+h3ZZ2ntCBXaVTmRA2G3cWVidvxDCYFadOrBO13g5s/ME90T+qIu+izd5zpnEIo6G28l6A
JHTnTWAmKNvL+4kWhUrGcI/WwXKd7bxrAAa+67L3o9BNfGjTmc6EwseukIWKQJFCMD9+TznKs9R1
4lzgeg3IAZjxHLVYATGx0U15RM5q5Aw0XB0rx/2bnH6gezRz2lC6HwSJkKH+ZtOuGUESyZRBRed3
mo0QQoOApgFLAv9NsofsBkQiQk1MXcX9DdOC8Z/Klxi/Lwjs2oRoY3dyHM7zb9cOk67TSo/oQXiW
rOSEUgqQhDnnNOdNrZEXtOMKOzWxNbQlg+0uwf6Z8wAz6thDUwBOoEUWn4SZFSZoAhzJKvuoMQ3k
e1ADL+0DXhqsTmrtcZ+Wh2J5qQxgrZmLjHPj/lw3BPcWHDl6+rI4WcboZfTvKnTcW8fKo/Wid//7
dac+Mx1tSP81li7OefWXy0E0Eqw0U12JtF3Ito/X51w35PZgToXzNEAiA1+a0Lc2NKd4qiotA8+R
6i4ob2f5wFxDEQZiF/g/Hplv0Mv2s31S5M8idcZTgupFVp8Mjgf6lF0yTfhJ7JoMouvnuGv2aYGk
YFXi+/IihHackQwc4X12AUBY3/bb1nUQDLrcKZ8AmMVemaWaKZRXMnGgUBER3GupbLtmGpVaV1B8
YGDpaUeV0vP0VUExCBv1vPqmcBnhvQHIaIKv4mnr1DkTdLrOs+OzvHF8V4OoXVBJM2ZKyfsP+KzC
X9OUb60ipu1YR2M2YbeJWp1RlaLU5YV4dpoYVeuexZyYLgWAzL77BoeHAjAZis7/ne4Qbp1K+DMo
S5d6rAEJGcLrL3+/+t5w9Pw2Eo4CPpLPg26TFECz6SZosTPQ0wUQYbgHyhxleIRVsdZCs08+sZ/e
tX8xgCD/Pip4lw3tEPmhNW6b78SdlDiHq9ddpOWiX/kZcZ7OdV0hSAD5cIQ6NGV5MVxvgW/W8hE8
SJVQg3YXARUdVCTIqvaMQ3ZVwu1ytW17SsSd7/2eCJPMLTlqIlEefaee973PAuMAPiA5qjl9/xLL
7rdelJXO+7EGoeAySFKzPaWR0Jmv9cbTo4+3reN1h/Qjum3J1w9RdPrZ4AACMVr+4ySrvxGiwokw
vQAlZ3gPFmp2QYWIV/6IDJTCYts3D4qvTlGK155yHp5PFS3PA09lwK/vC7Mh6CG1eFbJYhOWSCtX
anSxU9b7c+BNVMwAaTeInDL6defQ3JSzKkAfH8WeYhe5OAoDrNkeV9sm4+Cj5wvXqrLs/mNxeXhS
4AIbo7d+3864qIrAUhqLHqGlDFsldOfRisKs+V12dPJHGAy7Qlpf0azbQ7pdWO+oQ6Zwg5rsikmB
vZQlCi6/bU1qOSq6jQzz07yc6GQSlXJCbfpzWPp7pYmTNKDaYMCF2mqyH1F/wSH9p3ttlFDqwH+T
uJwm0UbSJ071D3hhkO5L7rXhDuMi2DaCKlP57IS1ulFoRZ+U9d616wbHfq1PggAfCL3C3WOpTEpL
xRuXTLGiQ9FDrs+JVQMLPaiNtfWVelw79q+M4HrXYLyirB7nh1rlmiTsECoRUYqK6CscGxGUyg6z
RmQ57X3FAzFGnPH0yBW7lrXYh0ufMDS96g4yR/SdAnzW2wnODCuZoPQT0ll0w87KwCHcDpiiEI3m
IkdYJ6MpvIKvTaC9qZhhmi3J7paRG0qba188DFfMiysScs7sCz5x5L0xa8ZjOPIzLiJXZEbVQ4qz
iXNAyUL1/Cwkl4CTvBQFHnw3U2M5IUrQbarncwiUHFmgDo/z4pnKrWqb2oM69l1e55CktDUGdAWi
xeZlkmfUX/66iNPfVs1mdD8G+jr1sxcKFTE83q6TZkaCeFIWLrtKfkWqRy9W7Cw5/gttoJNfokd4
Zdl5PruSEFp2t3Jwgs8tHDiYraWFz0Nlw7IDkdYcTt+6KBhNf7Lf+iv8riuzR+JXO0xFMhzeg0Mb
a3jMd1aBI81rPMCBvOSuqetswGW+gazAY0EigzkcpCQGGHTF288NhV4ZsCWDXrhnj1nEwDonsxDQ
z3hP+dkvF6hbpInxzPoX2RqfqlKjANtzu2NuKyMWQ2/1kgT+vN9o/S2Di8TIBnmWlL0t7JumhJPW
AqO+5AZ/dpqu9J62iaMMnMBNWHdqNQInDCFz1CTprZgH/B7PbV9i9J9JxRGlqXb8BPT+I6AR2X3M
o6FRBHsGaM5mvH5a89xEVfBLwqw7tLMhZqgPH+RWnB/faBcYenK+zQNwOjFgir4QmuO4oJEUWlC2
0dk9+z0QRaMLdaehngG/75CD5BJqI4XrSatTCNNgIDEp7a302t8lT4ujEOabsRK9YhuJwZkLEJWS
vnrngp/TY6jGwzSDhChypM3vOJtwp285rfEwMDJZlIXCayfZ0TW6sLdE939FZBtD8Yd1M4epdtyl
j6MrnrxitO2d1U2t6po3vuHYY33/GQBz5DyLFMe8j4vefDDJ0rCC4luWg4Gha50YMfeSZ7lu2pWV
9aPjl39ag0XD1AiWcsqfBP32YI7vugv+8/H7rzh4L0Hfbn6Iqf+Uor3RkU4kg56qGZUuBs6m6cvr
Gw/hjPeNb5jP3kj67kcE24LhQwUMybNguk66iwgc6nvjC7AD0C9CWNpdaVgpAtwsKx46W+IHlKhE
Aj3G7XnN/ssIZHyF0qc3sjsFnfYKDAnZDwycp4C+wCdz2SNFBmaBHhvuAjOVkCiV7AvT3WnRg8dQ
P5gHlQP/wQN1T0ssfYUPIKDRqwcYzlpZV2G3MWZiqtCdT1xXp2ByYeEulFNcrECPjtZjgloxMoSO
jfTJX7xKq+xxTHb69+isXV+w2JGZpY5Lftp/tM2DmBQQf6ajJmCASMJ+nxznP21XqbM7IFAcHYlN
nzlM7Zw6hBDISFbl0R1hsDjYBFQ0d6Sm27mXb7xhweUI1f87xlx3JLPhNZswF4lCIAk6g1U7YYKl
0vwVyKafIMlu/6EcJ8SORpI5Ij+wYySTDJZTU9Gx3BwN63WBsMPvB7TpAOH6mNV1S4OtcllwgJQD
IXaK+sr25qmgAQVmAlGz9C3YwU8JkTD4xLBdy1eFc7ybXngTLNHkTnv3Cpf4yh6P8zZANjTflkbD
5LKic/owqiIk8g7r5LlLz9cLhZK0vnT9jZsi66LlR+VZsfqq/FdYmFJ++bW3MxWP4vpMsc43oRfP
ZM85JM5YYTNd7SVj/Q5pZdobzK9yCXjEyH8Foe4m92AdPJ3NLY7YI6xxXTp5EZum9mwio/fS98gY
zNLVQhNmCs8dRUA0Y+iBIK1HTrUpXncVYLqFZiboPuLh+zWlkzVtEhKGmfnhH7UcqxhBDPZa3+K1
ue2ssBk19l+L5p5emE1pLBec1qqBE5Ijqqgt1oLh+f2eaiJw57LcdqiwH5zSe5eSEpTsL1NiYfyK
/zQEmfBLZj8hiwRJrOgIUuiEqsFYrhE4U+fnLLNmgDINj9EHoyUP+JCYulxhfSRONy/JRe6eL7/8
OnZ/ii5ZLWg8e2OeJvJY2PmIRfdvY3JFPARQ4pkw0a7BG2vTIfTgknGY2Imkiy91NZs44I5HY5lc
jHOBE2EsaTV+SZn/xuyJG9hlFXClTh+JrWzxEwWKdc9pEBm2sYLJ5UY8PzW/565X23Ck3BlXR4Hh
wLzWpntPse2qZfs+OPqzocIYASNRARmitvviTAOqLUYUeXgzHIInBF8BsEBH0+0apd01s00Ahyne
Ta95D9WL/FW2mDbxkNjHvmrPRkbBEzU9CmwfLK1ZKkFzzmF3OiVEykrOyglmbXmxEGu3A1qX8aFU
JtS7HChHYfHnril2D+IekoAhzPXL9cc+Cazxqomn7V05VdHUhA6KlsmaMlBcn75wehYuw7+ZfuFi
2r0x6QuLloSFRRMYUPoaBHE3zkCIxXs33Z8lq3WTTRb2lYmiRTXbcDUr4nMg2o6lkeprfs6ZoWKn
NRc7NIl/2YP2G7ozleXIfT+g7p6JA9//pjskLyJO6b4LrrQK2cRpe1YzG9uPDJXu5fh667TyQTG4
L2cCTI3q7OIBqiud0ncgMX+2cuXBh7Aso9XKtcPwB6G0t7WwYj+BhV1bNrpABPMa0azRyo/vWwlm
Hfn0R5iVzXfTDQJs6FsKju9fqSXhydbmksWg/XdeY4uJzs0BbfvCkiFHs1Nic1JOMI+h+f1+tWJL
9J9VGo9CSFxYQqqlZ67njHzRzt0OBEvVd7IZDYWITi/IJE2KthERktuNxF4Os1s6NUMObNj6WoDD
1grGf6ZS5giavVYQsTNxrYig9LKNg2WQXjvyzO8n53ImbLMCpLmefWNWg6pC6/I8WYbK1dmcVMZh
1rHOF7cl1Q6x0/1lDQxKx5t2Vjjoy9gXKPEruqevXN0f7ErH8zCz37i1FXDCjoL3KelNWSr7O8Pl
brqjnWWfdIqzhdc+3BlhZxzKNVxBf847OhLMv5FabcfTJkePrT0fMcREkHoPlaORnHr8LQq34FyA
EE86P0hGzKroO2aH/fzqrKqxvwZbTkMgusV0t5nL+rBc13aE/w0mx87WQPXpFwszhYgmHO37pRWE
2CdLKJ38dq42HXxTS5NY3jVEfb4xQCtXKjpp5uVl5E9oLRqpci5VvG6llFl+Ld/nqLk1wRO276y3
cHU71tF5vsKFrWOxrB+SAheCSNAERv1Ceuv8k65bB/68wU4PmGlHfvJtqqy4w39nPgMOTjm0eNo5
DQoMp05VTyJeN369OKS4rTV2CUjXmXBG7EOvtfSoPmR23do3PrYDEHRVbPxqCQxip5mQO4ovrAgk
Uyp0XC7I8UkXRdT/dN8DN96GIZcjA1dHx//rPHDw+mbC5e6yPX99RM+Db6NC8p3uyz8ckaqOob9K
PS/HuQYgtP9VICl0VW8ll4tAWwniKWI8PYzxk5wZyXsWuDia3Jo82L4KseX15fg1+P+LvTSDfKr0
jKoyH68CDE+RY6Qjj3ntpE5ffxCI/R559apuA7flEmjPUhxBw/0GfXKTxKMJSwRWIYp5xf6AZxJM
cGJFODRpwq5qkR+nde6y9GApqpYDHhn6n0TIHdGhFyV/tYXDmju5WIhHDZDg+zswTS8B7EnwcBd1
4zLQKOSaMWEJAN+Ud8U/kEN76ohYCPlRuVSTPt9ptRIAwWLe3EaR8ZbWo39MBS6x3nrGeqeS6Mfn
i4tRnxehX+pamC6zCH5R+GZ6wIFN2c4WplUNOWJ5hXzCc4MNtDD6RqNg4UQu+GNGTdTUQlNawrQQ
Qc7w8um9rNaL3jXSIrsU5Tnt01YfnRkuq+ndgBKA/b7PejxegRIW6MsRxeasYibZU0e3OQY4Gz5F
WFyFA8oWG1VTAeUD8l9MBvL9539ZQRoFgd7uUgYnBq8o+1Ee1DKNPe2AK+dXs5Hzp558JrGZnvry
DJf08Nn1Ov5WgOn9fJeF0FizT72Q09F41V62ADdfM50qy7bZdhrJhnNJRsHybzzbWAmG8rn53Y3O
p0LAzMj902VoU/7upRofK5L4HOymjm0JfCKVedxFolDTpl2uIcXfi4FAlyqAQHenPiY4ZnPinOSm
13MrZ+Y6gK+rk7vr9x8uaZDjfjXpQrcx+EHxgC4JuIQVnIeyV8s2GVP0I8BjiSqYlZt3khpVC5LS
Y6EK+UmP0ZuPD6ZO6+TCm7yiwmwt38Z0uMX62+wirC20hCquLRKI390JBArOnq26jV21RnQyJqaM
JFipLc77NJB3ET8NAIT9BYm7BpTyKuunYAhCI8x7V2n/Lhfub37vqb2sSKU3O0dswL1WQk623jmj
LFemgebzw3UFpuT05ppsoyQ6uKA0z0EcgFeUxxTAhFnf1veB87wFDSf9FTkKjEXrH1g+xoN33Aql
iBsR5OAZKGKMHFE81oHyLk0qY3Q+qNq+Bu7niXEYoD/i9mI46LXNCaf8aRgUA3zou9TYMjmVeV4S
aH/+R6rdHjbyuNk0lmTdKc58XZqfoGhJC2FG/Lq8m8M2QOMBhlKBnzCSWMTh3zDbNXAF+qYTaXcq
KvDL4s64fEbDnu3rYFlKblNsknI7V318pt0092p4w/xOEPL2TWUBAMkEXMwmXAAfQaue8PeDFkrr
as9GTUQiJ0BMKD2xTljULkV9+h7Q6EzBXC6O8WUoU6oSjLR3v46sZbCMmAXsUrXsDo2E0yXTxqge
rOyKBb378O+5RtDe2ZgcQ2axWVmWaCDEOz3Fgme+aCyZbU/UhSJrF4ysoUMHrtlopex4RkWVG6Ms
TjJ5vFr92Eah09k9+w5xjgTYy5edw97ebVbpBLKUCzyKS9SJGsOGBaA/qJv42sHkCQta6hq2k60/
ENeVA4sAaVIOEbOvaJ6tPQfjQInxR3T4CI+11vWqcq8Trtsc7SVrGnJdH9V1f36MsgkF2TqZxFe9
7enwik6K5Q9KC0gNKP41uXFJIsnfxn32Hg7cMdeUodFYZjHr6NKGZpiMcwVtOOVJI5CxSiQbggrr
R2qbD4Y/FwXKBSa7GkSvpHtGlhV2o2X/eJl+Z2bszVgjRCSkI9tRNqGEbv1F2gSkXI56Mx/qN1Ma
6NV+rZv7oqpHPgHCCSlXAVzXhK38r+ozNYncA2nqCJR4qS09f0EshEGLxH1zx6Arv5pjU+SkLOwX
KN9g6kSkGuTDRTFVJLwFvkXgG10QIfkls9XvLndYXvEG1P2W4eNPHm8k5azlXY1bmVNZv/JxUkB6
VywHa8/B/qtdCH9xVKFqrloRczPewSLB4//pLm6EV5EB5z1sGeHIGcLg8w7c+iFcAIBX6j+DXqWp
2nsRhaOgkmhTyg3oR8q8uXx7/fqwZE2BuqRAMPebrPWiwTOwbFuuJop6/ki7EadibMfGth8BCKXN
b5ml5DFtblpjYHNDC4rLLxU5sHClE5SilICxH5Xfa7xlPavVI20kaH9bPkpl+qHlyrSBPKNO2hYT
dEXa+ZhlP3L9qGqDSlJndTW4OTdjLn3TgmopDSwzgDjV7M/oUwZ4brkE8ODc0q+9oApqNA0PTOd3
OAXcDtaK+v3yuQfaprfaPbMPJeaEmSpypfFazodxv3I6mE5bPCoXxDaOQ9Xw0KKMt8G71efqt19O
hAq8UlsZ533+Dp/0fAPpmQEIgoN4Lwd+nZYLRdUqBy0wUpLgm2EiMdL+segfeJoEgJ2nbBjmXOdW
2C/Pu+LIJKxMjBfXuJMAzp9YPveAxbtyj5asN3oRBIn/D8W/6Y8BHAbgwJNwUkFbEfb6AfsHnsGC
L4yuNNEfCATLtlUTT0NPkNw03xUAO4gWV/sJms9K9SsGGHnbUQnZzkObH8lNfEBGTuB1T04k5GSJ
lD6MPIOUAbeGdJQUA1VlFLAnbXjc98q8WcKbeAlAQsaZsmkdUOHgi52cuqpZs4rQM8KJZdgrhLvG
Bwb9VXK4LVawX1cYFTnPYx3SRkvpl89lxhrt+D1piSML/8GRMp3hzykh1kXXmxTF+qwhyWxL3Fq6
Xk+kXdXEqJmg/eYfSZvsI28mwsYESesDTyCDTWdzvLgug8YiT8DRtftA6Lk8UvYWaoL0coq2ce1U
J54zLzmXYJfP6k/xBrY4sGbS/ZsbadfiOZDO/81PSVQs47SMow9dRBBe8zb1NwWCt5DCmzj6cmqX
rv4NmYITCreWgpbnSNDiecvNlzwAXBGK4ggUDpx/m3Y313Gmn/Zd6sFvHT/5cS7LKjjHN3dO3IP8
Nld0kPW0Nd7r2tLKoy8Ti05CHDCULsSZIkC4PUo67lWysoIUjzZQLOE1fKFkRRFWy9iz3fYC90Aw
PZHUy32zatH+M2UpKSp73u82xkajgoc+DXcr+uhSyiWdkvfqX1+PUODZLmJLMRAhxRMNC9cvZz5R
4J6Q/gMRxbviQhp7IJSg3kE7ejMBDQq0UiKb9SgvUuR4f63wCmU70v6KKqgAXqBXWJCNmXmftAGQ
R6z0H4F3IyNbm+X0vVXxuTcnyP9/PQpa0kAXOxxjlZRqTjFwf2duHHADWxGuv3BooDgJ9df36zLu
uT5SZ+Q+gmtWDhqvgU9esk3ZFVek6ZyUcEAt1eg3i6RFZWoh7cArGiSx8UbshR4OlEV9+TIXghw2
I2395CZCleGkNqnTuncdT5HtblRLCmV3Fp4w8xfpVS9jul/9jhOmT7X4oDi5sUVe5uwMeS/vI4aa
qcsMAU8td4S3UtvY094s8o9wK4iej2FbKswXjGni4Ma8SfIpBfIswqm/qSbNzeBYQU/42SzvZLrf
/Oqrgd4yl83/ffXcJnpRKjUHz0oBRmKaABWbvzxoCgCeV6xX/8mtPZkQ3wfjWv7a/MpL6saRhpTJ
vMZBySRP4I/ZmI9rgnT1+xGkMjx7tzLTnnSClRPahGx9yt61s51jT+sHOoyesYGcSkvDeYtfRQjY
iA4uMEKYY2TJbiQLwSe7TOZy4AM7i6fr1UbmIFfDPhqwdIPAHvoJ5geCGIau64Vg6C2KHR58hABO
YIhQmUytVSwNfDzzuV3FflEBcREwPaqiUF2r2BhWDR1XQTT2hjFTKluWq4EEyXIwmGA4dhE3e+SV
pW1cqE/4G4ZBoM0+A491ARRi+bRGnwvdZBYOriEYhnxvHvZJSF34CcmRGPMyhz41PDL1+4aUfEc+
tgdPVMV8fn6K8CAXgyQ4UKv/RUEM01zTqV9jQc7wurJ8PI41MN1UO8WtPhesauGFqBKLpL5Th+PB
Scm3QtoqrSdQvZCE438PlasRlXv2G249K7e6T2k+YBAfuJh5VEvZXi23DxqDVPHWqpaEXs4nERUQ
ZfISIpDXYhigloijKxDeMXe9TrroJoGMYcmjq154qnDVcPUzYxjtyFpzpz/l9Xg/uyMIttKI71rc
1ZymY3offY2Bfm68LUOHpai8jvLk+hU8rJE0aZnB7YlfrInPYKMaeDxeK4D6l+UzAVVirEnaCJoY
koPrQpFWRILVY24csWvfX/F8nHanHMEqOL1X6jSjGs80z+AT9TeRDAeUTSvwhiN4nWZE32e4qQCw
1HhjyTj+28ueCx2KUqCqKNMLBRkru6GTuVsaSLiqGVvDRaaBqSempANBhvF+Lg8A15MxYcjTn3ak
06GQkuvBd5lIrJdFxd1DoFQfCPGg0Kw4yxYdq9HasM1RVY7hM373wBXnJgBrKXQWc1ToYVBoaxNd
DmyAZv+6oIQm5T5KySQMRpZQvLSGjJ6e1+E0PVt2EG1+H/MA1z8A4GShKgxHlkUIpuOPuq/niIWO
XR+gBYjPs3T9oW2Z+OZhQXv64tqnYwGfCy/q4Mo0qxt63YsHirB4DtB9MLom17+/kkBPJ2ALWAh2
7KdzejFBN0pUyEiz5pf2eHriIAeTWCevdb0nuSb6u7aPxW1dKFjYCJoI3WUZmBJLHGTodH+kLLdz
zwPY9t/LudO1An9jV325MBkBQCiXn4yvK0SI2xiyZghbvSYfAGDr93uNpHAZpHgB7J9kuW3hR8+i
3K8MJ1BMUN+jrcpFNECIXmnk89xsT/RuTb0WBphJRR1w9wTL4J9tDGkl+COEBZA0vFt8v9oucbZ3
PETFVxgE2PFCGysf/fE7X/7L75+LjV5+dLcSDOj/7WlxHVPWwIaPb8ANy4BHkxXLm5JCa7iRFPLy
ENFF8OWS5pPuvrTl6P4iTTJJlfm/T4e/6bsTLBkovvNF1RR+CWcpQwElVjtCP1IPUJxuMSoG/Nuy
MwpBX6JjqWbVOVUKlL9elI7c7HRToL7wtDHEM524XpPeZckf0BlDim8sPGiWjzsTQFGLC7I8U7Ic
RbgO9s6ssaZwmECGrK5tomCE3wamBR7i2DiFzYMlkMDDozgqJdS3CgXY7bqaCApbYM/M79RjJz+B
QicbbsE/Fmp4jkHpSoFLaGE8gtPN03/FCmGWjWSDqNM+2hZ7P7NaZd/1TnDBWcZZfM5eGsol8ELc
/HaHF0yxR5mr7vxAcGXNVzvzLIUfl1fDfuW1pOw3MeYMYIswvDTUKivNme/Ez4GlCGHVZZxAtLCc
/LS0Gs8N9wEFpMf3ejKWtEda2Wy477MybxOBScdCMc8WVI5I6W8KXyPNr+2HAJJLGYDJkGnfGjRS
ZPBEJkSiEE6WuIRmkSku0UV0Qnev2GWfkDlyWd8miGmI0iQHCDLZg7u8wh+8yBC7WjzZii+M9eZZ
otSggnFfMCRBiGoPVHfXNEqk2SJVduUwSN3iHxIxTKGVZpxkMB1FzHyXMjd/6b5Tf6J9eS6bWL+3
etBWZYXoyRr82iCZoe+GQUXBZKxUYu0e8ykp9kXSCFnmwK4h6r7Gis40ZfCDRuBujrkNcE9gn8Sa
5BHbLBt34WOKylnBoZNIMDtXcFKqSzHqXSj9PrkApooFLMARGMRJnf/KIV3H9ZIc6F4zPrCGyVc2
uK8NpLyVNvOyE9UC73cgaB1+Hd++AhxRMfxrct+7Sc44DggsMgp7lZVj0vCMDpOWRm/kViYgrkmo
kofjz9YzOFyZoznp+/3h+M5Y0JxMnW8L4smr5mthb1UK8g8lpzPEs79Y5hCPjyhVWGXPKzERN9ZP
lABjIlz4FPZ0z/bSL8aoaluT9PoWCCHFU9eB0BVBIwGgZbMxlCgFiA3Zpz5ZakzKwcdtXQKNDk2k
WnlfV4hq3kjSgfeERb+8vju8kWCa1Kjn50GIxGrAylH9oZG35R/2Hpa2H11JI2QoDCzwMOx/wEMG
VN2fKvaRCaOvLAYcvyJkih0xSHn/KdEmPGXVx5j7ecl/Glggm67ZPPEpmsDw0gO13XXhjOVebtRp
/8rraZKA+DgFhYWx19X8uJDS4k2ppYCgd8tUSCvdb38HRzkRNJ9PeaEGJYNJvYAL5ORUmdkqS+Of
2QksXSwJyBrlQD59zf5KNdT4inDDazlx7tGfthF5Z0YMLZu+L1tUmR53TbiPp+IJH6auloem3KJb
ZOrZH4nRNWKndvmDzrYxvo4IDV3Q/igpxXjtHCMXw32ZTuOQJgQ05+MaauXVxK4xWFbrcgYdQ6vk
Hu8/oGZOgc5VaBzw0WRdJy1ttUiXNb+UVRH3fkuJmLwythhVTeHSkjVbKcy8/BefLL6kwKNVV7qY
4ZGcDrfEdvVUhousCuB9hh+K2OsTvzAFKZe5qM0WB709bpzxW9Q7os97nvFrqyjAJhadd8roQruc
+b40s17CUepMqSKJYcuEjSLd0NcWD8UhXlFECJxpQL3HqBybweZZ4O0tXRAeZ+Xo+5vXP3rSJqCk
1WlYU2n54TyTWeBTXBZHUJu4V6zQM1ijtR7la4ChK8yZfB4ZHeLYF1Yh3jCIYQBCmPWSdpaf0sGV
es7djhHw2PMswadk8y8HmGhwRrF90klnaM9DCxUHOMfKBQJfV4Ik4Sj0B2PGrq9Lh0W3p+8PLoh3
Mjo6IClKhBG1xeUiITj+QMHlxgywSWf2zwGw2LgiAYo8kEtT8D/csBpctWFBlCoJb9EZDiUHaZyb
rywrnxBJyfIvWaYUsbB1tf0ax81Irwm4lu4ImdxU4oBRr5bWO9z7n7nFZZMRR50mejZcN8x2vSxx
SHdSeC7+rWOUDV1muLJhzIXka8pZat0ggINm+KibnzEMWvxL2yUQvkouO/3zs40SYTopYiDjh0/5
2xvnDzyeIIJZJDvp19IRP6hMIsJKwgXviUVAFicuwGewrnkhJYNGyOoLZYnv3B77Db/HXFEdDrs6
LWGU3Z+ll8nMPCaNLG1Tqb0dU2IiQXQilU40UEDYFbuh9PN4jHn8N2NJOToPU5GZCpBf/k5iAz+c
HrMO0JvJclbyFY34nZLXPmLrC84VCCQl4b51Y2GFpCGpEUOyEG6H1kthuJnIYYTX9sVftyqmp0KP
QfTJkiiFZpgu/EhapKhAel/g+zRBu75s3ycbFHpnoix4LuvNqUzLmFlQfwrM9sA3i7yKZjZ/nEpS
plauIcjbf9LsEEKCLChqHPqji9uF9MR3SqS8b4ULNYlEjyZ4W/4KCtx4mVgiOZ4de4Nr1oOse61z
skiY5LDICc+UcfTXZNa4ggBvvfp6PC/1W+y3GgjvZw++6LvNYDCYJ0JDUKVLiJkXEvIQ2nzd2V/H
Iq9gBNoTJGYS0NFG+GvkPV1I8mOlxqSrOV2zcVyddz6K/FSC44B8Zjqjb4VofhBFBQDwXeADDMzW
1GhdmKtLGe/Yug0OhiUUU/b8ic1mDJAa2Bsf6NEImQh9F1hiTasgtSXtT9a+bZ7+bgyR1HJMHK24
QQBRFbWa7sLMwx9TS7n2C68WPF9VKz6x3flBmVfghjUECMCWYo4n4EBzFevHShmOxY86J+xDzfxp
EJe5AOn8Ww5totnMZSqJI4j+ltzAEKU26g8SLZdmsmXq/D+G/x6Kl+tUogdYWny0rcIO6kyWeTZt
9Pm0JjBQZX3Z2mxG7oue47+1HoHrHb2kKteivsicdu950ExxJN2budDwGlRF6L+YF/wH8+CWlEnk
D2ev1PhQjK23B0xNS4UGTt3QV3jv9oYtnIYD43I54klf9vGgybyfCq+AFsfLZDgE4XvGCyyWaEVZ
RI2If+yyI626ejI6sk89hBZMVYPxtzSPD2Zl54qruUcFK1rlhhoCplBW4KHgmEvDgE0f+1xpvYNT
U5PtFUTJySiNXBm8MMiCHGNk6MpgiZN3Kac02cfvNNSHofcFJxdxGc6C57mCUFonIGCc6PYeuvM3
bOgWXy5rfJVl1qGWoZWla+N99A1AsGzIGlZq61pPxCaxDx9k6N7AwbgwDD7bHyssaHuSNBq1BQ+g
tuR/s73VstGsmijY0nGfQMdH0mDW3SSD7spYBSiVpg2cL5Bb0eIlqPkcm3D18GwA3DseZfrPKO8j
4xi4dgOARYkpPMR7pDjJbA00L0P93rBEtnJHzx4UTHDCdsng+fv6bDAj1LxaIA9WunmFVHS7y74P
3YX8C5oVPjrUwzwPP+lqrj5zugqEjUaT3Z20k2J/dgXAaGsQ2YFentQuI7sbkOkyu9YrvsHXmuRR
sBkV51fc0CuP+U0O1ZtT1NinoCdWsGqS43IILuM0iyDBbdDe3l7ECSuDif1h/c/6PjLz3oVrN0S9
g90Kbfe3Djmog/RI/k27mGUT95HyiQbD1Cs7E6eqcM6oeavXOasJUY0wkSYHoxAfwXwdPWJhxDQ6
qeItMr/19WBqgwAnZfnSJY+G9U15j5icn7ZCNnDokvL+X3AtEDSIxiVN2yaWQdevr9hettzNvw1a
mZwAdrJ7WMjssfOXz+nPtJzNcnF8oz7f/LqLFBS7uXBFqCU3TnpJX/LdL5d9+9qITq5J14GKalyu
pkPzpCalgNbTC0wxz115/IipLcH9ebC4tnFug3x/Xh2U/o8yPrhGI5Wp4mj5kaTHt3iy1xYsLWzS
LUZV7duabBJZFjQNme9m0gD2AA1ahpJx/+VBdjFe0FB9g7l5hLI6Ey5RYo6W7QMbFqFWMwLBhEps
ATZRgYAwMgoE5skhOmYf/KN4v/E91QwYADEIn5TKoNled7E1c0I65AO0xwz/DxJWIbh85iKv9+Nd
P644h5W2t6rl17adBVT70NuzDmVhKd2DwybbH+grIwI2hBMTiLNDGCkMxtSczEWb3yXr9Od/bCjZ
JiAx9DRHEwlMRqIzblu6tZJ8oknck8Cu72se1nUsaF7yGyX9RVP7k0FHKJ0eo06uD9DLNAjFQ6yu
KEUpwb8BfH0s9R7ZGESyDFZTn8eUAvQSb7PHxonuFRmBXgxEw5KwPny9u2KF9/TS8mnMk2JUE1j1
bbuSuLhRoWMFy7eBZbEUieI34SNeISfjfyuT6vla1rN8O/3cO4GHqrkcIRV3vzGQORQxnTftWgfH
zNuj+ccg4Un/FY4RmZukaYVpXDdf0GggBhXS6NipzyarJXri/mWLDg99mZI7+IoVkcW4XY9naZsi
z4Nrn5we+g0EJnHchAe2UTjjbkN8QWvdc/FL9nC1K0PaLdS2esXbZ6oLQU6rDmgujAQkbNYLtCCh
hnn/wHo3pj0EGKVuIeYEyxZnd/Hudpjq0663edNUpgbVdHoBHS31XyUn9x7+WSpj9jJwkDXqP0eM
jRpQnNp4ykofp4tWqXO+X21d7pdB2tjYitboLdGDiRpVOSPh0Zy2asH+Pg0XHZ/0AaSYq2HKtfDA
xGTgTvUPXEI+jxUXqDwOJCuw32/yxBvgAQZ818hB65GiSprKpGsKAMrWSMnteaFgn0l2DcEhzMCy
LVPo70VG2C6HvqKfKIMwM6xzqWPQsLDlSkgTCclK+35B5UEx/76cgX4jz0GWgW/Zv98CANd8TzN9
bB3Ebqc3C15gxjBUo56yA+roUnLKpX0c2N6d3Ap0a3Vb31tf4tF2NzWtZJH8kJhDfIPiibnQNAlm
zgDp6Oy/lrF/CcqlLk9wB4HT5wsCT3knPJqUqpntJwpxsas8XUOw7adXFzfV0enLrsBtAuFvdbBA
2wZifFQ20v3klf6p2bW8PpJfcbvJcqlQ2GInq1+aeNKqv4aAo23lKBGt9WUVdlRkyVFEBMS5hirR
pXErqQWmniVhc34hW5OoZzFnCTTfv9Po4dpZO/MNz9QWc+wdlsHaAvDlRZJU7clr2Dm5rUBxEwVR
FTOJGFEpl9Ti841qq9vENcg+21y7Nm1CiKdvEK7P7P1O4Qn40qSEYR+C507G5zo0acN7QgpISS1H
3fzc8GSro1CrJ2n+h8qtjcm2rsO7InE12grZWeS7sZJYXiGUdSUranXRtiRDgzvr99M5ViiTKcOD
OFmj4lKRw06b8wDjsQALQ0zE8bn1RY9e5N66gOkeh5X9tUfM4hBJLg188OZvlXHlWJ/yAe+Krr68
m5SPcXsMNm7WM1YeV1YWNwevk2rd1dRmL318hRudZIJgcGJPp2jGqsxB/owoTLi/M1vGXfevq+k9
wv544uoSOfZHRi3gqMamxGvOx37YiE1UUQhpt5WcmwWKRYhhG3FhPHVS3Jvfg9BYG/Ctm4Wn7CDU
CqGtSYtavGXOQfop8Dk1p42XbbtadKExUaNajkZSynaOy7JUNP4KiI3l3aKgYnN2AbBuRzFf3WLY
lLVMYzuADWMd5ktLiAy270rrxlR60B/f8s0ql3SZX+SKfy27nuP470UGuJ5EfHOrb2/W8MUAvm/R
3R7nzDfybzwnc6UpE1SEMiLCZg9q1qRXKMjVbKuFj3otKZZern6ODlzwX9elxoe3CSGGvftzCUfp
OZexzFwTztbf5wf2Pkw0l7/TF5mioMMS3lvncWe6oZlEJOQpzkZ1wfaD7PJHiFa8LScmtnrs+98p
py4NG8MqcrPXBqDFkxnkBEKXqZAGARfVn59BuGva5Fk6dep2HfjmTVBkmZsCFNaZWDfQ4PbMSbET
z9A8QB9lg0dexchU4sCGsTT3h2f+1YMSmGeIp+Fu4QKC0mzBuyJ+N+AOnx9n4fIjKnAfH60Xz+1W
xx6jnxzaUde9S7UFXeK90zf9qB6J9HRfUYAlCnASiYxi9J7HKHatw+xM1p5SkXp6I0lXGIMO+qi+
HkAINOcbFnXNdHxoME9qiLPCLBteN3gFPCD1ZPlWsiNNqfgM2UMFryRHz57DZCxHEsQeibOuNRYN
azY6vWAGXDqpk45Jc4rU8xysi+uOzrASntvVbbKvYTFGaAfmsdXISIJLhuQ4cjDIbhkvwegrCtZ6
uxJrSIa5HCWn5S4VKe91qmvUKgwMYcva22RtQ20wooz0VUdQVrq34m7Ma2ZjEStoxldO2CiekcMQ
ktyk4hucBDcJvIWorwgMoGA6CKHWBe49ktoZUhSByiF0s9kxUokkUvtA2HJZwHFyD2en4Szt6ttb
rANFJgw38dKmJVNmpNHrmAAszUipb6I2A/M/Ll6jFqu4CqcTzWydyN7JEbrk4+J6HsFikuSl6b70
DT3QnPbbf0BGc++tAeq5vPxaVAr7u6BAUoCpi5RRCDndqnmKt48h7HMWGLxKtdPrM3PjMJK8DBqL
R0ZLiI1grx7s8r9g65Mf9VW+9WUJBu+Nl8OxeX2JGC4z3M0iahUkjEIeA7Vv6vKbewukm2GjhIB9
uf2jRUP6gbzAVwp79c/gByl0dtfLxUpwLu2JscscxTrJXHmLQF8cXeuKlKsFRgJxAyX0VkrwmSou
AFIhT3fvsBl8Rq5bqeL79atC6+mUoFlCy+df0/UXRQ/ijh0lVwPtHZs5J9J3QbFUmwZIGAnTuoi4
H/8uLqWQByfbkiINVLoQVkzeLk4qAalop1Ojdv617jjkXq7wDpVB1HqcjxYIoupVqEulPLS2PNhN
ZIXimhGSOK7xUy+y0O7zcynfIHrLFmPJ6Vf3XR7WZrdohKIz9T7iKeUa+VnIwoQlkpRjf2aErF51
O9TTQXVBcI7zbfo1SGdeGKmGtlos49HjvPUyGQKrMtuko7g2W10IoKQH7fDyqHMO2dNDJkVpx8oS
BUFU1f8xKcPjJa5dZG6rEx9DtJbcfswg3ssZ7O0B7Z2apP0St2G2Fi2QcsPGsiEVQz3l0GEEuWwg
wWWYU3r3lNo2cS5JdTtIWguUMUca4qlpTP8zl8Eq6tasSZ/fzOra6VsnMzuX3/nXNEZk4HBvF0gz
Z74XdK8kWYuW7Jnx8oEaEQiCjksMtnWZFsIRwdIqSP6qVajAGNvB7v4CotPsTvu/cV9h5c6paWfx
7kVJ6Q62n5wmbnl9cL/pIm4tjTmUahCX3lkFqFUQUpgqmBN+rKFfw6VWzOPl0rS6SpCKNzqdw4gu
nOUXFV3x43CBnnLC5Dfwup06f2IW3sI5TyA3rpXMmeHQ0cPkgbqhQ8cXIW9PapPQHSybDTOrtDth
UZrVW/oS9W4UxxzZHoxhw+2ekDXyio8WHZAWhjuh6rJfbl83mvifbFBim8bEwpCKlu+0tUdCSina
MecaE+VKT7fq12bWMyHJHUNzkr8H/U5+mDXO/39QkkTWB8Ub3PbnVYZyH92I/opfUfnGTTTMbwxp
UxjzesP9cgewasi4neLQAtcFlFyr9xpWrHjbcOzvIEIRpmyx7uQF53FnpM61sdPOs2ZlbnULpAw+
BomoyM9Zge6BB5SYEEG1Gq8m2y9QCasUXSl0Nl8M6UZt9hmA5EA5pxYE6ulH/DE3QoQwlIfJOji6
soBM+PcqOTo0DIxu22r6aG6VS+w0529qS+xCmJAppZKjFHr8T04fisCcw6NjGSL/GVjX3XoNvmtA
2mW2yK50AXvkvkoikCogvAra1l0IDgaMrBH9sAMWW6xepbXyigHfK9277qYw7kPxeM1le2tK5U7i
Xh+LA87GUy6Reh4C9+hRIm22FK5xcramzf2kfiFoUf2Jn/SlfggNWZOKhfcS3bpP1t39lfEaPTgU
0Fz3JFay6hNvqVFKSuXa6cZFGYMpo9GLJ1CAelNCKTeS0ioFXOGBD80MgJIH3OyvsWxL3dwAaq6v
/2WRiSLosoDlFVBoC8PJmHmf1C1oQfuaPbUZtkcq2mTYbv7pmGL81NhkjUK8tACZepkr3GE4isFq
BFGdWdPTnHhVOCrSXFTiMttaGVdhv0dF61dkb8v8w+i/3NXoM2jeJkvHu8WwiDZlIpV2sYS2u1aQ
eot5fkU0qp54ZmIqTnobwIh0luV776wQYQIKFjU+TkGSUSI40rUGt24TcxejYIlvIYy/4t3aYd1H
NmnDRutGzAzoykJrdqkl0k16PiRDtv5hJLuA4u9bMmS7ZyPDmJ2ya9EayW8WdPqN9ADi+8+5nqAc
OD42G/XriFhgezZVx8vkYx/VvkYVxGSY/yukzwVexBFZr3us6kY6do0/9i+K6zCVnLzBSeVOmXDg
PSHrVNepIZDxh3rEb6Wx53kJ7XLUhhuyLssONm+bXRSemsL6I+enI8u9BJFrPOka5fROPlNBTJWk
Rbcs1OFORekr8Ner6XUc9LRosHx6CXuvbWsIlQ2V3xPgvmvkClMkhoMEs0n4ODx8LqnVd4qW2fx+
57E0plurN3cXOxfz1kJgqZ5vNzJPYBV424gyD0KsxFuG1cFEWdnNCoFOh3bKJ1LQfQKjhEcah/un
0uGwCdO3S6kvGl7IaptLtF0Q50XmLdhKh5dYIhP8aSU9VBnrsseKaUllF0BML6hN5sbggCdje+0W
bP3cK8A4kNcdo86KatnkTbJsaP4i36plw/VLQdcj+uupQoPEnBURtoKcm7s8JkgO0N8uf6D+R6Yi
z9B8Yf7nJWQhcP5KfJMl8y6sWFqIYx3X9VA5XDVkYxX0IFFybSXK2rl4RpWMdZc9VDnMymXdAvgf
tzv56e1HQIH814ZBBBDt/ntsdWSnnStAWL0O7C07aFHE8FQwDeC03mVkVModOc2RPekjSrjheHpM
2UduL17MqtiCMgTmsZq73m2dLf9Pjr1NYk9wy0CaPp3gEezLBUeqwmDKuCgcLN5AeNl+aNMmVOO8
y2pFX/J73lfEI9oyMqsS5p7NtupAp/6XZS1/uDAmBnW/qom3p3Ey+ptKs6mzCy1FwfedZDS+PwWr
fHdJSz8NyKiBOkfwADY09urF1e+S0KJwPjD4k2KuqNXDHTdReQTTDVS6xiYITAst2ZH9LuJ8y00/
8lvWmOylSmSC1U+raaQl0yUHvXgptxgz9AkXrG+rSCcPhbW+3Gwmxt76AMIjNWiymw8/5oSBqBMN
qT7Kf571F60xJZSD4HU7By8QzDe7Xy1kyLA5+nDvNddTePTtD+KHR+CENE71aa5NAG4Hm5oRcEp2
CbpUwzRc/WA+eJzcGJbr6Nh7zRRjJBDRb/e2dvfo4ZUxTdVr2AlPlmUUlfbN3ukEVcZ9ccZlstcR
n6FzuD1f6nRhqQ40TwblvJS9BxewGxPP/bWbNZba7F03yuCLaebOwwSyyLVVAfUAw5LWk7dDrn4i
u0LRyvaMffxSVLdRNqFNMTK4ev+TMzQ8jpakDLnq3iVVxYaNwn1RIpGryOfzo0MJhtW0SQ4A9rvY
Ff+EQI6K8BzwMSRgCqaQ5CN8tUypYShCVTY0NWLnnVx/sJKDgwpo0bZU3kf8OiQWVBnKNWJ9eJNJ
El4dDGJRNxSWH4/BSZRRuJW9BCtZlYXme6CRl+q/3EceUq9jHNIMKaBnA45tkhsRQkPncbCjVJdT
t4/HtXNpjU/AiKyl+Qxux1km8xBjs2S+8U2573A1z1yhfejnZka6HUvWLMv411ByjX3Zf3m/3Mj9
d3BC1cDSyA2Rteq8WghB0p8jwdZEqVaHQDXmFJONUxNyc9tajuxAVtZmazrE3ol+cs13Iu46m73C
MphWgI/juWSZ9mSm+5EyyIn4K2xzFoUE3gvgBjiL/C02yIRS4TdXEa7vlMLJv1n0Vn95c4XUga3L
S63b3qLRDfAUH9V3TN3wDtVuRxZuPRrgcadadUBBphN0HB1TkQ64wJd2K4EqjMeBkR6PH1gz0Dgq
gIvaed12ZfI+A0qIVPmz1803mrOHe8nkiXK48fEy7up0pN3zMWsHJzNHl878wH2GbNNQnstw7ioG
GQBKVbhjgeSKfH4sf0StF7J9nG6s4sv0ld5UerggPLkmkhnl3WNERJPbOUEoAwuyRSBjW3V/uTOT
hgoQDaOOr7+9XsVWNrd/3OoYAHDKp/uEALsWtcq46SJNM+3QUzVJ9isNwpRj9osLGqVitdtoa0A8
e68nfFDTcXjIAj5sBdmjgPn3MYvNn0N7ESMIfAB0M/vT+MVIaq7yiIjRvbW6hx3JwO1tQPu14EAw
G6BdKsAOUnb2E2LwWTS1puu0L1QMNluEAybcvAqRBvbqDM4SwHBiMejRS4yL3pSHG1RBFNLXWArU
/XcPM3HZZNi5DuYlS0sBujIMkXZ5jL0rMOZB6TyfVVnTgi9dP1kCuICJc03pGsUMyS3KRGg7c9yz
1wsSQwyGy0z6VxZUU2ohH7LNHCN0QKs23zqUdg4dDGheoqypCRi8BdJJEzE+cHnINqaioP+oYDEf
jVbGgK/xp5bWUnIJmOrjxRhm5IEzWWIpYPRFqfc74lJ4EdXhOkShfgvEEWJqgcMm+4JYKtsGPHAa
pSFTtXuZfbvaCIJzA5vb1gXnj/E8BHCDzUHMeD5AcR6rOvsaJgk1oVN3euQpRvYBUe0kaIiaytiR
IvDI/DWzF+cm5+DAfTt2TomGRuysEQqin1vIaQBh3wnODvui/xieHlv5rB3begg6Kgy08XbsQENq
U09l8YGqrt/kUjVby8PCb3GRma7sWi/mQO0dzZS7XlKMrJ3cYFtt5AK74dEK+262sy2KivD+Ikea
PnOI4f1eRsuCCtiQo5t2vdPjlg89sETMpbgcK2Qm3lXXJK6YNqYH/E3U1w7QDFeP97OezDBQiro9
sN32iVYmgL5cCmHETfPOEMvKHKo8fe22Zl2jA+V6gZHdOYlxCbZEKgbpjMXrRSZL8GVcbHcS0Nzv
qlF7bl8PrdV2Ejrxum1erAYBSYIz6qy1JY4KH+yZgq8jD10uLfjzzsBoxSeuXH6KNJ/wBv7jpLn+
iauJXKNGHvLUHc4KJZGZmhrhu2qgXv5S3zNuiDGzTOGz7hjgBaLANBYnBNu03KyRRkQ7TqK08uUw
K2hJmemfAVzJSIiN2n/zNOwC2mHAecXHdVI8PHlff1rPIcFLUvmyiw+m2r/Gx2VtdMn+r7VW2b0f
Op8uKVvwwZk4YFjIlDiK39g79F0u0nmixRv4AK6gXM16h0/JlkXsLI00ywiE+DtcSZir7eIozIeC
Mj2zn5bu+yUpHoyVyPPFNdJt4mr+mqrpXffRU0S5JoSHZWkzLLTXC+ZEuoq/V98U6IZaBr1wRzdt
e1s16aVwn2WatlVBS0vmyi5FgNHZZ2YxVLdrstwOqsJnyGNwOokLM+oN9HI6be1r4/oZtHZSdMkb
LEVgpsLqv+xasY05YkpCA/Z0cJX+Hd7mqKHOyDowqWk0mNyjtz4r5swUeDSttLjQuyJqXXlcm95e
qDaoxX0QH84ClPelnFBP/b+M8cTM0hIQmEq7NLgy1b/OjXKUKpSs/+WTS/1ifR/ElxjMPPGtNP56
nn1G6x3r3ULYpMUBtrX/RknLlH8/EzFzFZLbA/P7cEEu1DMh3GzrtoUy/z8AoyNp47L9a1pO+v7o
ljSkEI9/ObsWFEl5OwwsO44PyTK5qv4oUDDXbqjsIQxbSlC6V3BVjqBp0vJl15oRUjLfrXeBidBU
V36+1SY/smdTbZXLAf/eaF+6Kj1qf332BWzVUGN0DfVUtjwN0z4+1sBk6y7kC05SnVedYQ0Xktyj
ZrU8cTWIQlJqAg/htA6S+6ZyxdFoI/0O80POnLFsE9PqzZZFlVZEDuBfuH6b8vCGCdmh/d7oz45u
Da/nVDKY4m5P/eKpAkiD7MQ6iRnyCfKCe7VnCjeSEXe8TyGFW0IxAPpIf/xYVgRhAMffXRjKs7aP
yB8BGk5mAgNwbwdAia4cC64hch0rA1fks+bv3lJ/4Sh07pKe1b9VdD8ujX8qy9D9eyiYwGGEvgWl
Pz2cqPnHtETf4TmSPELg8Rb8wUK5E8XFQd8lucmdpUB2mUOnrHI/bIjFuJFERAJi85kJ0u/ZnGln
Bzum7bnsdsJ+PJGqmUjIYF8VGgUGK8oDtEiSbt4DarAhAz6n5KyQhDtGIurObRlRaeEUcIZApOK1
xcmAIcuQEgOlEkd/GK9GbozstnBfElk50e+dmQ9jf60HGuQxOmh2n/4vtHX70QF+eqzlxYKznR81
5o4FR23pCVZUlFpWwntjhI2ZTFNc3wlEY4C3rAPC4h+FUUXRkl4JY862jv+FZ4epciqKUtKyACRr
cta2NPI0sZlSqqswkdJd4kV6u0K3V8QmY/eTX217ljrRlMsPM60JnELyAvHgwmUhJHFPV8Fqe/Bg
yK0dvFBZVgFxoaJSlk4Jra2N/FY+kBwYUSXQaxZzCf/TcXOMaJaz/ETsxexAxaGN9Fhud8ZxcCvI
ZEHiyGjMugavZ0JxijgDe1zl76mX2M2ziQVYng/LB91g+ewZLBLysGDGvLCgzkRi3R/w5jib7rxs
T/q2GGz/yGjnp7RjKKp/PnwzNBnQnLQvlXa+T8Nnmc7ElaN5/DTD2G/LIT0Bm/+pfzWByV6sjGZK
2+Ol3kONaqNbJsozEbVra8c27EJCJpONnPcu9AbptIAfjHuL1pVyu9UgotUoJ0ImfIg3j/k1U47K
f+AHPMM8VWFtsN5QtWEFtWXE6VrTRRUt5Xz03tsXtCZn2KnAh6KrIaSvd3n4sHZ/ThbchCveLj+h
ZR0Yh9dGmYuCNbi9uwcGUPle/UurKET8lmC037uwja50s60pBr4aV+vQEJC4A51S69T2RaDhHTPC
F/QoZtgh9vwsgGXG3IivoNDuynfkYHIP9sMpAcvVXXu/ma5CXfWCjZlZ6/lAn4vnOX0nHCuscfUC
GAny3IW6Sv8CfYJ5lfcXnxi06Kng+K/h9nrgUux+lGEj5F4x19k04zA/Ur+mKXbO5wpd7LhQdYtg
MLBWd+OYqbEZP1vpswIvm2s0vWtzfCaKYCvLTx/U6tZQbgGVmBSDXkFNY2V+5g2th+Pj2Xq/mOmA
hVQ+g/Fqi7SNLw4XLzqDMFZHUK10C15BKazyBBnCM5/EH+0spYQgVzLk4I6uMBL5Dl8ImTasnir5
Yrw60/PQpZ9zY1qIeQOZPurka2cTlf3tNq7A3yMbFsB63EtDV849Dc7xo1RSoM+SRpXgRzvHkKmY
8+IunprHOCpGRyghaiOc2PuQBdm74dFPIyj0RHwOhge7dX+8UYFlvKR8tWHlhh+9z7Azk/eGcoUj
G2wwOemOyahjuNo8UzSwNdFcrpsOKIcUiFENItTjKTn3j8XS/LNuMWltd5UGUkEz9Hpd+lDJ+0DR
ow+oqTSWf+jPsQwHRxPB5kxYAgdV84/vMPEAtrg4gIRTb5zqCRmmIHLfMI5dc4qijiv/SqBdsq9D
yI67wH7K+/WE1StDkeJMV4E067SHpMmoDcBPoy0z87NhghYcb5zY7B8W+Ud6Og34ly2EEL1IKx1g
HZNDWinkLFPeWq93njBs2ZRP2YFBzfIGpLrL/eIIqtPOzYFPTCpp0oBCgzov9twfh+d98LBYNNm7
9vcjEztcUWerk2niRzGYpQjc8fmX9p0I4KQjoiTrAnim2ShxX8BQrHTlc+NJbUWAXeA24HdEXMHc
GRVPSVB2AIOuIyBVJZSBD+S0D5P2IqDzbMMNfOC7kAjGbziMjfCvomrtP3TazYqaIdrSRmDWXt0t
eWxjXK2fKl4CnSJY5XwgqIlZg9jvU1o4z9VPRkxDK8d/CQcjTpyVL7HozHa/WZc6UmL9O5hJaF/i
AJJyDfSlxhmBANTP6a8yM+zaA+0VKs3xmcdhEu2mhdLs8uQYwWJLL4oFqdP5vIMn2gEyiBZDWa+6
/Xck60DlnPLoRR06e95GIXs6c07PwbDXbEudOsh2lWwyQRhdOP66q5EOFb69RqE+aLQiVapR//tw
v80QHE/fXgoTgiv+SALb7+7nduimjW3yHAkr3Zcp8tIwOqi41SVAbAiRkl0/zx8tlE9hqIYCgwsb
F/98+rJSvQpHhJkVyHWXczp3rNM2u6MXNT1VPZbNXm62gt8TW9N4U/wP8a8S/8z6kcoKtKFjGDQf
U2OOThF/ulLIxZzX0MOK74MP5YckeGf7Gl5d9Y4RlR2d5ObhBRVOi+o04OvHvHUgnDkO1FA4VCJY
Rq1pKKR6YLs+hNX3e+tUWouRoS4F/o4aSlzMn7oUVWKCOBnny0EDz02zd8Rkq47j2f3/sQzV8HRy
7zXBP0PET8NyB1MEgCB2fFhEfBgpZYB3I4r5MDSHIPMLOOtIF+xPEW/uhEMCpXSDOV0qpE7Sr59Y
PubJkFyuCvsaqzBqQRY4enTNM7errOIDhxbw0QZFHvdRwP4+jj2YMrX27ek2Zp/njr7I9HxkpchO
aPtrLP8uCv9nNNJsR+J7u8UzkfXT0e3CF3vgk6JJpP3mt47cQ1tXIdV+ysgbjpy2Jf6KYlsS+syT
+kyISu3BexmGECbRciIOTqOtEwaHFdkGLeDQuWaTjIXlT+rRYgZG9fKjoywz42Fr6xm2bNg4Ljvi
z6Y+Bn1VTo4il3SfHgL/8aCIJNty3xa2JwE7dMzrVGbzWpRvx+Qx2kPSeR8obl0Ff+H5teX5tJ9H
mxdG6uUIm5xsDe3q/ibz5ujBasQ6vaHxR+/+1QSW1kGh7+67lz8KKdUT4tchnlBSAKT9YNjAnffT
KLj3lV81a5WQazQD2AQqzH4GTBJRONMZ6/WzxL6trYPVPD04rH/eYw8ub/rT7/bqsFUEGa3wwJ3A
lus1w0agVXg9FOxHXHf/Ey5rOMSEvXBMlR87yHScs8AXhnpJf08Yn5EfXxRLw3pmNP9SO9wNDJNW
ri5lKm5dk2X8XdHxv8j1Vz5JhTIghZsN4zLuYzOpwuRXGXJqtZy9fghWlb5TYpuiJ49c+5w4FNL5
2jQcJ6NQcEJhbaw4xuSO8hQaR5PV4n22H0tJx6nQUXawialNKMAyO6kAMS8O+2X1dCOwK5kcYV8s
4ULEQ/zdtQkwQ1RgwHiovDxGhStpa6/IXcD0ebpYS9Ol2jooVvdEYJGY/aRFWwV6SNxhjD8JX7Od
UxSFROoYD68gRNi6sBrTI37+cenDArJBxseJqkBt2dy8M40/cr2wW04/OxTQ5JDkWipTfRCcOYQC
NtZTOWh1c6D01I3nyHAMxu8pLX0KDA8vA6xRtlBdk/gepRGQHIUGh3oLOW2i0/H1P2T8O8rWrfzl
VmUdggSFvuzFX5qMJDPRjdvEVUY2l8TdYyM0V/KCxVLOqJH78fyzogu/C+8JMgQCWl5deiFDGJC4
3D7QGaGSrqvkvR0iPLumVLC5A9U6LlnQqKlCP9qYRgWZbMGxLrji4b5wKiTtBdNO31m4fRebKazd
dXPJzTPTPKjeqfl/rI0KaKt13yTbz5Nyv55hgZ5zKFpEJL6SNu4/UeovS0i1a+9zyXPrRSy7aCcw
+d3mRwmiuVqbbjSJlNCG4ONDhM1nfOzfWBg3c9s6nOQ088yUFnH5z7bilO83Y8CibOtnJ9Poy3mK
7kQ9Ky0dI3ZUUKtOfNYI77m24b4Uj6I4V/dXboSLtds76qurbUIf8vfW52xCGsvxxmMsULyGBMAy
vc05sug2LIUW+rQa3RzFcUFGdZ9933GPqVVXL3Nqclen1iotzkaRY+s7DryhrfBUPBTakCG9354u
bISN689Hzm2pCXuG8MD0CHlQdra6Z5Qk/SMVAC7U6YmpF8w1lVPfLISmiA+Q72+G1cjhq8Vk46nw
ob3uxGfzdE8qI6YeA+U25bZUWPe3MS0R9EYPC9xYMT4gaCb8cijlzWQ2ikhHVN2oWt0dWOUkXE0P
IjTL+bENsArOxvOOzMK8zM9apSZ7Dc3lThrUd9SqHohWu+ismV3bSDXgjmnJH0wF52VilQ5knVcC
y7Pd/3yRWqr974/75r9SJAkYH+CTnyQnrsksXQfYjIyiBulCJ91ZQ3f35TYxnznmfiH7z6y9z+4+
14MWm6SNNCMgtqytLhyCO8baMpNazTI4bkA3KeKqc0zcga54lGGuN2rKNkj7h++GWoi7ikSn6l/G
W8CJE7pCD4rBQ+roGDog7LtxMuaXMmFIJVjTl7e/9o32RNBrDN84IxNN+HdPG7g291br2Vh2SAa9
bDxFUViTCwoPvn86q6E0DWmnuJ88zNOaM2W1f+ZCL2nZQUocZw9p0vDP8eoI1d5U/Hx9bpyVyICp
fEIpHRTiLthlGznwXvEr6vwk/baOoln4d+hr/LcE4MbplgoAeDR1+dZj97V7qGRtOrUz4mIulBbK
h37k/wQ5x1H0A9STIDpwsEDhqukoP9/Sr2LlCCNyu22Xw/kMfHXGc0Cor1NC/b9vmORNyQgnbpaa
LRS2HGgScSZeWyAfPBByVdWm0Sa039g1TDE5Y7bvHmfyzbompGyxnsvAKggrl/0jsFroLZFpTvAL
u9DBNDZE4cRmzFRV37zA1et1MOuk7GmwTZJSgMGq0QPzXGpv1I5wvXQUOUm1VdX43DPS74xJ0Tu/
/IK9gfUX4bymMZ9P/RFpfv3cRKqJcWNElnoVlIFs281Ud4Eo87ELtn+/7lal6kelOrAqUMnc26hD
j1dl5QTGLrArR5YrKYtxZe7a7iRY5TG33gAUwRsbTMJwwPozkAf1h4WgnUGdZthRv3dYmyif4co2
eZ6x3uxSnRrxy2NW9NrOXkTslRCMuSbWg5wNFchBVys/kGgMOIDJd3/x2H+gCA94vzg4ypXEqyRd
CatwdIEoSTcMhTda6kDHAGHn+bGFS8uHx+jxG8CKcqwLIapwJ/wlVveH2qM7MoKPu03vN/mLRF23
oCq5YF6BDLu8UEyIcCDFVNj7sIznnO4pkrK+Ox08LnKhUBeNSvgfXE3hTarQeekPNfx8WL10b9Ow
xifjmckSsM+d1o111nu0D8Lj2Q0iY6e7ra8j6lYpa8fiT9EJ7xAvpgOPhQ7wLVx4qsqQXL+JRF+b
TWhperIZK2fzyCIdNTfUccHsMzF8NtiWaPKlUl38nrIPCI98oAIR43k4Cc7v9+7EU5Ww9gmb81//
mBNxsP4b2Tq7m7u2etGXx5xXZidsXiLmTsUVHXkM019YLL/nJq34hOK7swr8cGl1RRNS3y2P+Lwb
vpCrB+hC96MNVQNxs74pymyXjQP/2OcukiqAIW3wV/NjnotMkdKTn5XIYyqsxepFtqgdgTbkEWng
WThFzWAyZGEfQ7MZHKsrzsLEGW2Kdk3cTvvaanQh5B75sRHIaumvYhhYPzOiXZFwCxqIyrPxhto1
DOvPX71sJlLGD/nQrRzD/HK2hO7ufhUI23jk4LVMbNo9fA3kh0shZ9B9FSN7teVFndAJMvuKbjk2
Caex6qeXhUFslfPHu9r9qt+V8yf5wparS8o3sO63l8wX8VPsh3J7jJPl3dZga37P82Tsd8tVV9FN
Hb3FTBze1Ou3rwvEAMTwpME81SqBvmf5gZRoZn6Ipw14FB3+1RDmvGI5SWju09D2y4HfwwdI0EHU
lj8Xcc6hF8C22CclPl3+xYsscTSsJMr15nxHzlB8+h37rkATI9enNryCwXgKLzOFH4zb45MFVtLk
MrabMEruViVjykV2nx+vcBIp5WlJkvDsELsq+4Wp9LOtL5de6+6zMqTEN8x5uRmKmIA1dY0QrN0I
G6OnXkouRLEsQ3c68tM9fNHpqZYFLJUdL7pixtXLZVVlih1+kAmgB8x58OV7HPvpluLyz2c/OsAo
yaCE02wh4CIWTIviSET0e8NoK9fSH9hGV38OWg/gAftM0rWDwmNT4FvrnHCSeg3fMHbQrIaxw+rZ
a7KqBfSAXE46VRJNbL+Kb+IN9hYPk9yjncAOggzUbKSQcxeXVRcVnsET52clJypY8qanRiMshtUy
WuY8II4VyNNBtoN8aHFSdxuxnviQczQJ5iOGW18CCFBiwPpbpux2s36TWhxae2FV3KC3hvdyh8CW
4iM2Ble8eRUFhpPJHHL853zSmgZRdt/kLN9ENDZ/d8MO+HlEq9zM4WrEDmgI4pakakXkOmgcO3Z8
lNb46+7w1vkSUSu0TItM7VRozL+uKHiatfPlNSwcI0gQvdtECVPeTaYigxHH6+8er+1SV3GSFWAT
2P0EnIBGHqEnlq2j4cXg++5SF5SFtYfxqceuQZNvTUQ7e8tMKusuWDofVtKPK5fKst5uGzNymPOt
qYSauBTjN3aZVrowrv/ksNdncUqRdOTGdTyOPqF/+11J+le0zP+0yG82Kkdu6Eif6swGmvQVQU85
86QiDJucCz4uJOZ+714GNe0KkNAkxbo70XoAYWkThF4JPnbJxjKIBDlhWn9evSI/pCYRvNRNFcNF
M2euo3J4fGPC5aTXAAplAzrGfzhlRu++XovIHhHQY9N8DA1Dz6/A4sg2ywFAWvtSzKT4yaANFGRb
eZS8pffVqHOVLBkyAH9SnApGNCEex0+G1ZNkwJ6h/Pwg4n78j1rA/oQX5FURIfU8VOt8syi0Phyo
rRmxU316V+52q69L1qTt4vjcK2BihiRT//hGmj+HzR4pK5JwDadu1FGrj4OYQXmjegDk/05+66uI
AkdrQtcTBtFv20e+IRZmnnw0Do/jmN4UuoGjuZKd/Aei28TewTYWe45oyfhmPCDbmZb68Q1tRMrZ
Ib8Lym4NhgFQISg/52XYw8cYD77RXQpQxSldPJHe9QdJkMTlmiwXn7Urwk62Jl1745DPLmreCI6s
lxl0l0Ycqkb/FG+jaP3p2x0lQhbsZAXdPHgrlKlxWTOuLNtVTZMXo2mQC5JQYaTtsFLU7qYtF4CR
YCB38DQ8dv9PkOmVCQsoFxm1a1hq+tRwN8Ipy+edVOA+rJvEVf+JuLc99cydUdM0p6mQrJSB+wzr
HY4UtoXwedV+ifMntbvOu13YX34tVeU/rDNv2qsX/dszg/W/fFHHxY2bPu6QuaS/6PGjIyr8S8Vo
UzSAZjxMICUwNsBEhOY8Rwee9Wa46WjrjjGWUfYULNEztEVlrN2Ab9f1rMqZLvStj3vLITwWaG2X
XanQm9ESIi0pY88LqVc3Yx4OcAAy93cFB0yGNgWcCTqrnNZuiylj3kgJoD/cm3tqqxV0hM0P5KMc
XIYZisL6gwN4GDoF5qiYOIX6IhKdt2ikOV17jbGKZ3zhJyBYF4V+66dXxippn/YEzgSLNsVD+jze
4hfuRWW6PM7GPoIj4SdvFkI9A2ItbeMt9Q9evFqmFQBWsWYl77JBbDBUM/ngE1eT2vi+b2ZyhMDA
aW0qquNhBE8DGn9sBhuW+WN5wafz1P0zL+/dv8FXxsHX9I9xCsV+3y60f3e4eMhIOpmbDU2G+f8f
mkKnrWuXmvQgtrXeeLdAKdlv+TjUzhw2KhRHIV+JMMX+B73jmzfmkmEHbBoHLmsaGeK88NiB8UtQ
P5DV6IjZqQRX30Ai/rhrwDrT+AhxJp0SE4ZxA7xP/6qsdDD/DUxjxZAuBIqdxLTdfz+Pu46BV9aG
MsYUN2YMkXX06KW2laroKjVlB+mgLD1F4YdT5ZHcKeodA/18DWw6ezaPvL7Q3oPczY9ox9hdQTZQ
yCqxgYIOwkRKnEptfys+GPYXDaH76pokKe0TiqL7DDLXcefqmSTIvNKQ05EjqITJjXfIR7lKe89r
kF68x4841dVSSeyXyfHnbVhQi1+owOE72mPSGP1WCeqnsxqBS/E3bLf7DYneKyBQzf8WWRL3lnXv
OC3jhetSa6hkm53xHM0vvZd91qgCQmk7iPWo1Yk+m191SnHJAXsQM/URvbFHMY+7NzNnJghJeDa4
1LH4ZM55Jq1YCQfjqd73yiwOH9WuJtvHIyxbVveXX9oqt/VnHqF5NHj9ZqIQmQfbkk1mxZGXt25O
w8t3rrvO43hpMG9pyDWNALyR85TTP/RMxdgKWkX3ICsYPtdH70zkNO/3n6pKzCg4wwN88RCUnMu+
aq+qB4v1w7L9V2wbURvT+TtW41LBzMa0C0mycid2X4tz99mL2hgxQppo7Teb9lKKq82kx3FLUDot
99p6MjcdZvlgJtGP3EUTT3ySQTdBLr7hXBClG7dbdcUffVydcuHhHPRmMxgbhkS627BGEKooDaT6
R+TtR07U1rbfIqmucoDqrn3a9usU+BSK5uqjnRzyJnRyj7oPC/+4pI5tUrfiiQG2gsKyUjCYtgZE
2KO26G4MszuGUs2L0MRFzmjESQal7+yBOsCwsuNy8bsXHwoDS94Op65oi9bDi2SwGBiXjkRpt/od
/nKBTwovudDr/2yZUxEnt0jtC/ykX1bdXTm6g9MyE3R6HTLtPY9S4K7dBTc+uyTWWZpVK4gPpxNM
d8H6mL5RyWvvvqjxsPqi5wHTkn0J4OrPmKWOcpmLJeQQdH0b2MYoOsbYCncQlBM/7TJTMh5UkTQw
Hzyfp767oKzETT2JOyTDOqC3qvompx1gP5SJ4mePqJHxgmW7Ixb3Yu+dnCWRY3dZzQPqvn5DUVBC
owmLYxlipkjjpKxwzftpYkMPuoC3ndahSlgjMsDc5AWF7DL3QtEEfaoHuQrwZp5IlWtSp+5iUT0Z
VxtQ2Gt2V6bZ52hYghc1uWOJN24v47gzmQHWCgWS604iVLciVx+x+RMhzWRMhf2T13utBc1XQuNA
1DWPqmdJDuDcqhB2wX6p3SZAAjCIhG23QExDc5sOscFCTv33KnY/+YeHgmDoJtpSpc/b0hSMTTpf
4FFDy6qFaZoGwJdINoOxJhtHDYSZdsHhyzEJw0eeNjG4VW8CfJhVUG+Ai2HWyzMK6+p7DyQvYFW5
6GQIniIUPGR9wbQpnLdM+9A88N0uTRPngyXKyyxFPtWXZz5W8bDOPXPK/04L85sE9WfZrL5fk9dI
TMz7Gz4d3cJvZpsuXtKK0GvnUoRuWhnOKHttZqZ4c7SDbUXFamHmnOznX0EUQ4xEVeQq7NU6RD90
ihK5dW9sIJyjRr/2T/LHjwtz9RaxOmECkha4OzDwg2o3xsIekXf9AdMaQTiLsb1Bs8welu7rK8Mk
0CWZYBx92VQeAzGF9dpBAUVETYfRtszzf/G6WYbWAlpQfFEzoSd0V4AoS1EvAJEzEo0w4Bo1SCI3
6DqI8VSQ78D5Y4Go0sdjIUXkCYK7u9XjzxRCrWNFSuEw4p0xWjm4DQewqQwSvRv0y3vvY/aIzOiX
qYTrec8ZwZi+1O4UggEunNdAuF74duz8VsW5QUCPxVo0ydxzo9PZLNCG0UC8MTSEOLZVmGalg0pp
UUG9FTnVdoxDR7ED55OpNh97QU/s2ajALK+iYT5z8mvpqTTvdIapZkMwM6z5gtiB24HM/jF1eeFm
oZe/kd1iN3vvYAwBuYQNfk4eFuv5RQ6rvYB+r3+vtCFsRYwVZ/Y5q3asO5low2oQmu7Z5nsmRuYU
s2A7VKy1uUY7K3IIil25d4gunuFWxBAqJbHw7oqpx4HwYLrzmmy9Iy8gDLG8FLU1GtofjLoeslG2
d/3u6Zf5LHZ9aBEzWOovTuIQv/OazC1caySauYTJqUl39t4mKyToUQVoR2U39rLuuBgW1qSzM+rW
dMB97keb6Ux69t/0bQLduEEywTuGutu78DZriswC/xO48OUtxrHGBg2+9CY71ZYJDpWNypTvGnTD
wqSTH7CYEWYE3VjefkjxS5QUOwH/BAnc/+D9JzaUVmS0327Xmg/CSaLGMK81kGY2UETTGOLzDyTM
CM13qlyQg2OUsdB6hPu2m/FSqMImP5r/ti3zHchob9xzIi6b2MalrS/3BidyOxp1m9C0Z3ivEd0y
sKgOUmVp3hr5ykivK4f6V00TzURF50rrw77NPPcRDdExlmtd4a8HQuiWmondm7Y1/UwWlyZjH2bR
Uxq6jWQUcbFMPN120x1GDGZcRLz7c9+FdoP7l8baUNiGwJ6pLNFu6qn3OFM0gpjRBK6J4uAeS4Ft
FRwFkCbk5J3wtoZu5IAzOX4STHvDLbcmhVKZSIZNTCgiXL+zFk4N5tnmM560LBF/c6p6EM8DshTM
ji54Mp1nfm/VWmtRWc3DkawGb92dWEhuZsiXKF3slkZ1ymZ+bPVFrq+0/uv+5YiEhi6wPZTf/xG5
39edlLo+B+V4Fjdxa7Ge3taql80aOAPhNGGzn3YHD+Q1M63SZfuHwW0mJEfkp2AnM78TZyySF62L
qd8dvUc+NXTMTkhH73J4scUkdoyJJZiaKKRM/N+Nr+bCtI/DU45x/UfRPGAZvG34hhAUDBgUsX6j
00TOknTfOqPn6ydaSPbk6sLGSDVLkllNocEfgCMt+ctvd20N4L4dr2zpD9ITyvtkFnqf2erH/FX6
hJx0psWwt4YASi0QjrnmuLwy0CYdncpp7F3UQ9iA5PjYcYKHLgEQ3gx1lN/artF9SBnHUX3UT2KH
GlLG2YDIpoBDm6/FvGBePrC42mV0z5kYXollvss3P3rzBLiwXe+cYzQIvKQRGaY19Ina1jz08yoD
xeX+oas4LPJcS4KGp2fGsE0luqWC8x1FiWu6uS78jvlR82yr6fqC/bImIlIwwBjwLkZ7KC3YJ+rk
Sqv3gSxQ/y3jFUTJ//Qgc7OkzVNywLH6TatSsfktuFm2fj3oZEQ7TK6yAFLPE8g43Ki3pRUVHibU
1iyRzKtIUDJstDCaG+I4XIdrHviMhmJpBw3ZnLZvSJdpogYpGgDwLgWJdy62BiZ0S/JQioasQMzL
f4q8yhsMEecTyWgGpxLlQlx7XSUvqH8JeQCLHR2HLnbbQ9ELipv0zjnFn0YAOBMcIY0V6b4bxE5H
ZBtlbI1g7FcIqo0Nv9wg4Dj9BH7pv2rL7VlXNiUVi0jftK+/5poaY/UbMUT8TB1rlo5TcGvNH6N+
EastlrLw/ZpYvekAycZgdER/qw5JJfDoPTKq1kYCfqXUaDkPY0tGPn7rpi0LzQUmBD50TIDuHm4Q
+3XBqsZCQn6KsXvmY1Hm0aRqbvj/3n2xnul8glbXDU7T2lN/wMx66ITcZ88NtZVB410/dcZ3xQCx
aeystpzFODvEPAFkFTCoR+Ac4PK2++SLNtgZe4stNbAhQNIpougxtTcueZUMfPdKhYua/vitOWQh
n/F5hhB24kUURoTUnR60l9ndoHzG28y7Dwq7tOfUe0V6bJ8sCzrtg01eFkX8b9rhmEVbPYoPQXcM
D6xJ0QaUnuz2Glqgb8O2zxuzz9YN15OhmUJPpOEeFWSN+KNeVfpBpZE6QgJzjO6+H/zp6awrtChw
Z9I1cwNpeWbEFQKI1oiauI9qEG0R42gIKCDw3Mr9fPCJrBeQ7ZYiJ/55urV7cn6VE1gi6WAQd40s
JItj2O0m4p3HHIh4TsVK6Pbh3gEUP6lc4n/1tI3/ip4hEwZvfSB0oGrdIfxIf0OrNkgpvKl2tY5T
/w8+wEiVvE+q5l3vpaYaFXM7A8QpnlWTpg8pHrflwxiS1yzmh5MzdGXGecF6m/Arq53YRpJAgI8n
j3WF8F050o4HsIDp/aiqzsjKmJ8VOYx33th2NH2zB/K6GDDRRR+K0/CFIptV4RjB5oeXUzGgeHxG
cvclLZYJxfdelqaGUIAauGTECahyTGyfGFrLOWStoI3bFNDCp+vwpJf+wd8A25vmai5mo942xooA
3gzx3ExqRE/ZbK/ydsR1TIX4Alr2LI70FvnvRhY7WaH1Om+BnIL1YfIyn5bTWxa8XKxVFzLVVulm
u11mI05c0r4yGxpiCFrah4P29ptemWcVd8hk+nIGWZn+6UsS6j31b++5K5yHHwkUdIGh9xAho25D
8c7fX+DQRqRUYUC8LbifzomkLhjGNC1bSx20DpYPf/CnCvBOgAICN/ngRTCnxYQwJWvoA1FlYW3O
I5aBdUOFYK5+CWDLgfpLI6H59OAQxZVwy0Mrk+uuGtUri4v871wtX1WNixeD8LP4t6VLKMRpq0SP
zFWl0ByMXCxd9E4ybPPfFQMUqqUJIjJcP7rSHSF+4Jc22xTUG7wh+xw6pIgFeYNn7XzpXi/ncQ0V
s0TYpvd2X+t5zEiYLCHhsUoBiG97YS8UFXFi963YCwlmDItvrNJ9NLjO8+W3cKFt6d9cSoIWm4sP
RCo6cmk5vnWi1bvCn3U6m3sdyyrQunDdpaasQ9B123p+6mG/eknpwT2TObtnVadTUZc30GRKcUD8
4VypzQbvKH7flaBLEy44mN9ayO3Vi2az2kTpRhKkz3BW2qR9GAUcBHd4t7YM6m2SINyK+Nl8ulJI
sb5E0KQb7MHI5okyfwlDNDRMeHQIjY0qkyJamAMr039mBx+pR/E7BucfqYDG/zHgW+4rC3k14OQP
E9urO/92AgpOfCkGcsuzNYuEIb1qXLeKTddkYtcFC3bz6NOZFqOhqIB/xNuvJqXnestvfGgkZzSM
eFjyzwyuwEM92o6OjbKtetrj3dSIwi2pcZtPmw/PLxOC4eMErf7+9wH04Ex1pKTOBqwZydABARGp
0C1J2oQfFYbGOUGc5ui4sfurwmlqb6xe1oAR5lmZIp11E3jlX2sg6VJZSJpywyWriSrsa4FFfhR5
UHRj13pJDDWzzzErJFZYOA3ckSntffBBitAOt/7/vwmRMRW+dBsia6fNpg6WStrllUf4tMgek0ct
a4Okfhx/bXoiZ435eYcQBiCmvSw2A31YR8eVylroxNKJbqYS11puJgt9BzCKyiLLf2g+QVVs0RKp
RTe8QSDKSSKBZizt+On+CPM58xAzrp6lNnA9/va4y2rBL95qnvGB3b12MVZXgX7Tc0jjj7+nEp4Z
ZorE2vp1SURmGV1MHL7Mye1vd745qSxC68EaSRbtKEt2MaIJtuK0bR6jbGTebakh/8CoVivMpTdP
owxqQACnmfaRTN7n/s1fN3g/1EzdcVhD31OXgv16/W3j1oH2lFLtkXNAUnggg1G3JA+NgG4KQ/c7
BVXUwu7hO+WF47XXlUkDySbg3jgjlv6kvddVNthWCZKqf9HlHiL37QZspN5NhSq6w28EWds1LBZf
MwoHY1cpfR46WX5s/XIuV4bnlgE3caTqDL7EnC+h0iD2kAH6by7L73OLyKi4JvPl61lg48qiEmAf
IYIafF26uQNnLqTpu/607D8IhfsEQ4vXDHhC698ap+HKWwOuGdPsE113kpPRIUgKYPS19HDy07E4
/LA68oLc4m6oJJn3mF6c5zBeDehkktaFroWrCxyXQZbnXvjBfulJfXdi82xmyr5m/sRsQXQTSs6g
cR1CsgisPz7kwfaLh3fBOPAxJfxK8HpJktIbJCNA6KaURomNbB8k9d8YxCSrTclj03TauN5PX4Z+
7MSEuzGOOiWppiA9J1y/+yPogt3JdMq5aiUMxVT0/uGf/22NTXjKOrWlanONq3mVeo/cViPO2DaW
mc2l4j/Zfn6HSVdDYNhfIeMmUmv1iiSuznS/WZXdConNEunzND5ziEVtJmKJob4CXeUAVTbHZ0KP
Z/6l3cj0PnrC73OpkwRKrSCJQk9JGerjZKaL2mtusIvceP7Xk4Tz2oo5IL3jot89E9RyCYa3Lggt
r0uU4eluCcBU5vY22SryqslRAfMbw+GLCdq8de4wtGPfW7+VYK/3U9+jf7f3VnrxtxNg9+LRSzn0
C3lHOFQwg7Z3TDQ28eQnIU1ArwMCC08u+8auL4en+dGa4gBgLL3fmeawvfcP3UUK4HocYBQBACI5
+kqvhGGJ09HqHcE6EnXuWQLCuKSd9H2OCHmEbeJ+x+1ovbFpWRHaAUZhJ2JZaWzrnHe4N75nUQiS
A48xPybdCzsA5ZmImmJomHFbtldVjf63iMYEiRplCSmd2+kER50i8Eg5z9gQlsUsfZLfCcqUEqi8
8hFRNAR4l9Puo5idnkUGfosvx4EjCPS395j9KNt6TRa+aaXxMY3rL77rcu+kYZQ82ojn9x5HWBMU
EYAaE7u6tXWuoWfAvs9ovoSew1QeTuU6IqR9vhzMebWQmVmEnxyAle+bXsL1a8JKlKw5hdol6uZZ
12SF6gMYq3u5nScVBKqF9soR6qlLpaJrW8lFxCvubl9BN4zNl9EAMa8ymuLLMRW0aqBC/1VNvNsD
d1hvEo1GKPBGl6S9uPsGCiZVcQWkaZtdF+sxCTPkJ6DYc9KrGVoUq+noi+CLzu+7NQuygw34r7so
+esfU47C5QVEYzfc5dZ9m9URpXX4rGdcy8NjGUQYVo7kRhzvDspZrQ0X/GqO5h8fgKcs395KzJG8
q/XsKtIXOCq99lbk8WbFrQi2tv/jKG3fel9kJHdyuIY4BmpWe9QV2Du3qsw/+LoZFaWUlDvKvl36
LsR36xZJzZAWsRCRcfuoQ0UproN9mn6sUiZf7FxhycaRewvCF++PIn1+vF1ZoKlqCTWlrKYt3vdb
/VJxr+OQwmrk7+AgnYUJdjpgf5wYEcbj71IPu4GsABsBLYufeDyjktTEKtMvemdQp0d7YOhUkKti
btMsqlkr0aoLwd2JI6V3HnRbRZ+5IG4T0rXHX9Z7TAgvVl2LRc2kAg17dxvJDbhlgY0lDt4oQTZo
F9mDDgkmTWnQcbLySK7BrqQdv9Wja2ljzLJx+w+QY3xqDnMa4w5+sDeRjf5AT9Rz4kjyq4QbMFZx
UJrKjPQ0t6/l1yVPtEF0P43MUPMMgNEJaQk57pMW1AMALz2SObHp7JWzcdprrD/uo21YkkhFyODm
OJgttqsDUtsnIU1sPFv1pcX9MN5IpzDXvID3p28VpRPITF9BGx/whIRyWOLZOoOJe8Fj+Eex5lZI
DX0gF9YWVA6OrkhbgnCwGUtc2D8ZGPJbdIJG2A0GGoDa+X/j5/qSmeZEs1ui779lI3Xgijh8thNI
hYik1o6W9c9ppymX7s335xwF/Ddn3TNKp1X3JKVapvvgI2PM9EPPEOGQu+2epfQchTIpD9xjdpmp
KFSMD3Gpfa2ymWEloFB+um2taUF0C20Rci3URZrxH2pBv3MYORfDDB+TI9ZzbvEOx7x9tx15d8SB
1m0u/CWdUPTsH1vbv3HJUaESQAXN3esMODKxsBg0CtYRtLUCsQGtSFG5dPk/eCn6RxTKyR5L8fJr
JEY3+Li58fEXk8AQVPq/8GBAxoBEkL9Q3zj8gSqDpSKtkF0ZRqX+Tdi5SRnrNnMj+3qeP3BF6JFt
J8KYMBl/DaKWtHSySGJ4mRxqbsAcpNGW1S93GYcb7NHdMnR61Mfqj+Rp3O0bpPB/J3Brdbc0qzkA
tVkvqdgHDrQIfPm7xw+bLncQiEDYB0LKghXaQrZ3Fkx8YjZ597i7+uo3NdgCN1+IOarWiOhOXHUo
72MICR8nXAe1JjBMYfJwHtgustP2W0UEXy15X6xcUxQK09VB303RQl8wtsdFEU53WUd+5PMrc+Zj
8N4LrnEI3HzasorSraAv3YiFAEV68JjF7Ub8YoVeDetjTCzjYE1/kd0LCeNbMRLVMhUQ185VIRgT
GdSpIsqDQz6UYi9mxDdVpulYZmO+P0wMyArBrDiSRlTFiwY7R5kOPkVFQmGbR/pHmg9VPOSoOKX6
ZmhhVLhlj5tKhvLYM559xjn+d+8iSpdswXAI6VWm9oe0+wgkAJHNNmNYyW86sxp+plBKuLLYNgrf
rTLkJJJ/APEFTG6MQOBuZWLSTj8HCmZajLMxzOLNCNjoBY3HYJgw/sxRi1THLSAyooUAz3PIRSXm
4i2IAMkkf1OLPVV6emgssp15X1ox2Fxa+lz5rNxF3YhoFUTItD6lVvmxnzBWmsrPxMiC5e7tuv8x
laxEk2xVGuaVvIaqhtC5Kt4Kcf+1IHr7dmWmB1YhlbWoPJqK9MZuFdQ9qJOssPnDQAl7H1wLxzaD
8K4tkyumkbF1Iw9eJ/q1BeewWArU+dSnnAK15pgp0viRw/WySRxChzlGCTsmp17PxjsiCsA6QoN/
LH9vQLZm8bDfhJZ9e+ERyk6j55WflCw1sA+AG9w7R9zyoHM410EgBJjD/+G9p3ToHeWCJdvkEAo/
3Rz7b69AmU61MvBh5VFzlRxr1w+0iP/3FebDBaB3KNIpyJM6QT/Spgp/vPMN5S22tmQyffx1r0Y+
zEm1sDVDy/ka4w7RnBdWHBJPJtAA6JC/AKsQ7vhkec7g/rG3UcVWKsC9YnMSfZZEE6KpBBBMWEIa
1yz0JaVXgFayxIWz+E259BMCgUSGj1WoURD//fkEiywwNVew77UFnF1iD0xJd1sbTXC4hDo7TGK9
Bs5J3XxU94TpdzZjKz+DOeyurtV2s2/m8lRAPA4CgZQUqwzb4KI9nxRGEpySDN8+NtGUlI7zf5av
kGRZCFYLEB0fvSbJMgHRKe2BEB0IfpxXwkP+0dZ+sjgBD6QEkA7wQDflb9KT5y9hvOOamMITCDpJ
ANK8LhtlZyES/Hd4C16O226xV8/wA/YLv2aXL+flTMx2ovqSO9hQk8HRID64550xzRWT9IFLtnWi
NnBbSR6e3uq8GlVPojWW95GsW5NJJ74aPpWdBi5X51JtvsYTgHLu9d7AqKYb1xCM0mSq3OgQ5kIg
D3PaDmqQkpsedALQlOOJLgaZL8uoCwTXYgoZyC5eBj5mdQzmDtjZBFMxvDntQntY4gCvtcMRVB9r
TLSx9YokZFbEjf5zBS/n5AmYYgC9yMEDVsCSIk15ZA0VnLCi1DDXGkqUZRb0mEy77INk+Egjq0A0
Eu9k3iuZwxYw4QMttbfCer7gBsFzXGqjzE6kW7G31+zDWZYFuSoBobXWfdlCbFFWhYRbC4KGnM7R
Ax5yBWqfGMHyddT72RtrzOOadhvjaZinOl2O71N7NoEZIK8j6XTQyrdQqf93sP2LZ1l7MTUeXIIe
abapfLBKoiXq4GCyqWCtGbhcPcrmpXJcgRdjkt+VU7ksPCiUq/X+F6BwNn9cSq3IEu6Iwuismo/U
cvfH7XlR8lR7kZdD/OhWX7tmK2LP6QWK/MS48EjzInzSR3Lgj2NlJjXmcrbu9j8GsVee8Avn6WvA
W17I07E8HHY8d6RAZ7dG5+yDs6JcPEHsav3I1OZKhip2O5p15cO6FZ/VlXfW6DsQW+ORUh1al8PM
ZqJodiWk3c0M762MutBgSWGfPJot8EaifUiLJZ1FnLuJ0k7ZXKkTQ/5KINLB2Z32PG61djuvtf5x
EwuoJNOn9uMH8rkOp0j4lanHNxwDafH6fTR4Ghw6qX9Kf5GBEYfOaW3PSx+Qo9Tak0s5rDd0opDU
5PwmyUovhqtQVNaZI7xXZkxNxIRq4kdIP6Za5J0+5gygmLT/WJrHq5L+ybqUR8dCHoNFY+/pprJV
XSIZKS/NqJrRcsLg8d9CnDUXVgeFYllalqyLVMWJd+LECEWU4vojDsw2EWj8c6ievSDTM9QeXd/J
6NEsH5r7otdbsDY2KgtdQeAijPg+ktG/Nnv/Ma80tGoRFSy8a9Cqhrky58IsJO4xwl21xhswRV0H
PBZafhb8XERahcZDKN03poktfHpGGGYU9LzI0vAZXianwbotYdan/H5drU1NnFtDwOQ4bfHpZgeI
cocInKJa7bHtU/9koEnnaBhTapiy8A/V5AfXljij0RnGEAVH4+ldi1h9bogAcTp0y4+Hc3hnlJqf
3kOczr4gDz4rOfrjjlgKGs51hyNp3fZGH6dpUhPvLKcXak5g/8+S0O5DNX5r3bmdLgMRm7NUfDb4
CfpGvCJZqNixGDpqV/qERy3RrGocvOt1kvfnz15/6QvlkcRDIOwPO7ZEv75XTuwovF+Sa2sjY3lg
O879Lz2ZyHJP6TwclqoPRwditJk3GY0Z6D4gTSxHeYPv+1kI+rodN66trZRQmKCZ/avYGTitJ8G2
tzlZO0T4U09oLt0U5onA6iAlZ5gPDYv9o7ss/PYpFI9HXlBOMlyKUDCZv7mVxdSTSd1z8PYxXl/6
GE3zg99dTaMqsnL9SB3IHzmHMDNnKbJm2SKsz10JU7z64IBOJ7KU6OoNSaaBcYA/Yj8OSQibeWdM
R/+Hwk/iZLmZgqAU9uoxSrAFfaE93mC6k26rIFqvmXNPHKEkg8hrz/ZP+DbJRmyh1rfo2LuViWNm
wgOM4YnVvhucENHPL/pF0bW50S7yK8HO0jmteUi5NBbA3A06sLnpfMsQCxV0hAuz/pakveMUoPNX
AMGqzPuNSBdzMlMCli+ub9qVyum0uK+qDG0J2Zpwn413RsZjVVup3/QT7htPWmzcy4uvAKfOTVmB
xYwHMm4lEs3xBeTWNUneQ/zANE5LHsDIiwobizCWHkoSEme3GqlFgWsbhJSNyUkL7qS614mbt3Zj
KB7vlHSehc3DIUrtLBUfHj9vhgFb2gbnFEmgfj4SQRHipiuP0+5iHfqDul8XWrPpqG3a2x1W5ctC
CsiYkMRYRB6asZDhy/Fy5e+Qtkj9c8Fst8otjuJonuXzCmSo7IxyHkleyHC2jobBgvaOTvydFRGL
SCZVVhuSnxylCSfRoi8MhWhrdGae+Haa7hhywPe0wQ1H/+Bdi4600vFOEo5br7FXbFp+MtJbNXNp
Hrvl9uN13k0pNWalAJbQJWo+aUWAMbdghikyCBz/Ux6qp9PqSeKLgXozwXVCvWheefrZMIxJvjIr
Maq7N91IQ4ByOkJ+tqNieTXQuc03e2+K8VWjaH4vruwyazDpEIEKhhfi/NR53JXAfRxkJXQKmN3g
y/4QYaxdiMgPn8IC4bDO4kQ7BL6y4kVF4QZLwcPhC6BR0xT+L94tMo0+bayLdx42wD4UgYFoeVzJ
XoW9Ev9Ad83CHQ9uzBRQR0atSQtGzv9EsH+NwV2lBCekrGtxwtnC5s7c6gbMBysMTsKFX/VwDHZB
EpIu8PahaKztT8zPNzsB7dA9Mln9BhuQBSWlkIdL9AwGji3tdRZC8+4KpQ7JhXjmg6cY9OKp9Sar
cG2Ov6q8tHZsbe5nkFOPkYJcufExA8vmiV76xtciZusOK2MpuNjvPetARDs1HPmRS9uvrmHEXCgM
auJm1iF1zVfp8dqmxrRD0J2OtGTFMA1AQmcUG3CDFOFuYnkpvyn1pQ0nRGQzlQm1DHW9A+vHXDfb
2sgIAumtaYya2fsQb6tSB7p3tbQ0S/39iBfz8uSU51QcrVWfIB0HzWgfOXKmmG/DQL5NKRp593Y9
s+j5/FOsTxULl4dUkwoGucJfZvkOpdEzIjdfn+t/TWgqt2qL6WiLDULK/LGCrX+fSlKkgY3TGQqC
o0LVbuyK8vittbDYTFtEaKuWOLjzRQ+nX07KSDm1tLQ8r6b883+r4NUCyi+3GrbI808T0KquB7LC
BhhjV0eCysQ4Oi8eS4Rfw0zvtbTreMO5PodYRweXMbHNzeWMFlCJzYDYeUmdk4+7Xyu1kg9OKZC+
VHkHIL8CfZjp6lEWTStyuuwLYnj3mk/rEasiP+RvITGWLfpeb/mspeuupwmdS/CHiR3YvLVQwHK/
43uCfRdu8IJmOTwZHFYc30z5eshdnD2yLWf2RiKY1jcf8/rAM6J5k79h6RYpCRtqWT2wDA64prWz
PcdbmKvdJhm5Z4XKlMhoBU3fEU2iSQXDtbuj+NYdcKVHLZBVYnI5VMUhGj5lCs9bOsqsbNlJuZ0G
Jdh5FUFKk+QwW+9dA3B3hIS43l2MmqjXr6jBGe4w8eVwSq4VwUB/RcNNfPFQIrMlLPDolgyHRuUH
f67lpZckCIDAekFNnVvLmWnjmST+tW2SnwjGYlUFKAbnWO9mQy9yAr7J+fVZ/lD3SHVqiiVVJsWo
UfvteVJ5wcdNe4evZDD/lMNIDFTwz4gPUslJCfJx00sPaVc9+xb0Jv2FezlcdE1SeMkvVJPe7Gij
LJqAoSie1K0a3X/q0kibYglLVNgKJW14NVTr3a8GlPXbjlsE4nbYxWlYOkEPGBnLyaHG/i/f9zc/
voc4z3Ti6fC4HGBh1QbvvTZezNFLobRfYmL3GL0IRu1DL73FvOZ2QEKF7dhojkA5u3C/XvXoIA0x
he37zKSy25yZwlNmBCD0a7BniIwjGzrwHaJOreI8ipw6LvOHJYebNlnE63/Q/qeKjAjTdgSuUMt1
tZGGSae4SC058rUxyA8H/3Z/H9/wdT/e5Rb2Mofn8Wo7PSwcFYQ+J9V/4RtNxsj3fuOX8VhsAdT/
YGRnFWp2QYqse4dUTAy5R1ZUY1voPCH2ZgNvNFlh5H8rpzvooY1YqMYoW71XcAJs25jo7q8muB61
gKSGConKS/Ek5qkNKED4DsLzLxJypTERzjyzEzy4dPQJDtqe4YNULsW2YIeUby6cABuipGuKet/9
N7mF0MwKFXoHDCOHN86jIMqPPH5JHb8+9oQJTewB2u8NKMX7j59F5KvcLihQ7+0wYTdIkr2p4jYn
XyWYkwXDVdQ9gy32ivqO5haB6x1T+MQtQELSEbsg038SrOW/qTLhUocNb/SpRo2nCHvAzNa2YofU
+GiyoUMYT21rAL3JDIGtHWeBVnHEETjOpH8/QKmNEgvfoYv8tCrckFi+U289o9oKEdMAVE5+TBCc
RLIvVNjGNmY4eJOSRNnjIaq2yZSN3q9LD7RxTlEFVcDENYSOUxty8NrU+99V7wosl+DDHZs1ys6h
r00v3ljFsCLnx7BpAmGcirhz0bfYujfowFfgfs+MWivUtwfJSbaOP/1Zgnkb/ibxWfSXtvib8vzM
GFBrIYA/JF1XrmXT/IZ4Cn7mdvX6g1M/JRK/+AzgFWb8JAm79r4xQNWjBEH+qbS0bnts2UroL1+3
Sjkxk0SYMZxqNBNtcBn0d8btjl1KnWXy6VMpSwvc2DEJLpVNqWL9oBOwmxIX+C8T7e9m+hwGKIVo
Sr4aIlx09meAnAqAjfBkVHW+cQ6rGj1ijfyaOJubLq+F6CRSRPncv/CFDVsL0M7K+xK7MRlKjnMu
9LPlieTbXGaIYAa3z7Xw9eSKbHJ+fqQB9C7O5GMWEjIl/haSqA0AGSdWs4+ow5O/MSSLJ4hjBViG
knVfw0RmlvIeteoUUKHubQUl0Zkdn1hRX1FlHnEddMS+DASgY/GtGHnAtQfI7XFd4tl8txELwqOD
PO0Kb4oZnan1C0x+4SaC1bcxnrXc5JJ3wdaUexRpwMTul75jGNRmgPLpfQ1L5FaN/Hz2J2R+xGuy
T/TTKMIeKYUPVt/vU0Kt7+t5wV0ZD7RQfwrkfXQqMCZ6K/eUggvVkrX/m3HGbHMwfltuTDQQIVAV
vbHIxq5V3zBlV2OK62C6r3F3hFu2yhou6I9LvlEugHm3E1+dRcX0ZIz4VNNxYg+ClRLHnw23RSt2
tfmB/XjsbWz7CInM0Uv2/7qYdz7tVFxOr1MqQGyZkucMV71NhyQ4YA5C4khKclMcfLupP07H6QQL
gNXSxacCcny4Ywgl5MymgMn0C0Q+1Rmz6axJhlw9yn7h/tMsqY1c/abu7PfuZsT0QkhCeOsJc7l7
olTToLuBmhZjtqHzoxeVqJEHayCqu+L71ORSCJqxN3A3uJbv+45WXLDCuF0c9wyBSB+UvhuKEtrg
X8/OH1BsFqY1gxCWzwbeyUbHQCxUuWr9zQAvR2Ms2jj8PeBjsn1z+dJLbu+b4zOlqITZEfInG3s3
A5lhHuXtsB3MKOCaL9RQ1UCrikdzzSxYKYB/sTtQemMtNntddvv5tLJ068+/OCU9XTVINBqyiL5B
M52m3JlGtSTD907OoE2ZFh5IalW2FeSxOtuljlSkEQ+sXifSlE1SEmRsf04WiGihvjG3B0iNFGXU
AuJsjoVvzGfgnH821KHNyf2uSsErLYL4SS/JmE1NL+hsmio0M3bTlkFGP9kVi0b9j8+9EReMYI1f
z09zwXzincdQLM75uieSYNAD8y3VsrdEc2EfXfQy1v2SuV0ObR+2nlr5GcXKM8hhBmRAPf1xLTue
3eKsaSXq8os/oOtpLGIv7QRuvbsGK9YSY1faofJvHM6aI8jRKB6MRYTw3RD1AIqlWL8B9sl5ppfm
rFjqy50GzASznxMNtNEPu78OMEYfefUDOCf2gHl4ZN3xZG9mfggk5SxQ/Wtnl8ubefvQPmWFHIDF
uNj9CVV28ctvbMtp53NaRtGzmwbltYBhSFIx7RuKpwgjsmfRWTPUa36Vrfmx1jhw/ywNlU24PCM3
Uxer5yk1z6Cj+lsgkE4I2DXCbTo4vC6MmHOIlplpqnYbsJ9NNQAIqG6jjqDjxHb6Lt+QsqRtoT2Q
A1E4sMLxpz6hE0cpFULAFj7TToeIoiJs9jGmYD6GCKp2roJ/JvwGaaGBk3zE/0wTYYE+Kd831Ea7
RYQ+o+y/iBsnmoXKONnmC9j0fKMb/jZ2pw3j9kQwbDwXlyFs+Bw7N5NF7aZb3e6NJCj4R4KjWrWM
haQFi32w8ABWXrPdTMhujP1EjNsJeGUrembUjehZEOyVyhP/v7xO5RdQq5DROiA6Z6mDf718IWWM
llJtlezG963Qya4yjnUdoNAt5Zpq+JEjxdk06MyJdFS/k0pPy8FU0Mwz9n8FzoD9BMAlrxzVzQ+G
1pGMBHR6rClXxsAmt4Xx+YoJJ8c4+cVG84PISGlJ4+09YVwBn0G19qmP1qpbwqlWpoNAOMg5LHPj
pKCWnNWp1bxkRHtxtMxNc/FDSQuk2oEjtbaeIXAmfsO9Xt87NhRYCSNwR1pQ/pPfcW12DTu12Jy8
HCdBok1SLEWKySvqNQAP1xNuPrTWEg+w1iF0g70U29HpM+bsbIvSW2xhGogSYti1VlYyMDQEh8B8
l8XguRO8qG0nCymUmxGLlWN+5EQleO9LdM3FMv3Du39OoXYEdY5BhPM1zQpYmTWkWJ0wMKSg6YCN
SaHb0YY0Bukl3TtyDaechmhTILIw/e5ZP6mGTpYEYhNMpyUy2L3WCpNEamS0V5HqWNsTPD8lBrMO
Se0wCxFDKdTrxt0g5tMNDIXOQ0RxSi0G5LNTBTLAAHOMXcMYdlAL/L3n7gOOdiaLe33R1Jr5QO7N
6RWX3TP35zaAN5ij45lXMey+8IekI/AFBr+BnzuMqZ5W0SJukkOOmaHuJQegs3LTvs7IuEmuWy4B
eih8gaMarYbW64JZls+qi6vh2YT31vnY90l+fRZcsep5pcc6h3AycY8unQHREULRBBoN+tSztUoJ
1y4k0zHKm10D6ZGTfvd5LqetVrflJ1Ra1qdj5xLY32AvGYdcdmIGlekQdYZD6wAGIb8KaZbVUCWo
7NR2sKUzf4A3NTjeN1tdck5SMFtWJSuFa7GXNKMB9cQuHZ7rTa20GqIC4gdfg2Wr71DxuVELiUPr
hQVSQdzNT2N+GJfA0UNk8FhzMh5YoGm6ukF5L2glXwbvr6trCydMoH3nZ9M+Huz3gcabR5ec7Jnj
rPndC9xtFdlstF0SY6QDPh31bvKtsChdRKt6ev6//KjLfhK6jpr19IY9O7j2lTWB+bgyaPPKDBBH
rTGCLulcqFZ3idc+r9l3WwfEygjNoQFz4Kbddx52QU6JV4GoBdggJXtUwVfJOVrlC3plkm0cbYr2
uBP73HxxK8eOvlycPsh7OhjPwIdsoUcnkKCR+ZSY22AU897RsxLVXux7JnJHYK7xDNJy/Izn2DsU
+ziBnzrGfW5F5URSUbiED+XFefukt5DQf9Ec1ZkDfpTeAZ1TKB828JKYtYSuPCGfAuNFVE79cpIw
gTx86gj5bAcyKE51OBsuQLh+I/NIRZP+/2BSFti2Zcb11bJ9VvdUCn50ZjjfHZedKF+ORSJBgSE6
IOboiNRWUsR74KmZwb9J2yar5cxQKSMsNCbIYcJVkV0mHvyBUoGYVDXY/dkLHwaLTQLdHxpcDGgs
k2U+/PiDf1cVdiYWVPV8t0h6BKm4jWbkRZ50csZ2GvaVDxT78RCbbXwhI/BHGf3exECvut+rmcHC
ZoBqieqvXbeqFK86NFDzA+FHjGUG44oNjcn8RCDHwI8N1nqVHdY7bYOwHXQ6fbnuSbpRlE/wOVsB
MhHtui203sIPCvBVZRN2nFHUuaAAu0JUWjV5IPT2HW8/ngwbHrS7tvq++b+jiD+dyVQMHHVvIH7o
5zxleAP14aJJI0v9Zw4bF9w+Fr8ah9NsiAPjjTpyv/CIA09HDhhZo2DU4FQAreEEpnt/5lVsrlWl
EBSLU42KFWDDPTbQr+7mc4CSgmcq4APoq7/XD+vFf1aDhLuedMLh4nREe26GQhN7vAg/EhQJ1EkC
EUdHIZGAkgVUvfMITYuSOXNB2aF5kaTpM76jJb5xqFMdcITNiiTtHk9Ul3dLP3cKEDPWm515tqCW
SRergSq3U+zyv17C898/YCbZtUcbvjiUdT/W7C1HhGG6nA7+B9auJ6/LIBfxfqzPvl5FoRkHPV1q
BBr+FBeWaSJSvxV3VrCXQLtJqsCg9J7moa4P/0YiGt6jpH/RND6YQkW0ThrLSiBCawWJf1NFkCZI
q5AI3OAIz9ZT6WtjdS2fcNt4j23TsrWaX/7Cpi1spFUiVW1W67RAJ4gP+vB+oGITwj5iIIjcSJ5e
NumjWVYFzJpZ32fo4KhYG57s/6w62PTLqys2Rem8qo12555YtPRtUO3+3K9tRundkXo0WK5kfUJQ
k0A2NIiwIZRcqmvyH+oy3etRl17NhGGBG3tx1ye7uQxKb/CSO1KHYHHVUH6Wk3P/JMTfB+lmtdEK
O34JwN4mlmS4iZcHwqEl7zXB/QPgwOdc9Ol9cytZKP72uyVm5xozFdVqaabgGKSQaqmDeHmc8/hd
xKFwQRpw9N4t0RFE5DrZgf/lwlOa0Wvu7UPQAamJZQIBSXuLaQdKSS3FOB/K17NlZS5SllVffFaA
K7Js+V4svxB5FWf4SVIOhHn7YeifPYAcCveGiFyc2mGpO4ESE4CJtdz1yNASWyE6g/705A6w1Xiw
ltnSWYxP4TuDb0Eb+Tk/s3LaSs9bR/RFjkVQKBYrgDB+rhjGX3taqDRxfxEjx1xT3jlnEzQX7Hbs
v/GW1/GMj2Of81ktFsM469z72iBJmIiRgGs2AXpEgmbqICJB+pSbhhCh5vkJgq8NxF0fZzDZVizZ
dUBd/PQxIn3Dz05rnZRypZqSNzQO+hWa5veJ7owmbKDmw5b8P20scWMr3vdBjHkNbThn3H6inw0O
autAYi83MyXBf2Dp6fjU230R8XyHyVe8JG1RncGteHocyoLRTuHV9ua3yvCpUBBaGapM3TvL1lIB
b6359Wh25muXWg3ErWp8u74saHsIHZrVlNHC+GH2p5KfsgP6wl29xhDN2yqWBNzSBXiFb6WeXokZ
0InwwZ+ocby9L8kQO86sAWqOrXAwY68WOlCeTh9WD0B38CHl7qgEow9zctsbBU05xyqbHXf3/7UL
S874pb66nkrb4235joP8SAwpD+3hoFGxp/DONsW7DfYXX8sTTxKYFdixjfRzvsZCBFvv67WTQUJO
NrH7nPdek31yotj7ud6LEzSd9lwL2i30U2klaoR65hkQwGy26K8JNv2LN7DdcwBEIuDgUGgUqJTu
TeL8Mv+M8Zb0HF+bjKGwnVtOOt8YXitSziSln/8DbFpe78TGqruVzPONq1qboWmsXScwsjPlzn4b
CFZX1VImwbFsoEL/DVKXAZx1a+BnmLtmDp27j5nijAKRFsK3tzcbmlRFOPGeFRWTd7eTrGMPHK/s
rhx3guiTnZTK1DyFSFo6H31J+7PEz7oW/D71QLv086unL3Fyftgd5Ok0YJ1lxQEwmYGc8fP51kiP
XNDhMA3iV3jdjU0M+iJrA+tXmHcjg/9g9we2vlaS2y7tp54lI4AN5ENKRI23HAtYwrUt1DEzC7c/
cprwjEy3P0tKe4HwR4wZFq/04YL9rnuJUxHo07xq1tKfXb5/6MUu9fCwmWOHcfNvxHfFwdr/+MgK
RbISysh02024HgXAsQIattNIm0TtZE08PYisuVSKyH0yXH+Uj//kYR1S7qQBGvxEZ6Zg84zpdTJi
OnbjRSrOZ6QSXWkx7fZz1+rStEotp2KUMI8k/tIAtjNsHL9MhKXg2r41A3DcVd9b9gZBK4S9uk1p
meAnn0xhxJS4yhJLgaPJiKnT6dMHBbLhFr6tWbxa9DtG/8MqiH98InDgh0SONWgzY/ot+qyGWUby
bhX14awfMHLgdk3I0XD+dpYUPPu529i1l4s+8bHBav+TfmngSa8d0cIehFKA1Dt3ZPSQAAgjo6kS
7ecO4xZQeugcJ2Iwm2tFL6QeEXC8VU/Nl7dxh89SbK6yOQLXfrxnQswEj32iumbMio4KDyvBndaM
BrIJfFb5pFIaR06TsIN3YdZ+wc94U3mY9W2CNC82hzqkcIe9IXh2bgU4WqIEftsb3/eLKznaNd+h
+Syiai/AIXu59ud0Tjztws/kv0dc7Sb+JyC579rrGb24891HZGt6KixzS89ARQT5vmZBkb5tmsTE
GcYdzRdfH1by+NkeKWWt8GnVTXqVxr1sEMvdwAqrFnDixqr7u0/5I2ZzDJuTPloFe4fLo+CWoWok
uk+yoTSE2bxRQw+JO4VvcDOae6vEzbeNXMU+5mQ52bNvUudFmIoPCtVVY1JbgrOAvTLD4fSI4p6E
3VTJUXM1xks5GeL6nrT/bgFFtOvISt0WD4g1sMwv34B9YLE+q5OsZAjmGGOllhCfoJyqRTfrgd5Y
P/fzYpP9WEvf/OZQQkSIBEDdRzRSPQkPYBHw8iJCwUWGNRbSKu//gaFHbQTT3nnQXXJQ9mpxMQdI
bIdgwgTDT8gnulUYA3XFPjnx8vmeBb4jT4N+B2yQHJZ3OeOOKawT1EmW5opHDZM7j0gwe2StvfnR
Q+kCSOlyAMDAfrFF5Mfv0aCph77ZMqT9wuo0/7MkSVm3tnuhkVq2G1kv7+gOMAfIi1jhUM24njwi
Fj5Y34DRz7XTpUkF+42LgF+HWBozlnKcWg/1D2K7axqwj+yEgDrBMmUb4ycNhLu28dBdP3tRIrrd
Eua6H2hAtgYk7HfnR4JQQIdyFe+ijKn6zuwAjAmwJexjTJQSir6/pVQqBDU/unVSh8qrz/PZFgY3
gYdn/0WhY/g9kh85Lv7vpLmwcPzyu8L0SFUOi0QD5jw32CvfbrwIekdBJ57CiXRI4bLqIcJz09HZ
IshG6c7DeucZgEEjCkqIYfZ9nHekExkmM/fhK2chvudYAIlHr8V5tLpXNps73r/tOPKc5CkvWv5F
kKmrB4gVAlzcQBD2N0IRYNTV+CHrvruIUgrHnnGVtT3Orbrofvs29BCvrQSbuE8Us1nJkKpD1LRP
GesFwJcDDC9d7ZzbP/LjJauV+fKjqJrfe2Hr8IlMxhgDeLr64uwL/iISwTBHGR6VRp+0/Q5nX9WV
9fXCXR+h8j+qtE3rhSYV8svNyRZEEiAHblBgnEC2kBlBpwjALBhoA01N/4BpKW28VCLJg+ZF6e+9
cPHUSZYm83jTTexmIjwBTZ1ih3ryPcLEyxKSsi0MbToV6jJoaOQoGKUgJ+PlsWDFCU1uKIVB5Z3e
pqWoghANkdMjw7YMt2TAgIPeVjJeESGBuv2L3CUlnKbOVvKXDjU3/ipKEhJx/Ed8W0Nzu5TahuBd
H8hZgFz5dFupJHjZkddWlhyi0NV77GZomIQkKho2nzVtktOQgT2xveZ+o3xl3cY09axZk9+3iG9l
XEVHiZBB9OI4Ps+d2xmcC0E+9AmOculm0HYThf/TC7D2ml/fJn0HYBBMo+HnsGGIHyZ81EKPGIYa
b9frUqn1My6ThXJkG4k8SeZUxrhPUNdU9ccJbvbmEDOXi9+MdPeAwHeszkFCKnMEfdJHV35+q+bw
mRoEp4FBiBHjQDW/fT1rqMxZdMYCD2aGH2sumgWgBulGVKgRiCk2b/2dOiDzgtioqO2I/yZ4usp5
mSThWw5qfrFkXR2pNOdQ25e+X6uXn5fF5PRDqqghQ8CtpiZIZ1MwyraNLZNZ0td/mPEj1/paOLJj
Fsxck9eH7KHmufeYMO0WTmonrxZkiflYNGSinDTc4jWvpbKmF9dKuJqEqWwjigBHYyIvlB/sO5Xo
fNSuNiCo4GyBrpYsY6kQYSr7BN6Zx+v+WkA5SJEeaC//Kzz0s5ooquuleqn1xY64XVTKvkb91Ytk
zt4YE25/LPEnm495xwktrweoDNaTUQYQ8Qmux0m9IHS2i/DEayIKkwaak4DunXDZSmX3nNkklDKM
tQAhBSRYHogY7jU2XW0EmTa7P6dJw4Tka7ELTvd4XvVYP2QBdbzHlvd2BYYMFB9vH0fMNaJuVeEE
vLphVwUHC6GLFXV9Ui58liOiTtlBmkBFiRG+NUv7TlbRVBYRSnGbCHB2fbE7CosNzus4XKz8vUFj
FBhGkltnZTEHFFdE/REUdMVTPNyZ7hTGcXE46wieeXzd5m1PU9tvLmvnizavcEd8WJZZuxz00IYu
h6qpGXhuF6Fs3KJ9fh+S+MO2SuqKTGj4jZg7+UgZs9+WWsFobfXjNqGKriNPHnl42XrVwv7V7abo
PYfML5vm6qhiBKPa3V6Z+8V1DH8nD8lnMol+JdQUyrg0Pu6nyDA6E7T3/jEWQo7Zy0W6lcdwheFp
od/5Si8UimLdVi5GTcD9w1d33rVlZphtJE6xYvQcmtuAG16T0nHc6r+CSZALdAc1biMmp660YVGM
IIyiIEpkpkIZ3/3a17iJVjAqj/g0DAxGQR+Z2MtNlPGLBdJVn1Oy2t8D78rZVNoYjyGYPS414vPY
/ANU9ANHSE6A+obBKltT+StGV19EKprYH/zKStZt3AuJZqXy+n2cg0suWozA6pBzhRRBwY4HpROi
1axX9AxTQ6PU1hncn8h4gDqPQjdhPaBLAvsF0ITqpCkFwdN0g3tbhAYRg6njBtZAlh2CGW/x9gp7
JpFVL98UUqtJG5n+iCCqzlri7AdPu3tuTLhw/noxxB6uAdu3i4+GFeddVLuWEXyNcFhFcFzuYL7+
2SkQ8UhdVZ5YPmymK1phPeaq+gZEXvHSTseCOTs2WQ5T71FgPYEYNMlzDzy5RJKDVWZTJ3ECU85T
le9Om1xtZjaU5viPfCzLqV7yza+FPKDaGU3zyic6+IcNohYtygqUUYG7GUcjhB2LaY34L5FWL10i
GDUb302FiRgJ9w7xQLufMaWrr4mFtlKWcREbozuJLMioXF9x2Ins4At7t0o97E4pltwjkwKR+jyd
mYW2+UykpqdSBu0FhYEXdKczmOAulwMoJgWDD+tHZiNuJ0Yug/bfLb72UV5EK8ftWR3NmwnFAp7K
KTZeVLB4xcASB/V4YS16RYbqoZRhmzwJUG2pq+5jCPJsx7OPle33mdx5yjNh4YuVIvnza7+iddkp
JaGNKlJRIN9MAu6JSY1cpbYRu31sdtIJshQ3vVHtsNExP2kNxOu2ATMIcEow/A2GGC4HCa6dY/bI
teWVn4/0p4E1U1R3bhQbKxEj+3G9QptzM9Uy6TbTgV2H5ikIcSHg9hqr+5wuOcbxJDIxFF/Tw9v+
3g+/JoEJ/wT38NOTZxTlh6GGaIfznmCYHkZDM1GtwcBjIVDTudQ2hGHdLmpSEFsGDfRuxR5bgx/Z
xVUJDryBggJHZOwKcixXKF04LJeemS2JLKJjkz/2/1tDCaiyH5PsJ2C98DjBIAMSqRHojd+Nfiwf
Yots027UkpCCTCzlU9C/DOrCyr5qkyFoAa0aHmeadcsWAJKsxCgdp1gS5AzY4+N+2hPIlfvNooMg
zzhuaJBDzVUDj2q1GaZTyND+DnB4PV5ccCd5weA/FOj0dU3WUDlEf8vzRVaEMF4tCWMomEOcfLl0
PlRuLZdayaicNC9/585ufXWlYYoJwAXpERMaOLREJiX+5ThzRnH3nhzfWNLQYAN5lbpoxop6wPwl
H68ywwguYZC7RLVAlePv9lbyaNpe133/sCYMPT6X/rqhR90ZW2zbPgubvriYsN3ghwNo2gw1h/tQ
2VPckq1Li624hrELLRABVrOiPYi+C3+kTUwp3PWuhEsEGjkyCciFapyZgbm+fllwBhvwaX20+/sk
5CNwC7MIwcBGxe/8kWC4FwaLaJtPdI3dpCWyR7VxPwilvkw/W5eCJMkS4YEeGhuAzZ2wQL3NH34T
iP91ySJ3am8TCjP1wuFiTVOoJcmZMVksnYcK8j+9wOkxjqTi2TCVvg/Dt+fL7BcLaPcDiUmS4dyP
mPxBH89drjz+3MFzU38mXk2Z+iveqbRGQNW2eJCd8XOfMlIJ+slAMxEOGpESvXGBLyx1t3OSUipp
RUSMq7UNwqgGOBqk0R/SQrl8dnjADq0qkXLprD0d2NofQLFzvhfHI9dSrMcGLOVb1xnQivG7/dAq
+WMqlx535Mo8H8PvTnvNTdUz8qb66ccLA6wF+ZNZyOMWj1Jv3x6e40Mae+tBsSsA/2N9dhoZy8Rr
xXa+0SCcgvzhYS4Ahu8+xNDnn2w+wMDuXp7IbSISh7Lv8IEx2qJgeg6AlygskS4Y/UWNlDIo9P+2
QHpX1U6pF+JCuO0BptP+bXES0ilfHuc8Q0EzYvuWo6UGVY3ky4A9J/qw1Z1TacFBc5bfrBxBiJ+t
dUrxdXALZv2QadGlyVa11ruBhavyBzFu1jvhBBobTA2dsHcwEEQbFQDcMxMKkrNGT9aRnHqG7pYQ
7PMPeQ4kGLMf969mR+/IRP8VfSMdwZlrr7CkalSJZeR1pqfK35ms7LC6QfM1n/Lt0xDP8ph/b2QH
1OfzRF+W5/5hBxpFdRrvLzwwDF6x1LpWW/4whd0rXvcZnMTJmHRrzzlc4y9Uz2OghkbhkxJ73TJM
j7VqhB8Dx6HFE1LmQWxs/HkDNpEFhk++Z/+b8KElVjUORMIviZjeIHsT5Fm6W4Z5ej5eZYDY9qH8
UUTD5xd37AGHpxvTqYmNMXBYC4Q/1v/cA5ckkD2s7j8v02SNbvpdPpifdhJzxOKDDEdnWpVwivzO
SJ73pjsrxCVEGIJ6LOmHYLz5t9jiNQxuIJcShGaVcz54Wl+lvpv69bg9P8fpAvoCGK5RjNyE5wD+
gQEUrH1EjjEQPbbjtSYZoHBolyiGSkqHpmCKoPWps5McUZY8xYqEKsDnBYxaQg/QJO3APP1re7vG
qBorh92HTf+tEIBjBlsp/OlRuZca6MNcGVz14MQoE1Ra9HGXIyLVECtTEiV3OL8Aq0kCCyjkvCfA
TVEHJsSMDooP7yRnbUpFWK2pDUatzh8zy65GjOulNkH+zEVmFc5DicG1mGIkwEYlMfiX3VHZ3ddf
RdGE9JhkotTZfb7MmpKoASw3NHOndJA0SqUgPYFQGvunauXzDt7pw14ulHb0kQFZz+nYMo1n8Mp4
RW3BmitqP5jpfOjSSot2ud8LrgTF+ts0823LGdVfLdQPxQciT2/ADke0M9CXRn/ijOLoYClHHRhy
BIzQ3GwfSeJzIHGeZ2McMlhX8/pBEjyho785A720P7rAEC17HbThVhRlkBPakHhMBLaoh4cZvOdM
eExA2I68lYDzDeY5XZac87qsovmXhcpAcQHmZWxSCl1ArPyWc2V6KM8rVOkscMvhJCqOERXi1oor
V32cZe46B+S7Gm29fmZ5QkfftXWcWv51nQo66IStsWTaEddPwFD4e11RpyhTO4oVWcSm0+cEFK1j
G5hVGhWHaJtwpONMWD6p//DyoDLP0+WMA+v9vS4YrRQY1vR3yipT8ahZWC5eCu7M78FSmNP4Jq9Q
B8Z4qF6LcxXzqGb8r54gauyOLN4Ah+45bK654sOqJ4VR6v10NNJtw2YMzDPkgTYj2L7HeYdmh/XL
LL+9XjLbnWdIvmTTkXZ2tgqMA7p8CpmqLKXpFR5KsCllWZyWDoDvn6noboLRJKvpcT2E3InqVhD7
Hnv03CkpbyBBfx/vH/+CyvccdrHZGLzrdDo6NPpdZoMMJTdKCUhiKUCoLVZh0Hl4ZJyCh8s5oeNp
pXFyAM+NgI+8IO3f6LWdhMyl9Z0/96VWqFeQlgV1OFLDEpG8UOI0GB4RrnOWhm01kk0OD9T59qiL
ck49ZhJ7gv/iRuUlqFcD/j18e+jzpFdS747PBRt58cPeqVcPChJ6p+9M2pL9ys6hnmTrkRmmoEq+
37++Dn6sTkEsEND3x0RJHVaKc3WqojhkyLiglYiB3nbA30HlxW6kgQDY60rnp3zaYj39/7arJfny
mQeCW0JLoLAa5DVxhQ5DizQinSxWj35gDWpKepaczPXdK/jIhxecvjNH6KIl/J4fO89m2/dTMV7e
ihX6JGyT44I9UDsjk1yfpkWcfXA2bfKn2W3SugO0O7C7sq/PuyL6i5+d50j97Z7AeMXgKK36m8V9
dv5QpxaCRqfQIuAZTqhKiKQ53yCBn8WVhS99uFUVHfPf8rtbFOdlfi8gHjaOhqhUSwC62aMJ3HnV
AwZOvsSsPeRrn+R9TI+/AXU53zL+HX6aI/YYQPfid1OJZBtXgHi77wdwzA+rAR1TKnG4B1ssQlqz
X4BYoVq05sPMmKYkCpSQN9wT8G+Srp4Rupf0ovOUy7+ls3/gmJrvW0zttxRtCRvt7cqYChvnqwkn
svp0QUwjaIjb+OLhxlVmF+cK2lQjCF7HjdlgMCmu+YHllmZN11V9de1NoLpLQJnNoTcpn7DhDSWA
n1N2HP/7deQrr2PHpjCaRhglhZcoa873L9Ovzf1iPQBOLwQjzB3C0cf+qN1IEI03VBQoMQsNd3Bt
Rrkq7yI6nep41zLhcED/5d4jnY2ac0QZHpVjhC4WlHfxt2kU1g4lzEjPuWEi1ZgrARCul6sWaIq0
B4WtcyjsXnz+TDWK+SrBD3+xxEIG5r2SkClcHsTVoDASHbxYs8x2+mkm72JvRLQb7fqwdE/PwTKn
wx0iKjk9rXtB4JeWg8X9Bc50vXOxQxRyFdH95no9VbYVgoBYrDVdsK3UZ9GqjQ1abeC62robIhPy
fy8e7ffGrLnuKBahM35/OEM2HXHh6UaA9HPqYhkUb9QoCfPGRaXiUr/1Z3ADbRg+ft5EnYpkA5z2
jjBBoOEW/QhMypSHq7sNivjZL8EPvxihn3d5JLdixu/nAVqfthU9vgsBar4KBmcOknl6xnUF1mIH
1LC6g35NvJXCBkULvdNBsA1TRPwh/AXHTz7hc3WPn1H5JoKmMdLyoc60166wx/EP/WfCEoD0AHsE
WwGsCs+IXh8GtPwVvJgUW+9R+hUuv19k7SSV6j1vA2vnl0M+NZzUweKgkwkWxT1Huxi6V3xfvRNA
uC+C/EK9z49QqZW264UbpisxFoPOYyP7SOIbVfyCxTxw5y2MPPjF0oDze5brv5PZfDePDlskjC57
DwqtfIaRneo1lDtvCXO2VQUoen5LVTRjlZZ6N4yH12PkdKBl2YprJYc1w023i1S4obt4Sn5IKVWV
U/DIKDODSxCOMtoDfPqvnz0OVi88nTEed5425UkDWyWSvYvEnbLmr8/3S9+KjHh0enrzS+FfzZS0
s5cfW15v/+HhkhT/u1egXLPEMykW+ToChmkj9iBVHEujG5rFysj54iRR1GEb2h3sT+PQownF6fBA
zHw+vj+C/eg6UWJBqMDmLYE+nAoZDHson1ybM1cIi0msc2O7JKYnV+FnnkDPyhflBdgfhGqBICs8
0zBKO4EMnRZiFtk0ID8clUxTsx86nNFooTZSSYmJxNThwD5qtewM9KB2htNHajEaDI7V+rJ+tPA5
LiLLVNXHMjSfogpaZeScqW1YqxhBSezVUOZPYrVH98RIgAk//VmhI6bVkiEKSknqF62swEb0nb4H
w0WeMijHbVBzmlAk/4eLw5okbSFDQXoByIpn0XWA1jXs0FYs6gSNt2naLld8f9ZJSBevfQz85aRd
KuyEZJFF0zT4kGrJ9sHo/ArSePLG9InkmSfP6tkVNXTaP6/6sb8suMWvpKafUvitIbeduKaggs31
YFHQSEXUanYYqiyXgVBmK/ZIr2pog1txQ13OTFHTki881iz64ZIu6d58cNk5oDNxCaD5q1B9dy21
EPJ12Hj3vtQi5Kyl5hY8CI8zUJY+pietj0qjKk0EDMcjfSi5d1kuKjP7g0lz6l36oGKJuHrqtSjR
rzSr2LwNmcaG0lXuHPOgs8qBrR7zpjh2xywqlXKay8fpNwGOivAMMA5v8JSVexdQ2BmK+cqzO/Vi
3pYkF0usPFjgxP5TnglUUB8RtMlZMRtsHniononIKKzA8ipDKDUuvQ1V7b2rS5zcQ52oVZmONuv9
Brpe+strctcU8sOjY5tN7ihbYP5GOIIsk/NDHmMDH61pb6C7EJOezve3Aj4N5I+ETM+emfqud7jY
7kJYxT4RDkApdZ6zBOoNJTGwfLHPBDwy6OoA6BU6xKnV2cUltgjYgApMRLg0dWpRiyoxZbvmGAgf
Qi1YFjqmBy41pUCZq0KQdJi7F6ebMcvCoTRib/Fy4Y5CdFJUmfG3KBDWWl/VFK+xnhtR2VVqVctE
IhLkm5v1QIj5XLC254Y/R9LiJMUt8fwKYgHLO8m9PpLsdd6lXCSmSjLAAZT7Pyo++g3XSg8QUhSF
/fjeVrTGjJjPaHrz3FiO/cXFc4QbdSSubqEpibsITAQCRN6T6Wf7DrDGshJasWbbmJPAnUNVqTrO
4C3Zin6LEG8Sok435yVRyFWxSD7XB5sJ3JHIAZPtOb5wpuf3j+sGA9TdVRauxzKpoViU1weZ06SU
9N1jpCbpAnPqH0iH9d6/sg+xF9ocGqzZ7y1ETzSVUwj+QDi+OpL5fAqAYT8PmeLavHeSKBjxTXI9
FN0x4zNXbxOOOeSMKkl0MvR8QFV0p5XoeqbNzSwQTA5p74j2K8IqZJp2/91zCWOX3YsIMASPCbHQ
iTXgXy+RmTPdfiUZNTtS0Ylm34PkMxjCQ+/jOtcgGxtIBrV6GZHbKQIPYROkLNkiX4EfTe34M+QU
l2DFwbxS109fqOVMzJpd/pzyG4qfe0RcZsK+VB5YzY/kt0tukWkPpj4apQ4+P8GMuvW88SWgu2eR
nbgGiykP+cFKM5IrvWx7FsUOlAALZuWii/hS73lT6zEhJMSqqp2+pnxvq1FbQIp2jZpwt0od8DwF
Ch8Ds3emdLhzVDTt8rcg63kSIeb83p5Vfg1NpbsPYA6BFEmmj5xoY+xFMMib66x9VQoi7yUFWkgO
qSqVqBaRqxM6XsZLK5M8Y9ErqNGIbqRmxqxlx+iYJn8xBNVJl0e4I6f6td5RXgB8bHLhtu5ZTfos
uii0+VtLadRxMbhC3Fluj37+eP+6E1uu9cU65ozV9cB2gVj5ALCbp8MnKGbjDMbx1S1C+hSzFFCw
Vy4pBRgmYHiLhjxK9IJ01idHp6ZvLKM9/UoLM0zpYvGs89BAW5wopBqGMnQApHEWLSPCSKhFG6Lm
AHhdkfm7z0Fwog6puC+cLw3rToPYhwJHccJLEqe7GGRmOORwytGyT1xVaaIpiLiaKhurPMu9DTxC
N13oqTL41jCTsEa4q8kwTfSLmwIdFuhOhrluapYRkupsVmap9EiILim0jmNOsqAse/Zq9uS58tKj
zRYBUi3OLys+oX26bQLoqJL0fSvk+otW2Y0dZR5jJZavNuD3ye0D8ruyWfdrHYttJeCWJnmMCYM6
XYq4x041OhR++fLq6jD4JR7vgik0WfUdVxSphghfqyKof4yUE/gTJ3vpPjerJy/i/GQ1BSq4emEa
hVZWD87mc/fWHYw6O1m1cFrxmYCRwKeGSq0AcfOoxkrPYbRqKPGGT7BOH2/kcDKrGzoOHnOf6Egs
Yf2BEoRSQIIePeNFQy62j6gzdzmwm26NQOgAJMiYLXBSWC9gh1jEnl0igNAGpgVSCoVxu8BXO6Rh
MFj9mXHeN1R4pRaEHiQ5TIkStDVT1nhaayqcLBMxcrKU98AU3wxlbG8PHCBhrV36wJ5YHCKlyLmp
Vif95vMmgzu/qB9qzotEudA0auN5T/OSxo6Nb6+yDUBdwifOTY+WQfuiz/41WXBui/DcRtD6oIKA
OgnwJJ743VqGvF27kBnaLgT8i2qt1SvJoOke6k+vkgnez3e1e7NMw3EQY73iUyYGDExEjznVl/fC
C5WGviZVNhtIY7NVhiRXmq2QSGoREEllIDl6ROD9wil10+TCgAPnm2JBrml+bNc8h2Yr0JhUuW0M
D/VTog3sduJGtf60KKNRYBUZMRRoX6DLnZqhx/8N/OFld21p2BfznNaQ+ZMnPCSrWiqfBzuO0UHg
FZrBTLv/oe9Vn+L4fAI7MDAhVFMx7uljM2nkttr/AjZoigMBz47rDeTibdCY7tL0JF/CFfcyF2Vw
+QjzOojbg3VPiGx+RbDNT7jpocp7SjPUcoYXJQB1Y5bCT7YH1EWZ7zvgJ/ikz9bBxgNpfoaHJaYX
UhIZbXTFVTojMx7UEPdOZuvjhMqwDMJ3mL29x33wpPvWD1mJbEIpo588n9/XqjE1VWq9zVKjDDpa
c3F/MiukpumkfX0NkM53+4DrG1vFdS9ZfCdB2C3t22Qta+uCdBhr2FJRhs1WCi9JbFInjo3zTaI+
kiUsm6OHhrHUxq23m1c+V+eLmxp77lp8Dk0zAj8xpxlVnpvAWJM4cyYqJmYxl3UeLKENLYTe5rhp
tunDqliljc2XnI5MPfTiieY/jHi23h14lezyeCzTgrbKMNJ5ZR4AOkDRcjXO13Jrcq5xvWXLp8U6
uiQxDhgptocqYwfEKnamEFSftm9HZaM/Ovg6RcdNzd6xPsFXG9E6bj4gVJCg0Dt/eIAn5mFhEQMz
0x7vzgjh6di8Mg8JKiAc2aQweP4KxcOqbHGT9rsJ1U89IYBQeotjwuiCMt93oJFbBhmcYAjtpNJo
vV2G6PqDINASG4RZjuy7INvQMAGG/xCQWLGyWaJYI+RYdhvFCAejUn4jIKa2DlevHZZCkj57lhGa
UoktHAGqxzIwqgjYAyj7Jolrwr2ao08MUP2ep8TA1B98dWa4vgRm/GGvyIhrArEQlShwdXhVub3v
jHpz32+ic8AgdY6iVhkFTJQHmkx7QKqeJFNL07CJI9kvcNFOZEOeu/l2SATd/4sxionCAcUbWQhK
5bXCvUXgK+BMT5WHyfMzOgUiuCzOvBKI6CxMQOp6L5p4mEP6qW2QZlTHtepQ06OE1oLuVgr5aZCz
5BucudUPxZmIgYZDAblRtKyw4aMEAf3dCbMmQ6Wt1rWHdZ/mPLYijiDpfrQLVQSXIQzhebjTHpLN
J7KrF0EWa4UPc1/sCVq8BVb08UMXOlK0topGKKIL3GW/CpFfuj+edPH0L5mUvbJ5S7LQbRZrlLwJ
pXxUumdxMFv19h1iGox93iaNIigSnsxUZ+GnkELM6GsvaOuqBpJwi58ndlbJ6NRfDBq4zuyvh38z
xV2wKxVUJ/Eh/Opt9BOA9kZ/2dR+zSeJEXm41p3vHJ/RhPgX/t8XuTua8JDK1vm0Efn9mV/Wlj5b
JhkskSKAxWWVliPtNAcOBoQm9LNnMB4vt7qY2p3sYDEVUokPIwlQ0F16EpEguBUgtGqnj8ekDdHe
9J5Z9bITdkO0RRlxh+X8amRh9nGe6QezLIKn+hFVBubHg1OAihRhV9ONJnojJITgI7LOlk2S1OmD
MacpmnhpOZV1Hml4B9P+zQi6UaAT4QGYKRbdbnlEiIPwaVIyl9rGJUV05LXt92VPK/GEFcUgWl8V
ULMQncGbNMdclrlggQwzpOPhc1yHD9ykqmY8/btYQcsK8nAt9tAb9tbXW9HqbVW2Vp2rrc5v6klf
/gqj2e5VpMQJZDPuXpffGfoLbrTZ0OdrhWLQ77qLwGMdDecGnQezG+WI5am1LA1NeLxDeWBghBhV
wkb8LIdJ8WRCmQkJSROo8cFOwMLE9HTeqapRyAS018rtWuHUC5tEYKubJUVNNB6B34QR/5BrTF1V
geCStvjGUiF2AI86utikJOUWmfGHuRwT+NG1u7OrJ7igTPqMPh8hF8WFdMc1U63JwSvaImBfxn8/
oqENv68R02mruFPwj/O3q6VsA5RlFGg31mDw39z/y2AaLQp9SRUyTP1amwL9B9Iy6f1Ah6o2eyzS
nccvlwQuO+Qqd3cjPDeekfaZvZx7ibkSjLhTe03HUKHn/GHvdacU+utrjNWnPmiP6Hft/BptSvNs
dy/NxM2Kei4vjGXIyKmcAzJ2AyFooIFaJxLxVpd7zU/wlS/6Iv2rr/JrFTb63wuRMVzYlEnT64HJ
481k1qcjPv4eGqTjdOZY7X8qIwDwVJASCf9eqwmxBjDbxwS93i9J+A0VqinUGEvvkXh1d26+9c8R
yspYXnIIbI1A0sSuRiJqtAqs4rfBQ+hMjyq5JHtsO6ARYA+Dqw//J050sFAolIcokxBcwaCWAr8w
YaZcC5UaCst09viuWl6+HwoQ3Qq+E62bvTKwjlsxkbaNcWlRi9pINjy1aWnQToIu3IrMm6LSV0zt
sndT6hICX3nmSd2nZV6JRm5v6+OOGi2r8qZ2WUi23AtL4cgUoGtnEpb4/o//0xZui6yEg6xYKj6E
IFRhW6mpwPD/w1kT8VG8ARgywTRQl2Wh2hYWFcC2R2Ng3HMSCK/7NScRT8wsU+bG7EUkKd91zf65
n1UxwMhvx2sl/zBMuBgtEE+SoaxyTJ6Iu0Q4uHKRrJcr1P+gsolnvojQyq1iIwjtR3sgOrbXhyD/
tq/bYeOIiGFv/WYhoYtQWvj5O2QQfJE/avoCuEoFUYc8lvcc3vXSGErB/lpsnptadE3xZiK26GNg
OaZBfWlbHxAKnqZx/TEUP2D72TgDfi8eaC5C1mMq+CHjoMNnyG6T8DwwldWnkfKb4qpmerOTVTbj
GnBeBWQH5ogVX4kcwf6iy+Sg4nDRHlmKnJT8aVVGsm25Gio8oEIY1Iw1nBVlEW/1MDqGTfQiyBur
fuRKm9rDgNseqbp9wlmZd9Hgf/EPIEDkOsVuKv4onwTx+orTuNsiurS0H6Hgneh8TspbxkBHrkSe
YhsrWKYOqqgNv481osRTubdM3eXmS8rYNeCVnJI56GNKBqAssbLJXpWo5EsIZnqA5pp6ByD15wCW
YXDL0uQ4gGcC7osw8spmATIr1rZoEgkAVPJTk8EpPAKSA50J6GG5AJ/W4ZDkgWkEwmTd8aZOSO2f
oXa/3tYnWJNfGX/6lYGxzYiabzSSf39shljWlOHr5Tjge6MBDFp09PAREhSWixIVgbG78Mby7asr
/NvMLMJ4cFNMdjrqWVdsabZ9sOU34LV46WIA/t9dfvbXOY6DJOFQ3/umPcnHpXtC+uM/O23EVQ3m
bwaJaDsSm0HxG60C5aDBcvGfr2QtRBuzulu41SD9XfyNBdA+to1xAkxTp8tgmSJEUE9yJ0aInCLT
UAC6Zlpx9mlEsn6Sl483JoyJnX1zCD1w9sp6vSGxgh99SGxuxIhsU2wekwCXYh6G6h5TtmWFZVgb
ZLlBDHMie4T/MxdpkMoFeyuzW+h36HfAqHHcnYfpPcMjzbBMcjx5Hq/vm3budp6Vq+Z/7EMjpK9r
O+97a8HPOA2SaafNeQE0wLBkVnneDXIHdESlxgPmmqswQ/QwSIwJhvr5wMiPCQMuEy8GtnG9sFpO
y0d1Le40J4nUNlndCuVwErs5gp3DUb+PYqmBtFODyFZn3XwGxja2HWKaeHjt/UrTQt6JacskzlWP
/ba2YP3sO6jlcOsI7RaP/hFMWwJaqa3n3p3H60rod4MJqzDCH7jDhGlXX437qYiJ+0XrGCr5xYlN
zwA065TnEHxIluCbLn0HLwp+9B3R4j/scuYQPJVJJgDnZ8Csz5/oSmI0BLuBDLCytpZZOlwD3kid
zctt8KspwuhZdQYWkwYLmg/rNI/ol5s8Ti2dMbcdJW4m9XtA562/jrzOxkkshMdKX4FA/YGdYyJ5
cmDdrAroDYqVkKGJ4ziQzhXuafOfkSDDBrExfoR5bmMMAmUNx7WQNImUWbMlAuk0SOEqdLZJvZFo
45MfhYln5vmWVlbwAPqhAwuR81t55Y3g8Efv+WAJTRslRhvWaEUCiKOz+3m1NJmIe7cgD36ruWlr
+ideOWOTNITMyre+HgA6uSv3EzjUaE/Paq23EuD3SdN5br7h6V7wbwdm7HwTqR7MPHlJKmvCaU0k
1oaoO42HJ/jqqBnBtmt21xi8DzogfV+d7vXtDdmWN9vv1GsQLBF2Sd14Du7UonnebVkLcN0OTwiW
sCBHlzlMGLVvZyAhz9oAWZckrCX4zH7SOnQSXkF4kYrLWCixLwMp0j/k+DjF+vxTvxJ3mif2p7Te
XodMwwJUKoLb6t+UcbLX4VsoBNN0cZ4lDGPZE2ggxk4KBzxugvI+hnWdcG6pMJjk5D68BXGulrpn
EUAYHFjWsaNb6Dr+c/FzNgkeKnidZJiMPyOUcx5IBXN/AV5nBKyeni6wPRwF8aNbT+mzhjcSaim0
SRerijoqY7YgEZb4hC2ZXgcvguNtQEr3M/gLDINqQe7Z2qRaU2Td6zlxFYoPWJ8QzNd+FBrzUquQ
EYbpdAKgsRNyO1ElhOWEc1gDtTaX589oqsVL2qbALh39fn9HBWP4t0nbG1Q6UjLOqfrjgjgGBXLY
rhpCYCO/QzwHHS7p8eU4UxoTRUYiX7hPxlZCiQ98+iGqN0q+HCk5KvyGeock6KsEJHPFiVIPbZHy
hfbxGrfwPuij+dURzFWWCT1tWF/OhtJH2FfRfPE8/CcfzSDzNxSSWTpiISGemvuM9xpkgRx6qgbW
TwvUyQpQ4tIzKhEgvEiRDvvz/hEC0oXvxG9IQnciu14HI4vlKPc6G1FBpI6ewz0FJNFdKwfuN6Al
N/H+qCVEmqrItEMUvKzmCgU11pNj/TK9TLJ8m1O3v7DDkwMeqlpKg+RC8y+S1SampdbHkpg09TGK
S+gr+CzGTeRMIc8FjN8n+gUr5vL+3KW7mVq6axBStu/BaYpgur+CjeoWPij6Em3Bx4QrWpnKNdI+
qToXboIGAO92CYbpaA3I8QhtpVDg6vLYHSGI1hx+TSMeDi4Wo7r+qU9HDxwZW7jZY02v2cNFNJsa
8QPj6+Of956zF71bhdVER3EcDyUkVXCAnWjBgYFgbo69+t9m0FQTC9AetA49NLV7Jy5kSaKlcDUv
r/Thn6HGC5i/32/5owZwumCLw+kVohNmKhkR8UYszWbbL1FD6fHF06zxU6UA6MA7YEm4u45rUuKL
RxdpphxN2t3dv2siwFwZO3NBb6HwqrkoXWrZf4UR2a3QuZ1udQnNfSVmrjNdN9c6ECr3W0RUhV0Q
xOf8R+0gExOauj0s9baiB5RmedDmkEr/aRQBasLKzZTfnUAr4qTBMT/HYEjfY/inPPjj7ptS6/iP
hbC/ej2QGEb1gQIhHxro6oFBLk2Gi763qAzkoN/kdcPmxzgM+4k5TYmFWvtYKvPeanxVQCP/HJFL
+Gut46QTQYQvwc9XZ7NDQQnDvruNp5HPQCeZSXYLf8hq5daXP2jDnmqwQSlcPcqAfCiFEufVccJC
Jf87Bs/JfEicPvu41HhzYP488mhG+HQwFPZeZYCBRAt4nHJfV9Qbabkz1cDreHZdy91eixJ5jHH8
SQ/6LIIdfGMJUQjGK0sQMPf1nxL50C6+QlULrjufoVinwccFU2R4bzJws0GO/6mRBwN05AORhEQ+
2Q/WlxTNCRmfRNXMmoXSyJgtLFlq6UKdjr1c66fUVohbQsJ58svzxyJM6HWU13gPpshkvSvllLF3
Kl0arJ7yuuORCCa+IRvI8n28W5bCr2sF6LuXVDjWeURnqGxP+z2DiDyXnaK0f2PvXcpLnttIpuYp
1KagD+vobn8pmMCprMgwp7E/Lg//7XWrykufBl6Ezi3qVTffYQ5t2H8BdG7dBkam/Auq3KbS4nK8
yaH//ryejsFH69dxmtzqKwSXDmf6Q/7TADp1uD2pTDV9lIzpZZFpq7sAzYR6ADcE4W3X7JFRY3hM
stLMFUP8ZCC3eRtCi0jaapWx+sOjfe0iOXMkdyyd2pTcu7PXr9rh3wzRhKbBOKA7N8xOmzXM4V+c
3LsXLdWkg/LBibDZloi9CFyuxqe5/mDtaVGN+i/+Jcd8/DUZEyxCQRu7njb/v8glsL8irC9BJHAq
rADo+1vXszNEXgJyFiPqVzghtf3dy2L/FETsRAG8nq9sh7xvNIMc+03CWtHklIEreonhmRUjCwaZ
5297YtAn7k/O8czXFlhq0/tyKO9OjC7ZLXN6jmMaKfYRoV55BdwBLf41JBAdxBYzSB5K/9mGx36I
T8gIn3/OAOfhmJw3rwrHv7LYqiEKrcDjMFHG7PbgTLdyf8Rfr/7J3FFdZlKgwkknt70uvVPdYQRP
l8GiRlZI2ZP36jF2ZQzG08VhSwS80ob6Nx3kSPhostNNwXKrIQ3B8vNVnc8QFs6vtWGnqozoUbWM
KJ4TpUAQYY+X7uglyOf9hQ2YcQVixl3fw9mSb5SniFLZDRJFjsqvs0IUnfEKiINsRBTVpWJ55rzz
twAO72/uHO2xki/vPFZyCBnuuvjzhBKonlvmsRrvHfBj/ymPWuVwa1V9d+1M7fD+u1JtEHQPR4NP
fontWfMgTxOvv41BbfShu5tAymkHkW1xGwU/oNC0qDEumbqL7MX1w/xNBKtYF1i+essNzGuRO1Ge
MllH0Mclo+ZgO6l6/hP6wxdW/wD9PivfA22z4ceSoRqRATNgZHCIkDjJLp9KcCIgCIVaFZKE5hTn
7L9ZFeax5fywzanteWkQ06XEgPu1WTSfJhQiZbypFZpL6Qarvj3QNP5lzbSz1yMCLzC6AySWTQfe
OlQYNnnf+Jq8yqbaTy3TwvbhBeHV3BOux9t5G4vGPdQjWx2TutheLPEjCGzc/o/mD770RgJ9ozVE
NwMGIC8BwL9kDmKs+9zZ2CXSPO2GOPikAGJYizshTesPS2/qNfkx/16R7NdjQfzBUmC+w9h3Odgt
mBCXWa7zerTrMMOyvg3Y9HdEKdNNii0ivsaIAdimMrvPeoR1o/M0bsKnr44UjufHiyCAss/cxbLM
PhPd2OXeCYfjD8WgTFsmf3yo3k1veeudrRjOtPm9usYboIDbPRgM8/64iqxE530zf0ntCFuYd3R1
nz7jKSVA6TwBwohT7zWygUz7B6abpqh8lNNl+eYXMPJ1DnPfz1fNkyBIf1ziuutnjPxVzWzFb6nG
iZ1gVHhg/v5gOJN5t+yCkhoCXQDyfC2ZdbKQtssPi5Dz0hVTS0wcMQoPRZdJ3+0xn7DNRQJiv2GJ
x0SQQaAgJak0Nklx6k1wv2m/eyoRGBTcYICrj9UkgyDvRAcFwGhPbt9kXCAFOjP+Psv1fsBYRENQ
sNDncDt52jrEY7KAdgg8TU5Pt4JDM+HLnWP32Uj/R+eJRrgvBOTpzehOj1tdPXk54MKGzsu4enuw
R8CLF43AHkqDupauhwoHBzs5/WUjvD/kSqfZIRdUobmIHLvnJSJEQQVGY7eE7hL1IXTOVpaEfo9X
XuFZ5Li4jOuYOxgrvux3a6gYioHsoH7NSxjPyCppzXJwyisFBjmjgika5qJ5Kn4idfCH/Ap6RFGy
pu28Ed6jf4mKJEgA40HQfTzxK7o21sRynRoa+Z48Zi0W9JfGLiJ3aSC8SPIUzkcDIBrijeWO+NGh
kAVatPdX9vb5bawsFzrvnPtvUmdFl09CL6Y8xY0DEVpXnsILYlxpnoi2prUUUi7NnG3gEib9NKhP
zZ4InhgOO/BZCUYSakhzjknWWZgAkC7YRVoqMiT2MzVeK47AI0lOb02h70M5KPkuyRW1etJBjBiR
xZC0ZHMSqKsHhuOH8WLNY9yFikbxwmjhKn9g8aKq0BwzFVxQFQCexJScMgPAUhsKKFko5NUjWX/Z
FEfQgwTXLiTUhBty+Tl5iBCfUpC3EYTXS5SkKO0oE00flCEj6CKDpCSqsniW4MMxRwHBTDzYfZyd
uJ562zJKzSxuZ1goQySfRWOvoeVDpBeP108jl3M7tD7DL9U0MhD1ovJVrnwzWPyauaGBOpDpPqZE
AwiSCJ6ktA2+4KJs8r3yU6owpE/V97LQVBkV+LhsQHrugQo7SLSMBijMTYQ8520cKlcNM73POami
2IXamuyWumxzNfhSOBCC2iHmcUHoO4wYHwGqS47c5ShIYCMbb/5/D2zDHZFRugtq+UzLd9p1It6S
el9f3tHHl/W8GJ3DliqSi8MIBFEIg61r68zokZWvk2y/oK5Sx9Z/8kMPu//NCVrCXeNpSs9cWtqS
Zr/E/sJkK7ye4QIdmRb7LadlXPwh0b8Cz+/k6UOqyxMm6AhL5embbQoC09L7YkUHGXyAhEdXl17X
V2Uq7GFWBXWX4BXZXD7pB/+wEsOiX5RWEthARzAoaFlCjYkPN2SnGMELT5BtZvxMmvgazhxbNwBR
BceNuZwm8WDuG4kwAmyc2P6RA8p4zrJyODJ9bBq0iiqarNoyIrHl9m/6XL7BQ28RxbQAxkZl316g
/ZFpqlVOBSLMyJXf9VApfUmB68mQIGrk2P+q+Nem8jBO6zhaPB/CqnDOEnlL9RgICYt1Rg8cZmDK
JfSOn3jo36UQMwfbLFkWRUaXVc51iSUKVbaGu5SAerH1iua956ZA+FLnTJI6U3dxEihvvOU9FTLM
4qafmca9bt5KvxYaZHoblovr6P1tX2ia0aDy+R2isxViq3kT1ouOc6sgZKKf6+DQEC9LwrfwBWXl
IbHvd+g2mubudaaH6q4jRCAH2MnXnN2XXrcJTqmEumwjHdu7BfYPFikLn3o0Wjzof0ZVf/8aR0Lb
qcu8nlUXIzyVTyymrjZmU2335dRP5/O9euYQU6cJEUOSZV0hS2tGhgqu/52LNP7FuCnxK0BmlS3Z
44KsBYJCBiy6b7weYoiyNAQwIMNwUagQjGC/NLAs+J4RqqDYz6GnJrvG/eXrJvJRENUnI4p/gdt9
BYzpEtusp0043SZQ2neq2sZ3/cPgq4uFpXNAevy/yuxH2QbvbiSTEDLZVy2pUeKc1WeU69QafAut
4zxviK3PdnHtAvXrX3hJ3dc+b8WbXdj7C6Ibo9WUFI+Kk9vmb/sm0E0nghso89InIxIM4oC82rT1
QaE1XD52RcqTpsSGCnWd9k27Cej/CYN1X2u5dtgv6+cgAZ7BNnpdSTQGh2zQCfp7A8UjsnmBcSbs
LLeJOL8W+S4q/vpWjPfMySMlrgdu4DdgY8PFYsXd9tbCA4N+jmWkmVk0ZOg8GvqzI9OswX19xTti
e7pLGePyu7eID5mE8U6aTPM2ci8irj9hjBh7ozCe4KVkHoI2/d+njL5MKMyguZgDO2cuDbRQ0W/g
6eJFlj8mpfnvfzMgDLKjkq8V9ZVra3imhk7t4PupzV1M93oWh+FeLMZ5ieApTOblEHNrFb+5J5+Z
AXUm3gdoJwGyBO/YA8wmZqwaWaSYRTAGRp7RiJr5xzp1shuupuiOUZo+a8VOOsMFXdTTovH40zkl
dDcV4lbsQWBgbweIVqWWBNP7M33d9gSXzJxuh9ENQjSggm5EBvHX+I7ms1pTW7fenz0+udj8ZQbT
YvlagazWqHQ6F6kcgjx4A0estDfTIP+eKywBvn59WXnd6NLmOD/IcwwxRLSh/IPIWFfhNna+X4Vk
qv31L903mND/jRnUuPqklXTTrnYd7zQWT+4o0yE9WOeFedzRR6SSzld5WkSuQMysNVc4d5spnm6z
EhgGV5bJPnDHBcF8ioHPNzZss35cCA4WVZPYIY8Qx/DiK1cv0gzROVrgDcTDVzz9gwPBpmYz/Wk7
TJ3QD83cAVCt3siMBqVP+eKfO5EJF+PyJfDiuFJDmn0ZUaqxMZyDYYbD+FxGloFycrqZKUD15yvO
Hglm6vwer/eWN9wkaxwBKOAOb0XOUOtizuUpU46vpU6bweKVNldYubqRuqq6ffmj1KEAvHhJh0ZF
j41eUSTVdNs89g1yZnW9P73AGVuAtogByQXDf5md++xEFa7Qekr4uTlLPvAIMGWn2JxR5tsePqko
lj//JH+9GtcvU+mcEYzfazLf6htm2DYl9Z2koVV0q3a48FetzBtRO/kw0SXwdngd05mfQ3EOZbd3
p4pp5aj7hDfyROp798YFwAJulVfXe7EEoe+9GuoZ7uIJGrjUAa4qcmoBE3+BpHEGD6wz/+DTKkRi
VbAr61aDPVe2/mjRIYX+Y6/NhI/q4m3j8N+dvnRz7lxPr/jnw3T6WR0dlQOKvUMUF1RuXFT5OGEZ
U/AslFAqSHUMakyr5cNPwERaYoHgGwPV7G2NASHSNXLqAYZqcsO2EdEZyogOV0CZEqD7Pmd5+UXs
0z1uluSKoskGgznl6PsrKGCO1TivsxSKDQmXLDP/cVEVTJ4wz4PBIMND86gGdUqJuwSxd/7UFOXk
f3Q4t+WUC2CiDv/SuTzOcgmwHF7pJ6jVJAnI5Fe+5e4Jvq25WRH1dk+SVG/5MPcbrP77LVh3FUTw
ES2z9Bn/NEfFlsDauy4glNiJlfHQflggT/p6TKGElPB1tm4mwfUJlPZfH3JVWx3bsYgzaNy+yub/
VYTeCnAuf5CcM4xkGP8c8TXG2BMLN9nqM1RAXV23/DczQwYrI2JaTQ3vJ92aeOSBnCfGihWNiNi4
6UR8xe93sF9XNtL3c94XX3xWFZiX3FDf3nR/+k0lzmD4T807fwO48lsL5XVE5085yRzWMslQ0JVL
Ej0oAfeq4XQu5tfMAObdZ0bbZt22Zt2tAZemov70wdPGCnIRaTbexYTd/+fx0WE1tIdu/oTnhvB8
9BRK1dmGHHAnd9kQyoFzIwf1g32/auRdF3nuEMqXNvj5Mo7xPl8Z61/0T/K97eS9IU3Paic2abpQ
ELd/M8qnHwEOQeCR11IyiuW3SNLHYYjvXeKgSoZBnLi5emYL43Zjwc9+Di/PNdyWvBTkAlmYrwGl
l+RJw8zMGaXk4pibaeAOYE48AJMAINWQRk+hmctNHBzPsfnWSpiLM2UlyJHRG+5HXMo/bF/4+C81
adlMBDRPGM03aEX3Jefogj5jA+0w3WunMLRBNvxG37PRD9QKabG3Eu1fM5ARIxBNSJowKAqO55Tr
Elc6Io9WHfJ4JMlHkWsXl5stghy0QAT0blGJsgtCpYzhRAgdxp2hx84QQ/XMF09WOTS7YylvyUby
ULcuI2cGv315VYuRAKJ3ilJVfLMKWoOitf2w9VG4rcvVwSRXb4nu5PQ9enPSDbHOqUgJoA8qv+sV
7WbmY1DOZk4o4T4fRATBrHqD8K5/dLbAXGi4q6gIj4hKLsfUVCt2i8Gm3g1ZW4bvKlvChwxdtIUB
jUv/X+fIaSlbPBX+mMzHzrUARgFYwK9jxhUpEk+vziuF5VuNk3WqH2axD970UBrtHwwt7ZVgtC5+
suhhslCWfWI+FYpH/85eeEN+H/zZbXHTq60B5mSq9k8efrhaDu+an8qeA5hnLkq2/v4JpfurlXCd
H+EQIZEKWTE6vRH4f0bEnU7rIQgJl59W456TlnUwQIp8g/DuTpNXEKrftjEeIYLy+SuOF8ynXbwP
nhZ94v4mjnATeDJkaCtpwv7Rk+15MJsUWkpvzXvGbjFH/COSCl4dL2kyJTrpqEmBAHU0wQ2rcX1t
BoRsSHRDhZwiqMkaa6dq+yY1RsNXt8p8DA+jbJM6R4IIpVIWU1SXcPlMbAEK1Ct6zE5KF4Hp8ckY
PHDw483Eq6OS5E0FErLnioZmvZtNqSBgIgH8If/qi3Tro5MENOEphmWG1O0wRb6kVfNhNzurrWBC
4WZMmdFZGpRRi17h+PMYAvbFeQ7DyHorx7SLM360uRWCh/pNfvteiHUX3dzrQ7qelWOc1a1JO9p3
9dDNwaAtyHQa0wUpEOoWD7cJEE8aJv3/mi0Rwi/Fk7ad4Y+kJoRTyuNm+NzEoVlO0Eh9wlc9icHQ
2sL91KOxmEjKD4IBz4Z62qEo7C8h/Zyn03YAgRxn75ySlhlfr/i6FBITBDE3BDKn6lF/AuXdmDi1
6KJGMLHywItzAOuF0bOohoOJ3FjD8+U2gjbhSCWHn8VgpnG4tz7mS8nmoHKW+l5nzNVcmnjta99k
d+tUEc82XpiPu4GhsRwGJ7Gh2DpHC8CMFM9zxVW9Su9EPmVl9VrrdBWqUmPEGDFeYwEhF4nUGTto
7fm7OJIF/8f3myeMfw==
`protect end_protected

