

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cn+MKgScMmuOXqDja4nBGV7WBeIF/ysF292lfgaKjpujK0iaFYzIB0eXWu1mkHfQiveaObVLOLk8
mrHpA4NCow==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lyXUbl1fNyCoynCsgKvsnxh4xSVW7h/6+WXSvHl9VdQRm1K5kCFQ2kx6cA9GQA5tjQws4LhzjH4C
jiN86wKYjDRH3aO0ipukeid3+Cl3Hf42WJLldVcK13r9M8WvFiA8f+TpNioyqUM09aStqFjdSjjo
csyM4N1L6gYZVbIwZOI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ocYp5Q+x2567q86I1MGJbRTpHjo6XgxppbNT9mGuUHy62i1N8b9FapDfB/As1HxRsllExonP6L4i
nOrPFX5dqrfhgwJzsoiJa+kQoi2nYY4KOnCB/Pv3Scs3TRpf2vM9w+ucmXI+o3jD4h7K+rgsIuZr
FCyudD/onJvsmis4CLUUX001F3EFidOEU1Q030HzWCJJNPr3CSJCNNoHPiRhh83y8YSpsqXjqNTb
qItJOecjL9k1mrcywbi+GE7p8H60wh9osKYdQVQMrETxJObRc2pckA7TWFtDMJerirE3KnEZvIsf
rkobt3565did5AenTYngu53T6wdatItFn3vIuA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vOCsY/SF8gPSqD/ldVKm/v7jmfpM33R1VJXD0UiCtFFOs1P7Tf2U4nhuNP3HANg0qD2YjaGQ6myv
dlR6lzeuHoYmZN/DUwZJGSaiuM1h6qmcn8qFSCISMqaoZHDjixJ9JrSXtSwMaPXqwy3RINyRZxZZ
n+tFIFvhOGXInTnHa+V/8xfZhzHNthwln8CBoCm3vnx5oPwRDkJfP3YwEDF4x4X447JPTEXORFnC
I+t/Qm3ldihxuP2e3EP3csValIaPqAY2BoE1dXhtaXAVGywLawKNeUCq9IIPVqj+KxyFneku6GTO
rnMbpLS30BN7Hk0gd76CeIpd158Kv0d8sEsmpA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dhHD5W3lGGtC4CZjL3T8nBhCONi7O+vACUFgJCKoGDg4NGC33+yxWhu78fODvPCS2DpLrPJfk3bA
djnpMpnwkBjzsk3CeFcPREHpRWWK8maEH4z7l4cbfw7kGO1b7+ekrWpBI7kV7eYckr9C0k8Ompl7
lKzWRDsnDke7Jkm2xJPdMkOOACVdIUAXKGvSGFbWAwk5E8Rp1UFWwqjmBhVrZ9mRxRT8Yg3dtQPF
q0TNwwUnijSFIcDGKDKuZ7CNTFcQuy/Tc8KslLW8lYYLxncygRHOjdaP0ohBUBQua3Io4qpRdfaV
InvJO9Dh+lNQuqdcaJvi0JXgF5GixjCSKmKlqA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Pz0913pmzb82uZOhWjEa23X64ev5vHsic1WjUUDytBBbAx/E1XSrB4wbUFgywP/okDl6EBGDGRvX
hoS0WBJe40mrnz7XPUgtp2OmS/NgcqGE7AhEty25v+Jxpgtk9CS4If7npTe95nuyFzYHVToQP4KB
6/HKuWIfxwjB8zuKPC4=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I2mjOeLUUoNbFKbqo1sWmTLCRf6eOvt7iqKURENUw3Qh1TB1B+bnN/F2rG994bfIQZsB5fvWkgKN
FG6KCYNjKLRpH6Z5OVJR6fOANjgDmnm49QXLpsNS4efTdEf+OXCcVzbqTKCiqtvuRScAI/nsT87x
y3rpJipze8j6Nlb8T4cSSjZaNmboEH9yPf7AxUPuY/HaH+yXbGP7PNWIOYU9iBJ+xgANh+c8Rbay
KHHeEYhxcnp20ptitbVw1sh77xQpfQIoY0Bv7zFymqzyeXKX7gS+ski/Y7A9b9aGTleTt87NJDz4
ncJx8n/LI8MaThS/7y2WYyDJ5UJrv2MXzJNvJw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
bxuslj2tr+jRPZMN7veIdYwDdDIVBd/k2b1tsYzRjILkm9zIxRMVZZeIljB7mzzHsw92OYobn3Fk
ihAJInqsxmMudtDWLEkZ0Aw0wQuDKXAT8NtShLNk1AGV2oZ/I5b4nEnrV2TGSxClo5Cr23QImnQD
YWdI/FdvZ3whEXB0NLv+LfiOOABzcouF8z12DGcKM8vIYDHpeZNAWecFxOwSlXMi4B/cPKH+BEQG
wvkHWUjoodsgSH7uFZFTArNwapgNYZ8hq8ZYTqjt9aYbL4Ez51SfinO46to2oUsuhMqddCyLFybU
UDTI7OJVknqjWFQfbW6/KWBfk3ADJ0svNfq4yfOop7RvqkDrFmJdvpRMhmp6faA6krq5YwTkqT7Q
8THgcFd6yNQdrJkIKjGqwOsZ4r+uyyDuuz2CXd8+KaahwuSxt5XSI6GSRPomc1HjI84wvgMupYg1
sPGJi/pEz+ZXJ6FklTzONe1yePBouqSMjfoPq6qvZpaH4oG12i/Bw6QxHzivuJ4rxDuGLmOoNf2o
PImlRMHOFrQ+Vek2mTR/6cjLHW4vLOBj00GLNs2qYYHXTjrP80l5BAF7B+PrIhJarGkEKRdmXRT5
wIA96ecZPt2Y1elLleZCWMFZQUEXhvJMC7RIrAmAdHIYEGXfa9pRk4iQYZPXdHV4uHaJRGeuFQAY
A+/5Cqw1d6yDRwzeOjclVr15mRTwnK4eoi9NNEiEhvnvh0HvHpzv8m+8lHR1uUcInSqFnaQuzcgZ
1MQzQDXAkNuzpSGzRXDDKXEzN+CfwYJrIC+sGRRilyV8nbzieWi/j+TT123+W7TSuVc+TLlaKoGm
eKesUIlQeYDKN4p9DbEYKNdDkO4nBKcrNsv0gLLO3nBkBVuZxm23qASZfAEGMqeZS6DRs0tA942v
tuh89wjeAdDPaLU7+b2gAix9PcIi2MkxeRUAusjQF6EmKSeUPHL6G55enuD3TVmCEZLCat+wkzRb
DIUBRs2F6H+DtFxQo7d++vILyfdSNeoeuv8y+6urEjI50CfPcycrrOE02hevAQkVnvJCRFlaBwk5
9/+4eNaufxf94ePpPMOrZkw5Rjb+5PA274gv17kLOm57GpUA+xgaVj5au/QCzUO6QS0ZiDCvHUE7
6VR61gcy6CFlUbQBT2T4hcTnGciw7y1I4aD6/jLjl0TgDyl21grSAVFWWqBNOfNV+qBJ2fNA3Ac2
GGyvDJgW1/+wfgRupK1FOJV+7bdt65c29cYTr0yRqMtzGOnOPDwbLzxR9Yzk99k/w3QjeiwVsgmZ
IBtoXJkg8ry5cxQT1ivN8yaSUJbsT+OvR6hpCtjtNSJyQr/akcDBFHNPkDBpcX80qKXVVnt9AMgl
RVZMNk4cLpzXwdciIUXmJxmznb6WLBQirtK21daZdv4NvIukGmg8C/amJ+8LkHfK3F1h3sR5eblL
MRsm6AgsUEmV/bOoqX642auAmyZ0BHJ9uZDyGxNMDPXjwEATt4rI1Vp5BkyvfFRxnOyuMNiLUUsO
UI5C4sDKq8UjyFqccspTcKBsDdqlwhSvv80LTPrX2HIzGXh1gnXNI4MqlDKkzzLUfjMPLyiak5WL
78zkvoHoqYFm22aC4FCgovq7hJROuiN7d44MVcchvN2IOdiLoYGP+42g7cnHtipRJ5jb/XT6zRSp
tSQTkQYdB4GKkkg9FQfY7kPbUkDrCkTY5BKr6fMHjizfEn2nZI3Aah5AjvXj6M+F0CjFEcNfa4Q2
cc8PxXJSoHGNHBT7M84uKAEoYYpkE2s5FYTuTB3uSnUkSFZoMT23cBT6rRmGafQyhfoR3CtKZ51F
kz2T9dV28g4u3woTn6v9IeiFHH2eNgZAJzw7Kj7iGuDQyC4/p6UDX9ZvePT6Rt7WS0og6tSPOt3/
8KwbDjVkRV9zW2csx5sJdz5sv2/Dzq12aiOaESXfGsT+hNQBftInnQrvRxNuQOFxpE27AZxZ9Hw3
JdryWQHdvSXWZD/l1KrViElfzUJsC5sAf+9WxeQMQBbBX6tGyReYLM8vEn/gqK/sogtJvHdTx5j2
jnP7Hb9/YRJggQ6HG8HI1Zu1pWMzlggSltr2G19RF1X90Ld7DR1aTuWBxKHrDSwK316w1PWMvR/j
EuvZCAXH849acdTjDGjfrYW2FokMWwhTUQFyKawjgrr0VVitFeQ3+hqm3v4YQa7y6E2pyrVTKjqd
9Ez0pQ1ApdJzPzuR/LEg1Bv6g2+twyPZqtClNiM3/QJwmd6XmOsc2SfN4ebPzlP8xwBN7548WeVG
3tAUxrXRbIGDT6L4YipidsqE9RbiX0YrVxEdkXfXWNmd735zpiJWMdc3IPWNyZItWoKwmRPmqn5p
cVyW9YR/vsJGhiiaBpd1MEx+U5yGNwXxMWgUSzN1KoO8Eni1zCtEjSBXJzYTdqZFYNROHUXxaRCH
bW3BH8jPMUxa7i96Dod6MjQleWG8BPd/2LZoyKcUhTwS3mL/jpPbbDyWi+ZjO/+JpNmPH2yb35cH
WIp6oSKG4gr8mWLblOVLpNI/VpC42E1SVf7KWFtozejotmm3/s0I5L4EhIWrzPn9wyyAw4qoxbbf
i0YlC1L14LW6qTguwynxaZtWa0qjYPYe4K17CfOMOeiLyLTF6QOrp0gGTvIzLIxLjmYgeCAqpEwY
y70rplEpP7AikteCImsJ0Xa1CYPcyTZCsMETnZmzasHz4O//zlyqJ77wCYXgPxyd4+vpWgbpbfcV
ThB2GldRWlndXSbQlUaKz7edrgF1HefjM+3jne97DLjOK6WtKsgfEaPs7ANPdOViV8pZ3+vxz2bF
XFsZA9wJSA2hRRxBoeKxZImXU6BpXGf4GJ8HK8cY8sIqQ8OGpSYCe2GxnVpuBt3dNOcBEcKnPWer
7GBLuURiJHWvqUrPgDHF53ykX8CTtjR02THmES84hCwzx7JnU0KAb+XD3nV6uu9K6XzKrQaPclpl
6LOjmtSZfQUUhJV8UyvRXdNwlkJlHmYjm3fmm3I773emeN/ldHGD9d/nIk7adXIgljExHtion3li
VPHwd5XHEaxe3+Lrc0E67lbyPJSuwLXciQCNQQ9UpHr78qhr974dc2yRKfjC+k0E4MCnre475PA1
/ymziSxACW/X/5kqvmwxYU/bOyblFUqCvDtnFZayUj7kJqpFoKH4ghJY6VFLDPjJ49YmEZ31dMEB
+QJ8QuVPRVJ2b9u8cx/4dRdKowuaLZNC2pRC7wJXR4tF5/eYEu3fS2eF5bk31Hk9vxIXovNwCrqi
mqKNXtM346ZoKyE16pje2LOGhW3sJV66d8WafWZSSA8th7/v9a/eAd7igdlDIWFaaOwFnXvc70F+
NNLaDEM854YQVn07XEgtnIxpGy9uEN9uqc2cDmPEZdtNqVlGzuB7ZvhHqGqCRXrpUAn2PLq1o/Js
IZe4/GcRCUfox5WJGUGfGpiIhx9HoF368TOY8HOd6vrx3lmrKYNbQjWvSP9XaBYVTp6mYg2SGTt5
1J5Cg1GuyoF3/f+dt6GIGqrJuPM4MP1TXXksN+q/0AWj/LVp0nTH78mzlV2WGY2j/MX3duSU9str
Wiz00bmaGn7RnuReh1s8/MrpEoeRzWiTS2EkLLlEgEXncEKDXAeO/W8PYdFw6XM76oixFQUwKc97
SGvCJJwuZ0ZxYafEuxx1fKAAKsPI5el5adQyQQwUFMM6LfZv47RNHMrE2j/EJkR+U0aezUbE0eMl
B5KpYrpZ1zwNlrCip20xFRUy2kJTXhSYlEmIi5bEGT6eVpe3VpigHIBHMT/nICvVV2h1i8wxsDYl
KrqiOcfnJNdCt8ht1LS+Pre1r7b6bMw4IVSwe8YUw3aHAyKQOvRYc30mSchJLNik8+Q0zqq3NSpr
LWym/FxTS6hltC+XZDdnz0+zFClwYh/pjnx03oDy84x1BVddm+nyYJjwiIYgrq+2yYcUSEB8OTt0
y09zvdrW94yb5mMnTUoMDtr33OvlFZRorqlJzVLrh9ctE7KXzBeP9clm/PSskGH88cI1KTERxFox
qdGo+R8S0PD+4zbBii8B9JJgpMNnhphCw91wLZ4bQPxC3i7dzjqyYA1JEy9gSLPZYfGYutV5981s
orzcimrQf69PgT9F4WZQxv4CgFECmXOLzcqSUL9q/KFmXSMZDWvH8a2j1BEiQHmlNHJ46MyjsriK
93+ELZP2IjoejyFw0ufnmETT7I6uu+lsGHZkkyj9lueg7Zf86DLKKD1nSB+hnXHuQVfJu8ISXyiz
bUkOmDo1buhQBGYdLhE0+5eEL3DyFGVaYeanpckSmXilecoSzpnW/1KUiD1HfC+YaLXA5LJWFuBS
82xunpe0PzpsCu5IHvslTCbmjlo9bsTFfN8/Gb5dpBcikVY7Ia12SmjTQK7gWM6zkmvkGCJUmPRv
aO7/5Fif6JnReYcJ4x/HPasTRyRFetvNK9NAQVWRyh9YyrLdvBKqiVTIPApw/4McX3N71MieTQ9S
d5QVb7qiqQucCVTmhfD+oP935f8L/l4ueCQj7OCcTwbJ5ZLJ/HGdYqMr0cSFpUBYu7LhN9ozQKld
jeKG2VuMw76TQRjzMUfMb5c0WOqZ39ZHFAiN93T0FH+6XYY+hpGeJ0M0R619fYcNaX/unacx3Yul
LkzzcGV5W8jCG2pTYyw3TjftL9ec0FSv2gCCNTaRoUswE4ziSNbKKuMq80sDGigJpZphPljR69WP
ADdEXCZ9FTKPqSlswU5lAca1m/mHr58GM86JjrI6+CKmlcbTNyL3tWbx7J2VfWlJgrJeolklcbQU
xfukjfnLpR0natlPkvPigVisnWk+e+1WRA9Jret5KJvo9ZI1YivWA2nO+3xOVvK+ZJ+Hq4rJD/hR
/+P7mwP+qHKnwYO0/who94YQJ7KrNaquhbi0VfkPWcgN9EMsd0k9KBJDW4euk8yYQuRCN9kctmao
MadltfBoGhplXCQgYdmhLDVP1ug2XZgL8HRYYuLPrUKh2mjYzLd4nhCSJ1PNVEBTabsFHhG3/oyO
voEm0oS6dUHSDqiaeJkQD9BOtSSMhqH734wU+04tfjENCqo24XRPdmEMNEGceCmVdYqC9l1VSK+f
CQBTS9JvxQi3FFR96r+HN4bD42yme9lpzVn+38pa/aKofrS/JEdZmXVZBhy9jVtvzvCctS9qhSvl
DXtjEtRTjV55MndQSQp9kI/0K0d1FLh9CBLsIl1oRhkCmUAG12GErvmkIIUfLgFmKNB5gWP4Am+a
y3NIOyhTVl2ChPgs4p+SNqVcsBFeIpRLMh8mb168zZciC47+3mcacuKTHaJQ+zi5O+V8sArZLQNT
qRF/613NMaRMvATBvp4x8Z44tWi3iUpJfTgciEx+6ngwu70u8egmvQaYn+/g2+ndSQPVYOfer+Xz
cVWeX4gLyqGPaAb1KUcLo1Wppg4Ovwmnty+V6ONRohOA7DnciKCGE//VKRxDKiWHQ1kYD/FZMRiA
6zobwGlIlu7A/fZUGecg/5K/w1qDoGQi4fzas2pO133IUhsTcUDndzmKnTjPJPh4aA1zRp8vVSKJ
kLTNLqx+HyTkIWLoCpm27I8koTduBMjUIadWb1keWdwO0pPLxHdNS0MIGFjBacFd+1msnDqE33ma
gPZHTIBL+GMjjr0TyvlA/3tsp2H1udrlD4+talBaYRRJgfrGlVLFQy3ZtxVmNM8rLGrCFJNNYbeJ
lniS2HrdKAVQWR9wrSzY7yg/orCYkE2dm7046j7SoS4/eCscOkGu0KAj39QBQnidtHkf2PtW2gui
j3d4/n1QHGW1vR/dvQgBal0ei4hyaEvqZxtf03rKqWMdDJeWCaVA/kSXm9Nq5e0LizcekaL3kGaR
/0TP7ObtRlIlwxTGMJGY1V6BMrB/vaizghx7QltC4FXimx6K1xtMs+I1hpdR020sUQQP5cxFebJN
NhcTZ/mah8CTrCQIc8DVYcue5mS17RqSLjivU7pWc9A6v7l6c41srV7iKWr/qwbWvsF/wDui832m
iF7oZW0Ur/VatrjCx73Q/h8aT79M8LROwe30L6JZYyOPFw+RxQWsLT/4q4BEtnmRK9XZ1B+3mcLs
+f3fKgL7+KuyGY9pkoqPhAv62eD1Zr9N/J/80jfmwGfS1npJO+EJzRQ/gdRgMmyy/gxuIwi5WVk7
8IvwssnxyMuMnlU2CDv/je5Efz7MvjF39623rSepkpY732vl2qLAzgbYqoDVtk/UiSUriQFfgzla
7kPlfllkHoOtM7NGER2SgjxmQ8OJ2dZ50Sjhn/I1tev9Zcc0lgQKo9KBuKTaKCMxscTJw7MAcL9r
Sb7xYQ/ZJbQpq23Hw1GxXhgKJ0dZFVs8zcpCO3mNEEfQ9ciQ6A8mTI8Mzc3OU8fbavzfVQqMbqoh
Eq1qKTSDaCCfsbXEFp/JxAJfpVLv3CVdY8uu3jz1N5o7Qb0JFO7faVZ03AE9sZPHCSHxxNqmGhU8
DsoXkEmewdZSNDvTVgHmNcz2bT4tfwdq0k6FS6K6RWBlsPFPKiyq4X+dy3woCcKXwsCpwA5tUJFs
/HM9RSBR9GGDH8HkZ0OiuQhLOVtM69Dxx3XZHxdol0U8vQrs1rxC6fwyRbc/aB71kEfM/X6vmmH4
xOGFmFPhJ4qp96bqsvHPTRr+XJWZ/46Pz20UOb24E0VW0vLMgL2BqDJbq9JKtdEOAUE2cOVdjQSA
Wmn/A9RXOUwsLfgSiE2KWj0rU7rJY5pv4EpCZNZZErSETAR7reerRTIZ3FguOQhdbj5BpNOfaxQs
p5jgAHBvI4wNHPipgEPacOESHi/1M7ZCG8Acnhayc+8xuCPA+8ajUxbfuhFWKhpznFSFPj5mB+b/
LpN8j8XGhXedjXtgJnTJJa9ANpu0ddrJOuJBcImFypWyWBxEb3BP2sDibbPsERcN5frdMm7QfAAP
a39y9sZxFLVLYFTqQxMcurKT6Dymrl5D91dXvFZy9zcA2b+SasHunThjxuGAOtUmn2tE/EQnBMl7
YAeuuT+BPLPB8ED46FTPpl0ZRmOha/O+mfeXLDAb7QLTuB5elLlJ2T/k6nbiwEp2O215Hq1X7e7H
Sl7rlACzre5sYAYd4xBjb64gaSfYm21bFUB1dB1DDH3+32QEI8yQyfPh5S68m6l55PS0soAwCWi2
F1s6uMQaKw460AVEOGTnybFY+F9gYECmafs/B0gI8+MlUV7e/EqXRnkL3XKiBVz4+AKWdL3uRFXQ
TLuqvr2pPCkGxoE6Av8isaf3KJO/yD40IaEr0VUiOjuRrtjEU9UYW9ghBsGLKt6CbNzut1x/QFWS
igt7AAjJzQt2QrmPk33tM2ce7jEf5ya7VisOaivrSxBgX68MbGJE8y9saFJtKCXQqoNyk/zIiVyY
800szmKYEx4Do/aqBBdpu8cdH3uI4euZoJo3qMlPssXqoMi0qrDvIFRd/dYi+2M5RlWZOaRGXiFC
oO9ZOXUel2vcSl9d9fy7lmw7NwDpNkqnAy6oXYe8yi2FusI3ma9/HC8GPP9GFusn/Smb7ozhEGge
85FKppdHx74LetpE5c5XRE/i0Vj5Tqx+fpylynnrGpa3PaY7kghCW/gP9mksn0At+EY64/vHPJZV
piflc/H9HAEHber7folq6Nu0xQipLKcf3uS5tZqRwg+d9CmmYDTsFhTK8IGJcozbe6VTiy1Jl+I0
aw1e006FDgEeg2n56+xB/eR5ilIc86cOEKhEWYesX1WG0jj6eHrV3ncU93L7NUNMICFGCrqsp8mb
rK46cjtvYEtsV6ZS0J0eq35NN46clyg61BtqranMY+e50Yr1j37ATph7yGySh5JkRzE+gYiqS1a4
vG6utZgDBY7yS5AKc9JalxrPzXzpcH3ZH3LM1+un3RMzkYLyXFfVRuP5NBLw+yKs7uaV2bMMusmM
kHGK3y1CnFGAi+20xH+Uzc/7HH9hJaR2IoE4LaKo3gzu5EMF672mOsG1AfsBGOwCLJxF/v50pZo0
X39I14pgrtJC3rZ0IN7fWPtMlF71Mj3F87II69n2kd3Z+a1VQOOtfYjV6jL3Bm7ZXJbhd8iBFEsO
vRH8qkq3LqwLgISb6oWY3QClv5QdXQoynZpaso7yOKr1MMomhkNko0ocLQvXvqzr4pXwIQvfRBp6
nl//NP8mB6ck6kN2SwxU/1/rkUuwlLODE6pwBL6bWZwwG8jArggumHbBhpIKgVwPCe1IXo0k/8mw
uXJ+3QgbTor47HwbM+xQ05pYpjR8K04QF8INtB+n4yLM9R/TjDMT2W8ne0o3riSxpsArQJ04Pt3d
UxJLGL6yl/FhB04G6F+J4XjYivwyeaa2DJjuP/BKGjGR3/bXkbXskbU7N73qT+r7tQBHuOQ72BNM
2VCCLF6wjyVHf/57ntFgzmSsgXRzXxU8MB3NFOOhaQ7Jfek6xBQauW2Yei5CPV097nrtWk8N2TD+
WwBbqwZHroRAtpEyPtaoThbOd8vh6v9WcZwhZeFxr9tdYJuisfXzv7iviN0tvwwGkmvfya/YMCQ9
Gc/RfhKXw/zncrwSwh61TG3qW+1Qv6W5ycZQWhYw0wZADSiK6ufaOdUyWBA9YGoIOhIzwE8lTGJt
UbLX0y2SSWgUMAjTmFlPAVYLf4Mgn8OzI3NPDmYK+e1tVvgiIRrsIhq5dmeP9pKNiT67sdaWx9CE
A04OR74qxbU9MPXfFZ+cnfD4GfOmdzyjMOsL42xlvCz5A/98i/dgrJYMTjrHtwzIYDrSQNxPLmDC
iLjCYDQM1FopPwHMTvpsxsFwBToMW0fqw2y2eOErmmbprPwq1acihhlIV6d8Hko9hcd3BaE3L1O+
uZ5+Id7TNBAkCV9JGQRm2/ZGc4PM8+/GxUprhiZ99FtXZTEjgBTj63zJMaR8ueiUFIALbnroCBpK
0nGtw9wGhfjnHd7gRW08bDgBNbMTX7BOxmcwpo0mT/FYQ651vAU0bM31mXixmuUFI15y6SeXy4qg
ev65WQmS6JkAhfbvWWaWlx18wKXmbVcnbuwN85+8eRvBZtgeltACAK3YeDOlgQjdmg6NlUTo70My
z5joXr1zpYp4VKgs3bnBINxRhxJgNksnE1IZZbOXGbFmB745FLGbiagL5blAoLcvrLOCsGaA+USW
kj+jjXkaYDyykCerGfXXKN++ui4+c1m62QfuEH6v9X4C9DYJNXs0Tuj8fJAiUXYGRAQaPzm1B366
0plbqVv8IbbtzAMbS32OJ4MWNiDHSvzVw4HyZrGXJzKe6Dw37o885PVjByVDgd+G2e9xBiwF/ldR
sxHDdE9KW6n2qOAn7wlVCkB7w91Yo0Qjyy1xBMDwqXlkTN09tGLQMwo0iHke65TllWN6Xd4fxaHz
zIRzb6mdBmE6yhCd/5HKGtDG3LtYUhr0qaI4RBASTFVVpvxGUDzE4Gwuaz10Bjjb60ng0AgJxM5h
1dhbCLQjIsylWESNtXnwQioXweBb7Hk2S6aRCK85M1EWkcOoaglYHPwQNAjaGUJOHUDQB1mxmIgc
9eKkukYoDXYDjjOwBmWf9dco0vcksDa9eepJhuqhwNotLbByitvlQp7Jxt1xD5HwhXRS1tX/z+W2
Ahkt7g3Kqt46Fhm/Upz3WkQmJk18npeJzu0XE+qX3qYf3XifGENEhp1MoCjyGKg2gf8wBenV8s5c
JX6dD/vHdcEIhpD7wD2E4CAA79p1totYgtoZY71wbZC5zBw+4O1ANazDoAXQ7S+uw3SFuMPkcJLw
KMzfSbVuqE9/oae+mn5vCggDqMvQPlIV/rYvN75qY2ZbixLwx1VnKZdX4sDnfvQ+ViiBqvrl8RHt
80NMhHRUXh5/m+Ock000f3S4+qjf2twxh+kKhwO1RLNjZaPzzjwuhjhek7iOaOR/cMwblkwgbm1G
Q5N/mdfKslwaNuaBjEXnPfUi6xYD4Rgm28ZZ0oehLZfEpOrSPIP2uOeE3SLkQeVk2W/tAVdoN2Rf
RYFjo3CXKJUZvM6jf1/91N1LKXC8MJx7g0jZQtFPnKZlYGjiQQvfOe8VZhtLBTdPh7XtgCh3ze3t
jL2i+76DI0Q63fY/+0MvLXMyZ30wmgwdVghNocjtBIcYna2ouaDRvHTguFaDX3OghybeFkEmLOLD
kWySwuNGYj2euR7pYKK7w2V31SyMWfDyNyFR/uq7Ce2ZlzUc1wC+l8aVKvCvKIqaI5tKDKQlSE+k
CRGWuiWIcFnzhrvpcUzCc46+/d7D2msGPSXRHgSgE5ykHXmPj5WgnI8g8jXz+wveci0fjwe5m5Pw
WHfcYLSBhNNUGbdMJAvCpDfoAdfU6O/q9nvWSB3bGj9ULYjVyKpp6fO1gJ9LtWU4e8Yme6m5c9t2
YJYwcrWEq/fKE4EPtnLjQ4q41NvFFA0zvuC2usEX6drXWwBf894vHfeWC5sttTfwwotiQkTGYOBW
igDRy12Uz96fh4NU/tMbYjfIdAg9EU1VBSL/ZGDx2adeCB5Nc3P3d2W0+2Gth957DIIbukFBoQ3D
qedMhMdDuxNq0kezI2gKaJblnRByXXHmkJl75kP1J5hKEfbXe38fRaLjKa//+kwSqPRzgkm3eUCN
Spl0G55JMbrosszrChiqgLYxq6At32FTvd0BsSjV1qxz5HYmjCqqBh/iZeeQqGzk/EJ6a+CfK9Vt
swLgduJN0zV6FvprujYTaBtRkprmdc1E4jgjwaLw7P/INL1cZb50Rz2IUhDIa0Ts/hiWQhxpKO9W
rvxTQulGKq7AoHVsqoxkTFR/sXToyQO50nx9GqmvWzN1qjv+qmTJnrOHRCzXKjpyNSiwQN97/WI4
/cubYse/WsIuxu234W4rm02WzWCUfDzolkzBk8JcYSdjqN1nmrrDM4iDcgIignSiZKPM2gWkljGi
KYYXlpZO7akjcI8h7AoMVWS+0qjgOxVNUYEoriI1KRONyjxkWz/E5D/t0JgF5sN3ohqn61rhqTmW
9aQXxN3tVRGgst5ZnSdnWd3VPF4x1dpJWBZ2PJETxMYhaXtLi/V12sc2bBN5iRTgAzd2zlNVqc31
NSm+K6a5HFVpopAd6nmzPQ/O8+YXUOpqF8R/1s3uBi3c2AOB/zJ8zv1xZt0rWj+ohd63UNj6TTiT
aETKEEAChsGg08Ck3fWXCuwWwzUWVLMr8ICPphX15fMw38g0KskBEDPzZE0pjkt1KoPd4F2NJd0T
haBEdR6E5zN9OGyqNVlcujSSPYyoQIWRH0nvMu7k3bYZR6R6K0LTu6v/iHUJj9u6tpPwRqDse/1n
c8tFW+j8uBG0PTPO1TEOJ+idRTlczaUayCgKQCHQ8s6ihVgVR3FNXYgkb/UcIbYmb6IyWKLeYCJO
nIoN6gq3D5ZBsQnpUKmPlAIJiFVCs2o7FGNwOHtgqkWVJ+EV9AwRxsg7PQYznRwQW1PwJipc0OTT
/Ks80WYXhjEO/sbux+TQdc/2DZUxdVcey0y+Ywwa326YHAtoL0xdOYpLG3HTwoicnDMPzF9wtHD9
9+ZOS7T8L2MW5/BU6oK85wQNwxICvZP5LReBOJ6LcABpeeVKyoPg0jr8f5vlrZrYhia3bfCfLLHU
y9C9LOqzW2K1dnQOpbiIZ/Ky2zER2zBBoSqK9dfPSnU3uok4H6HfEMbc5gHPmQ6lw24PsDQCUlZ7
bsg0xpXUtkuqdXCeEitIjXv4Dycbppzd3UQq0K/LEmXT1fSMgbZ1WpxCRvs2KKn1YGw0Co28lauF
84vrofWlPahQTGDM7OmAYTRBWaufV7IXvydwXLFp7mlgXgcly1nBUuSmHjw9rK8aQljIxEivYc1a
ltKsopJNSk8Ok2TyMqEldR7NbwB0f8cQ/jGcGzB/XISWR2RQqwiGbeUn+6HdOfDvvqswpTgWJkvP
uQ0exxpu5PQuOOEocp+uUXG2ie346gKvV3LwXqvVpfTeChVWPtzQYtNB4q/YsDclbsrq5+bMIqv1
6LJA5uTwus85eMAw6xcTSsE2TIiKUYvFZi/IzaviSIpK30/ZWgGgfW1Sh5eVray/WPCwRy9ZZLuU
4Ak9IBK0wOfI89YGcMuxTaH8iyUgv3yQ5Nb5kc7bJRU1SuqyNRs/u77qcLuGBjnL3b3PKvbond71
PgNtFuCr+/POF1VHt6m/V3UbCWEW+bPAmisymPHRYSbkk80aMEPpTOYfJliWQiKuffLTCLitFta2
mv+/v2X0bzCXTkUGRipBdtuYS44mvBRtbneg6ZzkEmmbOQB7hMalJOO0otrNOB9sKK2h2b5/ypPf
OPCK6cRPQH2wNj64poYaOAw7zyEMsDSyTrqX3aXPpMkCGyCHTyLabGrrX18T3P6LYSEIO238Dxvt
3X2NY0s53WxLrpyRoQnwbYMeaAsX4o+E2AOBvMbo3lEnyMRoIOwAZyZLD1qBINsaG4zoP0ZMRnQj
YLMk7Xt+ammIV+er6ixbs8I0Xk/JsbI5uAULV7aBbSCUiLU9wf/ofzwOIAhnT2zziiiS99qld4e1
ZQSB5GSOdlK3UEIJww3rO6zE2wunbPefVBpJDLeqHsFj4gi0G3zC08i5SgLMy/hUki7Yl8Zhi69b
EmFJapiorVerhHxMEq2WqmAf29WKzjYvJGJ0L78ReOcWscKsLYy3JgGiSHEyf7xlC/fvPr45LHJ4
1dBLi6WSi11gLdMNcowGt8NoUgMXNP14UO4Jo4PVwk0xOLHBDCpjZ9ETOJ0v77QTin+e0yRbxDCg
Ov4Df04O+XDgetgmU1Jlp5ftH4gbG+rAccJjS5acluhyUhxV0ZHH0RR8te5Xk1KvplfgETwdud6Q
nfq+EQnzGOdxmmRAbJ3VG7WU2XfaRMIv8KgBz99UsoNUtr5eHWl632/U8XhYQxlhZlEwFjRHSpm6
FOITsoes95xmKENLcEj/VTtNcFIzKys1vrUIUVoIW0MkI/u1PbqPkEvr/3fJZ/qN1os+jhbBkukI
cAugaSmoeBBorGvnis7jM0MtodSvznsA5P+wO7PWoG7iA6vimRPAJthsTkghPaMMo1+5GXrwNdqd
AguuO1O5TuEEk03ljGtZHRrtdZtptlOrmusNvvK+E56XbQVHgxev7VbjSFUVwzJHPpOVSTI2nJmm
MemKqTGgBZPm1ruArhrDwOqunSjxDrQsXSj44GjluJlFtn/RKhXjNidZ38yQEsFeQx9ws65FAvtf
alHpbl0yT8oMpyteVCXtH+zknCHj6mqGWmHih+LePpR6hdK9IVyuxO1bywx54hjgdne46VE/P4Oc
whXCVI6MJcYQNesn2gx5uD71fpIzl00vusXlR1ZvjsOSOzAIBwlCorWBo+NTyu6zIsZcUMVgTBHA
PLx5n7ZPvFvoS8DdCDUNGQyT1jbMypHKNyvIt7YMQF9nE7fpw2gxEI/Ee5a2e14Md0QsH6c+HVWX
EV7eSI2bFbK2nymy84dMLxrqAzUbcW7qFRAoXcuFUks89dUoV1B9qLqGj3wGp9HirS+c3+djyCFs
ga/ybiHsdza90WSGyeCVmp4zqKypAVQoyRrzNJO3wsRflqsuVj5rhFHEMkevr8uPi5Lk8fp79Ijv
4HbjBF6WLceXk/pyLVZTEe0uDnfFROypYlzKd1moOk7GcM6ERTIQKlLTJPFZw4FDT5r2SLq7FFlD
VxoovX5wCEloXybjHj4rs/YaO7CTUYBqacZhU/GAqZcMvS3IlfJs/1r1dto5mbD11nOsNoGG7Il5
9xRDYVFYFj/CHWnsnV4pOgRr2H3DIyttnN3vnddjoBIkCzhd2T1auZs/5NVVyPshKhbBbGj5Gq3K
HsWByLitjQnIG+3WEtShvPLSYvAn0rLTpPnx7AWTgXyFXCDSzjLve5jzv5rHkZEjDz7Xr+/snAE9
M1ocgXSf/VwHv+JfWm1UVU1ocr4Y7XOC79VO9m2cBESNOe7hlkXA4fClTnIntorNGYGy6fjJ/sxg
KxD80dcSYwNenmCiKGVjz68L91QNj46gKFbM9s3sqBCFpYDW+c9pm7GHHykxSiIkX8GljTaxPV+n
ItiE4WO4tc9HNZzG14NKk1v4rpz6YCEFuyThWYSYvq/QKfukyLQBgi875f0aowZnIgA1aPLeRi1e
CqYAqEuISRrnqItgXofhUItRT+OYu5Uw85GlNYpfIjygmiA/R1PHgJQ6U2l7gjZdkG1q0ti3vdDv
ymuOE7neLIWCsr76PazLcpajdzm55xNd9ry9JOhlWwStTNCFf4FrhPV72JHRgC+g9M4/3jCFWgNH
wqVzKdD3B2DVhE9cf3opIiY/er9hLAr0h5D0xRRMAm1cK3qedV6jLV9crPjyd8Gw1OqtiiXF3QNm
2ALqAdFUp4qZ2cP5ZBbnbvlvwuzEdtEZqylE9t3bVIiv3/H+MQPBQiRedcDRI6MUy9tZVdhpU5F6
y9EsY6B4jAJDUecYgLI6vxky9nMlXlinL5cgkgsVFG4lp3C6WXimdwWgXGgZ4wQDTm5Yq92fKiI2
WBX/e/S7LG4HDBD8ahmoDDvCk7WzVgJkfudG/txCmzPOMpaGIhEUZo7xq7XAFT8mQe8xnEBJK0dn
zKGmCGXWhNxbJPdDhMDfRxc/+BeK/BhVU62OmA3ait+UpphrLatdxV3xfE4qJGIb7ywI8JfJLc9Q
TUBWhyJys9AkG2UPsvc+6b3SwfwvGlvOQ0iD1so0VS9nB6kcP3MXIZKlIViQbys9b1paN3rDZ4NR
V9D9a8WwJRoqnCdTDgLa8KHw/mAsao4kIe45C1UgwkttgidMtquP2EnNJ+cICDTONXSyY2MiwawG
y/l9dXzH1n5s7I8IWCmOoWyk/GNSWih+vq2u/9EY+n4FHUQhtDkICBP+3YW0xui5DZqBBx7HE3J8
YeGd8A+SXqM/3R7DSrU5ktnnVRRdq0pBM/rk8W2l9+HQf7wTDABS0TonX2NECC5FU7aVguBtbhk4
g3cw4f73Wkafgll05156Skni8ecBknQmMY3kdp1gmIRZdfIfzrX4UNBKAMEd5KMQSYvtJ1iIT2ug
j0UqneJnKLbPY+jp1LcLfWoGM/QIpS05Hr6sJUDd8zBwTZjZsDlb2Z3ZLuH63yF76pGYGJBXbdE7
7JvORmkT/o+TZ03EIArN/P7dEMIG1lGNHSm7KKtpn068DOyJjnON+aSZRY9BM5Xl3Ad4FHuvag/X
lPgz6mA4l9NZZA6Zyu5ua7m4EbWp0W0IF04s4jkR31B00Q8zBvLZAQ1aeFR9iYP3BUvD8zx+YvOI
QA23dMSG7XNpYGMmYh4EspWIhi7gUOCt2NYyp4Wr+nbVZ0hfEg63p/4LKS/QRXisZdbyRdybpvth
quP1nUe/UOiTXTIFo8CiAfkziFTg7VwLze8dRe5aKY0D/lcGlYpTT5TINO7Eeu+FyYbDy7Ldf0GZ
mzjlDTH1LqOIdvDpX/ddtXCrZUqhThJUJyMbru1NofetKpaHaHvWWqdukht4iHv/HmsO0eUIa3FM
RmabF6BTdsmFnMqYUx+skhP8z0MC5llZzLfUnX1Hj5HrIxV5D9QaXm1KbmjlaPm2kkXyCf+FaKxz
RyJAnWdma/2a9ycLh48U2cBFSQBXC6Pfu+ehMlSi+pdAE2w/nH7ADJmpMRwI0p4IGC85mpqp2lpQ
kB75MBnDiw/0L8lhVQMah8NGsBSVJ3KXhrw/+c5vMBS9OVEeFdbsB3lSZjP1UM9tSeYUoSFNoUtF
GHTMXXbhsVW5NeZZB36pq6KBp8vFWcm3XYjfBvjNaqlUbSAkboKyO2WwRyKCuKdR75MX59n/pS5C
XPgX9C/eSHC6nJhB6QGbD+80SSO/OQ4jrbnYSmPBHZYd1j3RqMOS9HmXAsoDldWezUnZkz6eUkaV
1tuFKu70ADUkVpW9DpFsBrMdu+FhyMl+L6RJ8BBtVKHERmDMtD7AEhoCRwxGHDyJ2N8sqNr2hV2X
LkquldQ84ZBhSSavkIYTCy6D++1doYsuPYeE04U2Q8Re896/siYKqVL5D2+/rMFiyYUp1z6S1Vlb
bVIxs5cFOTOdW4UX34ULsqfFnrHab3oT/W1rVKVTcb7pUSheVPQj7iNstj4ri2PjkCl+HbfM/bi2
we9l7ufnJsoGHudvPiAmBDfVIV41cw0EfC9VffIo59fPC3bsBFfq1L78VpF3nPySsoXsS+0PTKTX
vuPmvOzpjGCQiWMH1cxBoV2d8tbxy2CZ9JVXsc4wq72iVB7JUvPMQ8Q4tRPK6DztqixOAHEpgBdM
6xiqXhXbTiVGuvnSAU5tbKbwAa8mzhI37yHqgHUbifGFRXFqHtQvDF0jhMlLcSG6qw/Fg+yLC01Z
IMXfCjwNeSEju0BRxvDxU0ONCi6QYmHH685KSb9LlipeCHzoAxOMeqHBz122iSYDX1RFwvxcaS5O
f3Nj9a4PHHRCfAcXq5Fxq2xWzC93dskFbvyAA29m8NGoHGv6n26FbPYLDmd+tbeIDKq/wmDMfjU1
XGHls7aQXS4laTcdJg9P+zJ4KsxNtvg+Om+PhwRd6cohObws9PhAe9rSKHvvHtBdOF+QDOtMqisC
0RNULjXwZzGALb2/OR5sJKdtlvmW9Tzs63EmjrVES5J2WDLSFAYwk1GXUtc4fLiuCbSPE+DvykRI
/qdL1Su2kgohLbqIj7488CqWQ78etU2dYCRo8GKRcQya8v9vaU0/m9Pu+6NMEUfXbnVeDoYIuXTn
VBbS2Vrk4RCjO0ya+ZdPotV9+itaHMC23QPZtLhrjIECM76OzNQYNaKq+bgtIOVS2C679B9e5uEM
d/DzgeBTUIKIZeoY0VRqMmiycp63ATW9epZuGNPabEfSjpQz/p1LswpgNXAsSXqUwpC6EU/Cpcg6
8q0MTFONwjGRwOiJBt1MMf6eGK2ZsuVmqPeGkDGFTQqLI3U6bkBPTZG6rrYjI9yRT1KRHfF5/XRy
7LIQWC5IPKe3/9XcwB7/TnefeQ0ZUrcZug2f8sZNCk5uvuI1lK/CdzPmAduJhrkFSpd3rxKxj0fa
wq5VxJddtdwEyRroD/0x6svet6X7DOoAfXXwlNuDEQ/gj6Zzj40Xx/yEnXpxrqdcrvY1id4B6ljY
a+51QQWwzOeLi5lHyeBl8vsCKnFQSeX6tvGYg1LpmbxXHmRSgdhKriRZqGXMeJ8DSjQASQ4Nca/5
YGUFhMjiwQoDOvDc5Qx/faKQiJyGLn/mtFSrfS2YrBxOtBFMDa+d8Aio3T/XuW+ZGbakkMgdesiu
k60X+wRsuK0kXhXNSaEcJpNGuwfz5RUn0qarJ+t7yEhJhTWWg/xZdN+r2JbM9tANZjgXU+petGj0
updx/pBWsSv6rAHZF5DmQbqYObWDY0TP5gytcml5MH5C42n5ZV1MbhQJR9v2ewAEhjdkl5dMHFjS
xkUJa8fMDatNzdHhbiFXrNoJ2J+aZfnQjC1ARur/76L0xG+PFFECD+pH15v9ohDEM5k2baP/hFDd
S/c1TeFXCWRj5iKSHPn5nUIAJBZOVB6S5SnOnIaXS7MfwSLkjOwIYMoZ5Y49mzaSXGT/VDxi/6Jm
6aBT3fzK4Q7xb1o/HmpguVIu5eHditRP56qyity9NbOrR2QHYMgb+CHdJAgNEGbipHpaifJ1vY4F
EMPpgD47kgb706U+CsMA8xBKHaylIdGMRH13dgaBmtxkq5D/m2Bi7BKfiUhsTY02CVrfvMGTT6wI
+AwRtlKRELzmFMdcn/rldec80edzSJbVuocASsyoeDfvGJQo0mH5YBhvQc27RqdFTKplu2I/Wi7R
WwLt2BzF+YuieEXYcticGpysk0CvngHg6Ho6ig/VZ14Qvb7ky5OJkpoDUzg1oskawQIWR2jEo3j8
zpJTEPfq9f3mTiPOO7IC3kBbMEWoW6FVCqY3aF3ZQQWYLY0rLcdQ22n6xelbSP0rJ1ExMrLPhEm9
LpyY4bYqLsmqm+cB72f930G8axpLDviT6kBCQAEjMh53mvCiZNAC+blHWegNEDczWYxiEOhs5/DK
YXcfIhFq9JVkQ5ltw9WOtW+lHX/seZnMYjHRs8auUJdNY/GxsxAsQF3Gm8zgnzkDcpQahkWoE9Rn
UBo2T28r29KHBYkCXaVLzIldHAzmYw5wcqNreYRI6S7Wbt3KYQaxxZL1LTdXSWVhPwUixmc+yBdH
IqEL4BXWehDXcbswb1DdqvVx/Xc0cx2f2+bnfNyFvDGSuSZgKk6KaTNkUNqsi//Zuz/JXuLVpiUi
OqO2PxctGcnIwR7wSt8mIvysWZAJzXj/Hmlcdn/dP+GJr/IiE9HGfAYcsW3gSYBbaDqB0FnvsZrF
fJQvOhdiNRiCtmCLgsNJVVCU5j9tdmCYjYdU61g4SXtrc9RTbM4cBdVYqDjnm1teeJJPz5HarSFv
/jvcZg+BzoQhSpkzHhDmqL/x7MFfCW1a+11guxhtQIDQysbbXC/yREgjPFP4+AoN4IKE/UYdVy92
eQQI3D3K7Cz2UmWLac2PspTER5M+/KTDgQXJgOAejhg+oEkF/oQv5dzzn12pSxNQ6eHtOOtwZBUY
iihP69aKbOML7l+vEpi5baiDngZIiyuLmMforcShUH8ds5HCck7wVG1a/o7CbI6f9BTDnIGHJ6rf
dHUAhLN/WU1OqJbWGP5y1NRn9sVSEEIJw7Nss3EBCUQXZJV7zphUn1ML+vl5+NDDBObs04K2IdkA
VFozB/eoGBw/Ex7zpss+s9lNxEf+8+C27a41/H1AWclENxYdQH4ozMEHBl6rluVDFQhX2qWjYEc/
XhsQUAuvv5wVhWS0edP6PnFheWOTHioTlT2W9fiYfDkD18nUGA5gDziOR+k5NZ3MRxQMA5R2qvM2
xw+u4hkgm9dOrmWa5DpJbdFbWGYt20XHAvF0m+NEX/a331MKjnMTkzag1DhEsW0gO98qAMn9XyoN
UwzbZ1PsyJhgv3Wv11PSqNDBbq6JS4JddpHvGuRvOzHyp0yVs1ZWYspW5p5xkcPoD1ICY6kD1oTe
7y7EmNcQey9xcED65SroK3ApbA2/PX8L83L9i8LyH0eeJfAKKTYF8X+zFFxJLoJSnAqeh7EqN7Fu
eAL0mD043Yjl9MTiOQmf5+OnFJh8Na+deynLOoKp6qopYEKvJarIq9tAvVS3pZX5UpXjs3YWOKBw
V7kcBF1Y5xXELsoEqLKEbxLMJkgYirPnBQnkco+0sXqr2R1X4CsqDiEo9s0yOhzPAdcxVDNeKhdr
+tM55UveoGYo0TCbEMEM24GCtKmXU8Zvgw1uuz+GFfFZOohRf/rhYPR/wYLPt/HMsQly4moqlFPC
08F+F2I7vpDNFH8D08WVkZ1y4Z0ZcwQ+TpoqZ+FeiFYadJGhtlYjH1kDU5j6y3zP3AOO+Ayknd8T
FvJaQ1Vf1BgFNb2pHgASjde6iC5cBwEsvg2HPMILPOKlkMPiukCMl1yygSHrs+ze0IqIRWK0zK/n
Sd7wwLR4tNYeyWLXD0nPh/9OyLknL+wIkq41V3Q4p/3AaAEblG5f9wUs0OiPR0Z58IUVlcwPEzHi
n1otLnVnENyix1A7aykl9C3dsqH4F8zMiloTwqp28p1UuYqVIzEtWVVljlkpuAknBHJg41aHFzuB
ncyV7h2HUoLIRlD+lyGFfkcBEsvE48kv/mxxOLVW9SPMULsobKfVNvo0m9/l8z/MxAmybk070ucT
vV+qLxHu7gxKKmoXcN5aEDQ/93hP6qLTF17s+Quy8JeD7G5A6yI+zJwxxTCKF9jvO5MZlYtCm0y9
aYpcEspOMboHqSg7Uj6C/Uyrrz1EIOYdupMm1iJfxSAFnXUXX5HGZTKmbqeND/kqebWPhT631Qli
AZhFFz+dLDjeqWVhry/KJXzzW+aExAOYG9dXqyS8AedzUmzzlZlrQ5AVwJjAcX1LZXq8CHVF3cgk
yaeHtQgOrZxfUkaw7XTvXEBHPG84CvpOptneVONi9MAttoKyl1+nK4v67x2+tJpGuOpVFBrkgzar
bp+m6Vju5BykHr1HCSZfdSDLJ6DIjcHWqa8+77Iv3vbqgcAO3ns21O0DowGnpWmueT9EiSgL1c2G
r9BTe7oBwJn866hecmo/3zBOos5FBBkHsAG25mQT6kY5EVTAMqMKc57WlznP0fsh+TGocmPibzR5
HGpUA+9UxumVBOT8CvH808Hvn++KtTWMPxhlmeIfExZtMGz7KAMXUxreFSULAa7TbOxr/igp38VM
KDoPAZYSEmlj4j/ydmPZWObrljzjVghQlHmLSziPYvE4wV3LS8d0p2IGmCWcaCSGTIYvezuwwkYb
FARkH4xtf0kM1QDsj0Zh/LdJ9PBLiForiA6D+XAR0JSh4BNyFyjzxZprEexapb2sMchjK0mjbBUo
lN5r++fVmnqdhvTVWBqhoDoXeDOHe52Q6J8XENjp7iyfIJ1NsSG919t8qmqRWwCOEPwWQUyV78TB
1JLWLWFaY7k6t5BrsjqNB+G0CCkjlpVB4wgoLDPJkgzU5MHfhQdeJEbsy1DfK+xkwS3cn+e139FQ
Hco2HhnES+TW+sdS4MSf2iEyjzgFT8A5JtRJSXqstALSqNKBEbNOJhltbwMOmPCKTDjTHVfFhiJt
EXYtN4Zb9zjv3ixne867A6ABZDz1qe59a4Hl1AGGnJ3mO0dNEA1URHoyLGBmgZs0UEzdEDBkRTzd
QgsQOTXxs3lhkhlMb8UACsqNyEt0M0HQPSXT663Iwk09itS0k+JXgGo+n/ZkxnNepMNVp8TdsW6Q
2HdJ/J3lLmDgSXPeIMq5Us8wcDVaimk76qnJEqPfQB9XmYyzysJQwzkNQ96REfAC2JKXugsoBE4r
kvfIhGhrPfH/wwGmMQZgPEWzDluMwZcXjTC1LVCTabcVVKO5Rzj1cX1Ek4rAC4nRtDnnE1dN8gQ4
05CjCjjwrpEeOv8zBli+4aMJOv7ajObYqr9F1YjyLwlQwLjXU3bqY3wsXt9Qt95kkfJToEqhFipB
/gcC7mmUHIrklrW7cC8hRJqAEOnZJwtOBWZVS6NCOlKiqjyBzJ4Cg+DQJ/1vReF/bkpFNzcxs2I8
xw0BmZEFt6hZLa0H4wBfmQVVviCb5vq3X3ARdusVHBYgvQTz9R0XB+GWfLBGFAODkBm6r0pfsTuO
Jz7lPzCBYtW9Q6gJGdz9SGT6/6yg5OlYM+LkjtYXjwSIei+q2i87zIH/dgu/WN5guK2+jzGRotd7
iy5Vu4VVjlc/W5nCDrepe7XvWKse+CYxAdQmqY/Yf7x+PnT3PGkAHDEyJ3StjWuEvfNGuXbzCx9L
S314LNvAOrDNSExVBhGthW245qIrzu33ix/yypWvxQCMTPhItfiw+y77JEDzFZ/I7SC3/6BFyLdA
OBCXJcNMz2i0qXsCm1cYND9oF4/C/nL5PjPntKaZ+AkTV+y++m+1kvlgyYXwIiMdGKl0MaQtTjfZ
hmSMzliLQ8NBmBSN0Xk1wKvx7kAlTmbCfdYzyb728ZSBchIX5gq9cPQK1nPs7rI/H4DiEKEwpx5l
DB9QMLo4Shb3NBmhGj3XXKwRow4hCTvu2behd3X+5xWequLfpTkoGnAxG9q2LuyTbWqmDdP3jk1D
2kT8PmdRFLzzNYsxqoE1wIFiRRdltv3Fhmo1jDRh7oNMGNTcuawY0TXnSor8Ov0OjOI3qtGQbvqP
cmOm5olttnoUGd6Ag0fVi+HKXE3FEPQT5OoC3aGyEzTsNHhuaMYNzQbd1jbkqMy7LNPPiYHZ2V/g
rzbYaeH/RfXs7xPq2QdyjWytZ/Ek/k2Q8rpwZER2xvtbwjxDmRtLNRFJHY7iPlLG7cIcSObp1pkv
C/IwrL19HUBBXS0ZC6rb6SjuauSgLHewRadmYl7ihNyymAtDTGReZaewgkDr5DFQNDnLC1ldMJeR
+CTwsUfDB7UO7Eky4kwOJF7rriTX0fhFSskvh9fo9EO5PFabuPC4s6DNUMcZHVxCENp6K5OxpQ/P
Rm+q1Xmj2VSuuPdGYn+61o6lwbzxrjmEQP37YGPkTZPTZUSVkkUErBrCCOdJ0b2BSTAJUQWwcoxf
FW7XbzZRi5EyqUHMB4o31b1aIEwfz37fNjd67r2oBiEIya9iY6jCo9dUJwZaSMFirAKsf12uM6tu
MeBUFr0mcl9spIUMMvHHRqWfTiWN+oLqTN66KBolzKE8FkarXdK8oPq35dRnnDD41BIkt3BxOXtB
OmQo2A4UxH+mRWhkdy+xYpHd1plda778PS3aHWLwqp+JA/kOOi9TRMZg8qtZIdMaf7SDeLsGRuP4
aaeX3gCQI/3pf+By/pN6mhuBdiD4m5nDu/saLpSqiH8RLAJS6PN5vC4yROU5cR/cuH4H4xOFNv99
28JET4c+S4sBUxXwzS0lcqF8kcdmdxE3JBPglDGe0c3aPKG76kMXW0grsFHzeqJyQWZNqX7pT+qU
JMIkfIlGFto+YgwY2WCrZ1oJ1edx2yH7TzDK38q8GHhNqs7F+1ATg0QFzqBefHaWmOxEF2wZySXR
TIavLs677sCXSMwLM9NJxMbB/M3qVWxQqggWe5NQVKvwOIRPfvrubrqQfGimmoTWpGu4q/Ovh6WY
pxAYKXU/MRFkaQUDAn7LVmPZo073HkpMnkNoZFJ43Y5kPCSl0Xy99s6EG2WgyW0S0r2qN+AVWVRw
G7AC23OusVwDQdP0naSq2u46uCGyVvVPF52EHgyE98C6kfRDDWTxU+odChEewz+kz6nAjrFW3ngp
axDr58Bz66rIl9eomnbxaKewMq6uXY4ot2wyuVhv1Af+Mu3cvW2umlLMUIWaVzK6pdU2FMQP4GRD
mkT5xrY8nX8ICMmjmI/ADhsrhCMhIhe7iBGet2ySVcZ5EKm3IIJO32f7Hgbv+mCxCoD4kAN+en5R
5XV2WLcXzLFpxgrl02misTxwjQ31G3AmBE3xXcA3VtR1mUMU6XnzHzpLZnr77MiF9mTrCCb1jJ+k
RieYL2p4Mthq0iGjgC8oX7v+soZ4VZ6j6DLyRc+jyoqMoJTU9D2ZHt2ZSyC/y8equfhcDjazTP1j
lbChm+SkCi5O/RhaxZkstsHOvYB+uPH3pTlSOwQLKwKrzAbpChe1wO4smViWCo6kfiQIBOVThpd9
SOmCHHvwJrT7fbtB7D8tT4hj2ycHnY9KRHKUG0eJl/R8mAmzlwOaB5iHFTJu+hzIdjr+o2D4jKEH
weqneARmXUb3MI88+o2Zf0aCSY8dCQTx9QrAwItwbnHpDSzGZor0w2VvQgOFKlAztAdG12+FJHJE
+XTdIVSQpK2VnfGEjoNWFksP+t+TH1RzpsvbnXxAvg/yZX/vi3dvKscE25e8jr8XybqYKOnMJP0Y
5KsZqFi366wkcqvdTsJkO4xuepjqVlrW4LWHC7W57SupdRkyVTHf/BKH0o+ObPAC86IzBh1uxcOW
w1/nCWXhI4M2reYf6H81nq27sCCi6QcRbsMa074jMh0Vwade0bPLRK1nJ+0xbbnYEI7qkxeGvKd4
OnQ1q31zBl91UZsRYGocx+EIN2FrDB0Q1uxKepTtNl4NdZBNWt0R5vV2SOLczNDUJbT5ABIKzKar
KU6Wdnl+36CywHhe4qJb3sgHaDCnQtuEgUTqKWT7Tip9LvWpsHapENEyOsRwwwp1Uj2V/fWSkv+h
S6gdVYFlv8kV3vUjxCHyZqBbHlc7bvW6GyyaTp8cGq2t/1BH0Qz9kWKKROYFKv63H7WfCPFxFZaN
TD3GBsZSlUXb3AUaMX0caDtd8AEzBQa2H2MJOaDWhO6jBjMGGMlVIr9cEWRxM7LVjr8N8NFP1b32
4gHMnX56IhZJWmUvp77uzoQ7YCnIL15RBOIDkhw1J6xdsSqyz2qjXtEx9SfVgRCWDbgDI+4350NK
kgpbJQMurW1eOuBawX1lDuFqfFT34tusmc7H7nknpcILIHnPbFfjyt7olLsXdokZuipG5Tqg8acg
AjsTc10a9Qf/MnLqZXY40lufcNL9R9SH4O3P+7R9R+rakTaAH0EXjFLHJxzMFqiIBPgZJqIsuTz1
Ai3KEL4JrkYP3Jm1H9x+/0mpbZ5xrfHx/eNtFDiQ9CH9zdI+PaV4vCExYRK0FlZ2pDVO7ysig1fX
UWBneJbYxBNU5dF6Xde633Zyis3FS1TpvcBw2e7ZnQHwZ6U98s97/Rpz2kbhk0N5InluxVPthKNY
NM480JrozZJ0LYJP/BeKktW3vuWzN4Ub3dG4WRsNRL7CtnfYy348R6kf3veRb2p5MrmwUwuvmQIF
cOumSxATNXdRwumNI1GTxYh8+l3FvNdAhFVRW8KuWGu4MGPTVpgK4Qwz90QYgRmh2d2wL6Z+KsjV
T2xUbrJxuO/6QIkadJO+O/zuxtcfPFFa8DYE+65P3ACegR/FlZMg/sgnuWJOk2M27PStXfIvR8He
yf41hddT5k/d41jcifYaY/MoCYVysGFlPMxlQDhVsnihleO6vLkSq3nEAC+Jf29NYz2vfPA8IjsL
Tqk4t1+ZlByKL/2J4AAjZhmIGtfgsLmZYCKAlBVHHHDJzkzehYtQsTitBwX8nqr39m40gQX4LDIj
NjA/7G3NWC+NgP3GZksmbDGbL+FUajaKvtk05qbCr+B5bXvHH5sAEudIcWlLj/Y1zbParR7YGSN4
qcquA79i5ND6frraMHkOjxFQviWifbXiHf3FT7PlPFVyCLp+hKb8oKi/2VKnT7Xovft2cTniEh2q
JU/dNG6K3pAMYxDGiAP3xE22r6YlxPcW3B7P7vGWvBFNJ3pYua03Qk4WAIl9QJnQaL+uEzen10in
o0TMt+jKq3xZNI9ziGzLxHKhNWvWtTIeq5GEcZkqjDHX4/4Wa6cKKxtLx1xdwBGMMojtezLZGrvu
mlVFcTu1BQafrgMEhEtBE9R5O+XX57WZ/k2zqPz5sNbSBP4iERXc1St1IpPPxr5hYmTgJTMNwN4U
29f6BFmEcSPyEXwONirJmBK3Ikf2TSIFBIiLlzQFJID4DmiG26KvtHWpVVFZIW07yg4uz1J7B6w+
YqgghcNY0Pmufg5FUs4BndNdOO8eBgkhsprh0Wo1kgjXlOlwF/UytYh7puj5iexQj0lRpfMfWuJd
Tsk/oIf+qhHCz/p/EYLclEavQr+4zKTKWe9dfmCthXPIwHDxSGAb3zIIdaoQ2Wg3m+/UwZCSWdKq
XGXtHRo471C7ri7kAJyhJqETJqrqNRuOd+yMY/CxpjgnRty1uXMO69T8dy5HJH2SDDgj2AuI8iP0
1YIH8HWUsbnm8JUgWUVqGk4H/aSSo38RpLF5e60aPjaihvMM+P+uMFTshx2anSKsCfcludeCzEZ0
ayUctAqhHJQyFkXBNTrv/tZOWR6HGwjXorymfJoeliE1caBl83tvwID/p7JGvJujtsNBt+TRuoMP
xv/ScL1JSlJMngGzAIAQbZLeKE5GNK1JdV4mG04RsAd6M+Ep8xnMUueZxppGheBsIGSeYTskgtNb
8vH30ahD/IuqvnotgLo2mRHIupd0nUwF8MFT3c25BObjqFkQRVIFGmJZ3IjBHnbwzxFpD7mMKLVW
deBx7jgoUvDzMTTy7vMNm3ROyWh/62cnY5zeNjfd21Ab3BztkiBBzUE0JyNFDvLduzPeUHWPpQph
D8yvuGzFuLQf1e4msFDzHo7V0h8qw+Z8q2TFCB6EcF6li57QlKWgk4Gmql/xgJ5aL5oYbrRClu9n
sLbicVMbO2cZLy5OMtiFRx3/Q99iQHPtkELCiXsuQJXEOGA58BrTFAVjTLSkxvmGzGgdXDHSemwd
3C9FNpJdyw5HUJwyv+vVXnrz+YIozZy7bdNnkBvkievUI2YSF8yE1722brQX6l8VBLYE5OX9a8+L
Sfx7851YzMiuelmdlHbtx4OjO3UCgFiltAqmC6gVm9fAPzaF2q48jZicQrUJEv7557qrStlzENhG
W7D2ufPA4nIh8crtmXmb0mpptGbEn6zpR+DB0jIoQckSQ+I6wcs/2b5MhHjZbzLrWeviEgvW2hy7
xzgvWeEwM4hmNkH70qH5HQaPksLejn/q54COX1aWgxiXUknhHTJc/ZjuHYouYTzeQz+RdNqjNBGP
bcouKiCO0U7swG9TTowysRYgME29ANQXU9CYqz6NVQaIveE5TPtvPNw0AX0QEX1FxteRhfQeuGIZ
hHGzGD6FFLy6WKM67EVmHpu+xRtGQfOIEHNItfgP8o6EVFLG+Buvy+2PBnJ2duCG38UcaiXVf/HQ
ImiNQud9Vo8i+zRi8i26WzLDiEoR9OkEF3KuSlrsAY8Cb+ixdZ2fPqkpwtbGy+btaiR9VFTMgepQ
Y2eczLcGHR3XmbJ5WujeR97FwCtVrbjQOwpgiqelEr8VSWzxxypxqqBLe9WWJ8/v3XT7mpCC3y71
GOzMcRun3TuYGRSt5Y0ghApoo8XhbS9fZL7d8dKKn2yJ3gHxOfBFxRR3/hOhDI2GDSxw1AfvCjTh
QHqc0b3CixS6TJZal8vZY/OudgNemyYssHswY3zXTMHc3+ApPMN+qGBn2SsZyK2A1tB0OdK9SPXV
ducamCZQRq3RyUkpwulOOusDP8cTQWL2mRnC8b3+o0DDf4+rT3aoe9LYjSk+fGo8CSj+PQbWIo93
e0/tuLU96K3VCrKtarxA2khQADtUT2olW6iNyZQ7IfEEWseJBnf8katAAJ/scr7cYSCltp8/5mjD
2eJw70uxb3ytKiFZnoGnxvn97jgKMnS1kDCSGoL1NHd9zvfc4m9x5BM2v+eQ2awP5Qk9QzFi9nKz
bKlQhuefYKM3LxV6V1wSPzD8WACLGWpN4K9cM2DEseYZab8K/N5yqsx1NFH+oMojy9RXzzkRht+Q
wER9dObVad+w3TtAYJQ4Qp3MRnJwK5cYhcLxlQD8YdztrtYgCDOqQMf6TkvzZ7gh3m5wxKCgLaCO
3C6JRoiigw==
`protect end_protected

