

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QHA3Ex+CmcwhHYj/Cu3wGvj9D2Oh5X/PuqFEaH2NXNQZh8T+UDvbmRy04SPk/2ZNtGxTEFpvVC+A
OCZnLDmVBA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EpCFyIVFCjVsV8JAoVIvFxgMicPOE+gA797pZe0ptQ+JWzBRfe+ko7I0AJCcVXyK67/23E/Rmn28
26K0nfbqlZMWRo08GQzdo2Pvg+0zdb5xynhVYesyBJF810yAmWPUXibisA0Uz4hy5us4urGRvXui
1VlpuDGRFz8HEMlbkMQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H91qDFpDLhLKyu2zO0jS/sr50G0AneZOioO9iB+qoJcFLnwgo0vpwwtqzJX6wbDVN15cu+R/IWxt
dEt2vBf8d1vLuMo7BshJZtbUM8fTrhTZcFoSdUQSe1qC2oLTy/DpceJuEMWuDApMg7w81zUOWyVZ
l0ZQx93l6uEMApiR26abzikEl3AMNYgld7204pP+LGkuQpEm5BNdhJ2R1igYEH2SLr9PoNXl6Ybr
Jw60dHycu/SF1aZZvyjj/k0RqWzkWo9OF2bMBdwweatK0hL4Za0tR1dkbQIVANMFXr81aRAsb+LC
ySA4CauSi00Vi5Uc9EthY+ZLgX5Ay9HkzjDp/A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UQgJtyN6NYDXy0tjNwGtkb8soUmLxZJVzWlNkhMS/C4JfTEXUPg+A6vy121UgFOz3JMSNyezviZf
Mfex2hTID+DH3Y/f+mS9lvkRe2ugr1UrbCWMuo61hHhoeO3FlSVy5OojiRVr0pFZAlcHpyRyAMDC
2ubNAtCqnKhJ4O0W2nXkasQr4eFt+GOK6JSg9BIu0PcXYnr8Z96U14IqU8qoaCFnjmOffa4iFoKt
fCItpLPWXVs7vpK32UsZ6CdWATv1DRVa7rvpoKAYhB3pTdLEGiZwBFovoFut6DljSNKFNe31ZoBh
ZvEnbvlCLpTfwwRuxQIxsF7NsbghGxInSwNF7w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GLlPz8clXjBHUAybAGhYboHKfTw7ps5cfHItKbfGW0Maog/3BI94ghpter+alXbAkH+8KTGFy2Ck
42pN270kZeA0uP8+FP5FX9Hdxx1rjSJSYnLaETC59zrF0zNRHR2eUpWdzjk3Q0IyjEcI0hzDMWpB
BTUA2W+6VKIt7CwOChCNccifqqqM2/lE7U6SRri20DGmnKYCeA4SLYKMVgbYiwIQ1WpXXJqIDpo1
bsC7dc9a1YP5bjwk8u1LIhPncODSxREUNUwGR1Xb9he8Nu6GvsazhQaKR+ckU3zv9ioeFohkv8YC
6S+WxXXst2ppErBUJHaQ9VRsWjop1VaIGfPf6Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NOuQSwyLor/NCRAPbb+hLF/fWkzD7blUj5CmRCbO6PxyE6eUcw2hCJ3syd0WNFx3AwuOr2lG8SgF
2djEMbP+862p4gxkXmmNOf7tGqVDHgC/fgmOIsxfkZ95hvRAcEvi1RVx++fS0h6KGuC39yN9BrTt
nmZ8JjVs3v/ky9THrn4=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BP26diD8XpcagtcJpVVq+RbpugiTQYYy381rJIl+lewz0g2oe3rZrSn4SemKHDAtULgIN2oNIFYj
pWqaeK5KLTW0n4xvkxIsB7rciQ726nTjcRddBUmvF25tkhA3Y3UhvL2S3bElyqF4lCnStpJABIFq
XT3R+Lyq40nBC3EXTPszZosjTkHBl3uO8EFhwXxLaoSimXXGgappLzUn6dp03J+zr78NjVyMcx18
lwiud2D8+5QyO+QXigVTSDyD/Zd1vaDmZ5CVwxsypJWCKZ2A3qx4HCL5RoXw/1eLwI03EXKqEgVE
P4uFzHRwLGNImIZpDLhj8SnU8I0lOUFiGGuDRg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132672)
`protect data_block
jymTfeAuyg5cflwDb3j+l+64lLxhS/MQBaDYq7mIYtiXMzoBmEoDlJCHszHzs6NXrd6Hc08j8jxd
oaADK2d9J1iCm0Goen1KABPNca9P+xqkimavq5AbEf08MQ+BEe7+kmkob/vcPv1odYf8uJXU2duL
Bqu7BTjE4rN3ryV+BzPGeJOOCYGKDSmIKw7IAGE9o6+pRx/A6lLiWY2kZbAR1NcLqVpjPEh/jm+h
i88IdpH3sDN+JyhM6oOTN08CnnrugOmYsFZipS5dy46dCOHN0H31TVsQOsvCeOOW7bU/4yddrfEu
H5gcH6PVRf8q7+Eo2kJBDwP9C6PAY+PipJPnJQt+b/0Ur0EXDlJn/yCQSxsFRz7GQRhIvxdIIfvx
NUj2H/4cQZkewAwGL3KTLAtuMDjIpMRVdc6w1CgXDUOxYOhEgIR4D6s0MiJpmJNgt9Q5dHQYD1dM
dqt8pnjZLhCs9RuiAPUTn3d4dN6TaEF7P3pRxlvchPvaHrayxzEF3+1VtcPu0bzb7304gN6d17oG
CeE3AqRAnISbYuM6FCV8lslrJ2lZX4VIf/hvsEMBpmPiGwIgAPLLAdrruJivKTzXyfKNCVw38myI
UTwut6XtOSZ3Dc4vsjm/7DeB6AaNYvMto5kGDHfJ7FYFhwBO4HdOq+Vc21atpV5ZmoRDY/nSt4VE
F83dNtbcVkoftcSjRJsWAziB8N8J5iVQkAs1LR1gVu54NHhqzHl+44/5D28GWQkrgJusnMRh3BCW
pDa38BSOlAJq+V09Plo1pgcfy9/i6Gy43pq76ThM/CBTnsj4RZcROAOsoBi+p703FtgeNnL+ommW
Cf72JvMhGUXI0Hfs3ruE3+JJqx017V2Qwwz28SPO1dX0RjHrFEDtc66TWfFPDxfHYMXl6z1flDt/
3ycsoSk96oHzeKPcBNI6O/jo1thXRTHXugaf9AK952lWzU5FfSR5RwluHfFP7wERJNqyOk5nktCC
P42lKdYMNz14LXkgcrXGgDYhHnfkMjwg0W+iQtEGjdKdCr189Jtrf8vvavSpVN1OogKCp5qOm1r2
KozwDA/k6Q85Gg2aV+oltZN8AY8xvdyqsTDMay7Tu0DCOHFHXkHoIiWNJMBgFe73xJl+2V/X1A48
5BfFuyb6A6aoFaAO3xGqHCdhrEcVFVRRAzEbY0GvrVugX/oJuIl8KA9PcDCRP23jpuBwmVYhJ4Ti
UPjH+TMSxuP5pQtcodBLmVszf66RFGZCRMSXtuRdGlZGEsCmbrxDiD7vb1A5R3qZQwsMJbcOQFbk
xARkzFPkB/4kQP+ksSz9GZ1Eb2omhH0SoMdg6a0FxS1JT69/sp/DFRvj5qE1iI7BRBbf4zzGGcNT
hcKTRncZ51gP3hB9cCY6H6Ef+iOTzbso9b20COXd9zzL+cd0IXEr1+1iGs97vm/MauZ7EfOcRN2z
Fo1wokv4EEFo/nE1DRAFEdXY/y9aDkXUM5lGzdNR3nCCF6HuTgHw6XFuQu2x9enoIkXsxI/gQ22p
sE021kxGHc/aU5O+9glqRzd4ymXfzbgjGDa/9lIb3ESe+nNM+9BZFckmK4NjasmZBnNOaNz2o5zN
s7ZDVr000Sn5eY7ZZMOLJqL9QtN6Lp7szp5vcSyknuhwRE/81nvfWeHStg+InCaVvsNLcllQzwO9
4tEytG8HRTuxE3KBaxNIzyQM0Gk0+cfcX06bTkS5xJcOdIzLtpP4XAHDhEts26mArU9PykItBgmH
0NDP9d8JLG37TVD/l8xw72GAQE8wKhcs0noHInG33paohY6u7raAlLrkHwajXKcicHLuCrCj+SZw
PB59VaBKBjTXfKUgjq4cURjoF5U6kSIyWEbq6Zxpj0y106K+9DqFyJ1INbPo01Yac5QfKr8Dok7t
qoUoCldUVdbA+TT4v3/cPoZdcYbSXG93WH/QMurdogUXjzq5yf0a1ja2pVCzHtdzCCEoIR5CWfRv
6BKPwDbFIbkzlbgtfj1owqyLon6boNtS95gb+kahLVQSs8z57NHwAYgdZXwoLENpTf+sRjfMe3MC
eLjlBUiM808hFvGJZBQUciPY9aCR86iJyQXtgSgr7XA0H6UP7K5b8WCCw8uZwDeH9WHBMVGq9XrU
B4K9uoskWpTIrexBJ/ByGHNGfwa1pj0mC1pyPlyHdTQhHxMaLSKpGTR8G5z4j0r+/GOFJvEVT3lK
qoiC9oQED6vWEg0Gp6jvjpVj6gHWbIJiKHlVsEIsAvFc3oev91La5u395skK+nmNyYDkQ43gk06Y
nB4lDrkhmSltSh27yn/BxVCJpsyaG36aPObxJZgeKUT46TKcZ/O7fFa46i73ip+Ladd+fRql4hEl
BDx/pTPV8ZB9Clv34svfFFLpziRpXrP4Ldp+lCyMol5CHGBVrOgplZB7g9eGIeKf1MFeyFGrRfFH
/29AtXpERCx8SXW1vGgHcZNNPSlmfl9Pev8mGUz7VGxysheIDCRJAaQOfCfcdQQZITf6zMQKA3l0
ih8pKhF0x5QV96QIzOuWi76Gl9/WhUwyWem+cmroTDModDZi/KHVR/WC6WRzfNrilraPNryg26v6
4RL6UL/GGLG2WJ7addeCMbJfrS2ZF3K5NNBoupdx5HGriTwSz0os6njafXVQ2yEhYSirrvLbZt1x
YU7cVe+QpPBHRd9pKji0Hr7c2Hc5LSwe7d2g0MB3GQY/IfyU5SlASkEQvKchZ+fZOF+cmxx9EkeZ
PWv/aS8kAqGJ2Mpg8GlzlPuDqLT5aVc+mFtSwqZyJ7rUrszbkcOkyZ5rfw9fp56VyGePwKDAJIz0
sm/V8U9xpfz6Hj/eSAQN2qVGkQEQ5WsSKPpIBxfOk04xHjrWdlHfSMo2z8XgTooYyMbxek40sDk9
Jo4/ukVICbe4JTuIFbs1Zm8I5nDJtYdgQj/kgmDfctiePvQsKua+6WW+PVYjroRhiEqlsFGHRJU6
Hn+8Z5b0qBQEMQzPYZjyq2ALbcp0Uv3D+cCo9LzNcVp4C0/DVzHBXgI0f7h7X3fHsApfxl1oBxG7
2anl8NgHXo8ewzroEttWWb6d9efE20tDKX2Te9XXZwPLdbVvyi5Q2P1jqUkVkhR3bZVzyxxmMjF8
dTmakmuxdsr54CYIiUmTQLKhlEXDmAosXnusbRk0E6cNJdKqUKfO09vfyW7aLYlKkj5+4ds5M5qR
vA0JZ4SaFb6uAtYGPYbhhZziKj7/wA1/WgTuiPw1OOfP8VqXWdZDc65/VpLiSZVc7QKiU0SZHk4J
j5kvcnnvcqk1ux1my9r7dQpqv9P6b9KBr3mOkuoWRskXgINzPRJ3XdHMAh/ZB5EDbjNIlI/3OTaP
si0O5vmeizB52YZEw6Qc7BuJpjYCIIHQ6cgaGPW2MW5VwKWUaAN91rYTXtBC5WxjhzVI/vo97fQp
jpHgi83Lo3MNLfZYJRoA572Xfo4s2EAZDY5ay/91mlzh1ljpBtujO0d0c5w9vLddRJPRFSWJkZaO
iXMQIpIKwhYOyNgmBby7cESa9Og3aX9smNl6LyQnZTmAdcdtKCFCGSqaAz1FKaVEZ0ueyhhEaqwi
Vre63qYArHO/AMU3mGT84hqrb25n2vnBJ8e50mFhOMH6EhsosBYaVj+lLNUfsgRQnxmnO/nTfLxw
Lw6f8CztWRfMqVc8TXm9chrxxMwiIJoG5IN7Nd3+1Gy/XFA+KqndyUyxnvPmBYD6XuF7WAHaTyEA
x1+SZEkCh0JzfU7bo3brokrF6MNMHQ9PFax1QF/P9kPf56mtzhk4KUgjFD8YRoeh5rp3hhgQKpwU
dsA/0+raY5Hm9OFW3+wour63J1jsgF526NTBZ5WhFbcCHgnb7QnNo3Tx/3y6M2ZU4U6x11caCAW/
PSMK7Oto6ckv8PhGuJ7HLISZ7flzPSYI3HOML/Cqh/y+Lnurz+5NUAuAzdcxDEPr+Ab7h3+cX0Vy
C6F5AOOUsNHv1ywNCKZfFdV7tyO0TXBTNyuET+fyUI669h4UKKhOhxSf2ukHHIqMHKXSycH1zN/E
0hkjRfN8YWBfj/wpFxssOY4rxmjw+BZMik+B+OTR5wysjXpALkOcRd6XHjX3Pv/CRWbvIcKb/Vg4
0JxW5rtBBpkoYg00GQHBtgNMg+oYnTlQChrqhCQtLASdvdFydvKv7SO5kk9hYf4bVv0XtRxfkCN9
2A1HCI4V8bt+GlARRI9Uj0vsNWU24nWtQtrmS2wvubrLqeInAFphKq1qUXvfamS5uh/diFsMd3pm
R3TIWyds+uJYeS3vdUeMKJQxx5FDk2mOTdyPzPZvD6faFSeI1cKNKEeJmCkPb9KYrOOM6j1GlBG4
P014vSK3jNn87BVaTLptmxz9u7mfKbR7fPvd1zYFPXruDCMTvhSHTCI1BtLzDXBg/eRKFt5MV0Hk
mJ9aUWBjbB/2J8cSDL2QNTrTzVGaARZE0BjbHeqe/ZyG+cynAqUoDfm03vXJhN1o8X1XadWbUq3c
s6M6HDSsSlVVpCYAQGOYrXu2ZxrwnnshyS+rLaOBEMfAOtvv7bJoztpx6WpxG1XLE63mHjhtwUMu
yC3xNbQEwtdSFsSEiehnEsq09+oaB1+aJKRJLqe7UufSKzWfLuC34zSyXTtvFJ5RhZzQxlCkw6A2
l/+MBc4Ls8cYSXRZOpNLycmXMzADfRt8GMjUAuC9zHvwya10GpJDXGC1h8cum/zsAGEQOG/kmRXr
mutri/fVy/ZPix9ubeFtw+9c1uj9ANUnWKrQCAe/MwSk47X7jd12Y/UXSl9hXjjtxfj3CMkotJRj
e8DoIiAVegul/yRgc9pSVB/m2EmFiex667bZnQHByegVGONLCN9jIAjetE+tD3ehYTRy4palF1iJ
c6Uc6WdgM3TOTz0cYVbPzH3tyFBdu2fkfKnRH1a5g1FXpYQBPiYT7PCTE93h0XI5ISk7IVLRhZLH
RyvwvB8ZNYpyU6B2SpTMIssrnTccKdyJ52ylT24XVnLBnrwxuxDlsQwFMRF1U4z9/TMVOHsOePWn
1JEJWr/z/vo/M36x+5e55isJMqXGjEkB4aEz8PdvNvLcsKNgQKCfTbWvbexwkI7jcnIlCprUjq9q
BUBRfuhDxXs08Uj6+YqIuQDGObBZvF1R2yt2d6/IT3k0OOfOSMhqBdJysv5NFO5hYClWkDyGSkK7
YoekDQ4jpA4Owip4j/67RwKFqneK/DH22/0Q3X9Uk1oLMoqus4oVcy4c6GqvSmkdObkdcaCODNNS
IF0OhLzJM3Uz0fa7liDZUwA9+Crh8s9t0ZlkzBDK2SD+l+oCXDuunM0ZqXqyCkr7JEnSE2BAMZfr
cVLb5G5MzCrqaQQ7Vtwx47WrEOiOpkczx44g6GSWV4RGLnohDLkSwvpSwHlTJfEsqd7JsMEjxCjO
g6P3HZrfGPhCYzeCDtdVRVujp7aKv0dAen5aiVSz0iMzJrTO5v0y4ENXLggtmpxEUgtKVQaHdXdv
ewlsT4ksu4fF0dSzNEn0fcew5OaoS51BkKtsMe8JLGk5Uja8logN4JbtpgRmvWuxhC4M9aQdOHJ2
Qisc42hXREiUtcdxrd4f5bNul2EDPBrnhpS3vrIYzR//X6lZfqzGpg4JGne+dVDsolYsfm/FDVOI
zHnOZ/JE9UblQsTrMK2MpZX7VhUZRf0+/nMdEHeWt7PmXpqnyJDRH9rDQPZGUn0KvH2k1gWDUBvL
OPWJczLJGzccYpLb1o6jEkZa2IjRELASAV7/a4a97DB/4L1sgGkuPbe3BjyB0a7pgxl8o8vEdEFE
t7QSryPeSDK+WVEPEzSpg4gV+R6zVerO9vqVYjkMnGw74kp8jGP6Ebo5VSWMCWTXJbeZTXTj6CfB
utgTcyjxwrwr1jzhif4WM26IiphnXZi8Pm+TXA9DMxA5cOSL7PPCaJwXZS+uQd8+SUbUGvK7ciEI
QrWr7e0GQJS0d7td3QuM3xKG0x3fCvzF+2cEPHH4aQoZYus5VZzTVnPflwO9E/qXpK0ehduiw4hZ
RZGtu6sfyJK+0+wfFHPfnif8OxZ9+JF3+WTnHANK0/RvXxsOF1BTjaBvoKpabQM03E97Er4VAdg/
ATRaYKFH4trhXSKBmmyQRSz5g+k450IgJrmRCmzpNHWxLf36DG1dGkqDdCJXd5ltxaXaEmCuZ795
vNhHNEEnsHBudSLi2IJxjOw3c0dR28qQue+tuSR/dwstps5gzVgfucfDZMJChMQyRksUfAZkAyeL
lO0R+T7ee6ayfi2/LR4cYWA0Td6WafDs1EsigYsv2b5VYsD4R59gTqBPh4/AZ/bh7RD8pqTZyk5M
n3M+Rl0n4VCOwBU7G9FZj3Me9iFO/uDkAjJf3+lnIf8YXmPbuWnSpqrj8S4kizmEr8GsOYXF7bhM
ecFQhI52LY4dU7OotXKW44A3kIIK5LPKz+rA/fpK4Uz4+8/4mS06KBVkyXF1/j0OdUQP0wLrml3Q
duPvHNrdLwrmftlY9yCyT9jfwtDWGy80uvuCGIQfVnOEoPgRcz5W4LZJe/xGXkaAvBWysF5auQ3N
mY6NMeiHfi1DIIsz5Im+3tifCvHwte/xCKzVBM/ynC9towms8jGSM6ULAOgmlWKIP0yVLGPTkYC6
Ge+d0uchDL1woeJxNa4xXpWFME/zuM4B8YKfbwE6K62krBQ6N0LuwSmZ3tAAVlzLGEl+emq/c4q/
HNW9pN6r3HXm2x5mCJ5nrgokdzoppUxLf8H7xAidmi4/zIAwZeucyYpFqHteM6ZcVTMp8nqN/xx/
RodcVESLUqLhCAEjpGcjw5AXomjsMWG607j3SDpjnOqDs9btopm59V1w/XrcrfzQvmIkLVJnXBKd
Ps+FzHA/8ZDMqBMenT0LGgnpHGUtPN07p3hpWs4ENV6ZZOzuYYKc0Yfrw672p+O3Zbk5rYUVTKcm
5ejIENldjY/qx0Gy64qa6lQajTmpHi9DTS0Q5FRUnnNo3vv747yeMWlg1ppKCKgWIMHPAgZwFIuq
ZZEl6xTO34af8roH3jfOCZ8kTUPFvIEb5ULQHrAiWok+PlYRPL7yGeRoclQRqk5BPpiZn7daLCfq
S3wkxk7p8DnPuq1GABXX14sLULF0VS+71/jQXdBieE2/P+2CCnQR6YCaB4yZbjQle+lToiuO9bTp
GIcCWaiRAEBFOcW4gJFfQtyZEGueuE0ccYln/Yh8Wz9q+wfSF9P9nvhXO/WVUgCdI0utrk8mkHNb
VAKOTfZhs0QUQDolRIyn4PgCm/w+CCDxcdrvPwnBo4wMAxrnZ9R+wWkZX7smu38sDSsrnUCGTbm7
igQYSwq1NuIGpLVjllOHfEYJDcNi3e10kG3EJAQC0u0N21GpVmDHGTGFBl8exLbDlxBjSg6cdSw7
UEiGUjjVzC851m6/arFSVfm4jrqM73Gc2mkBUt2LJUHaJL/YRY47aLO1tHaxGOdHS/oD7e1diWvJ
BoELUApDXpCUXUACDrZU31FdV4P1wawVTfIROY/abijU0LdlfpE4W7Xuz+c+fkD43ZkGs4KL5Tok
5Lo3brVkue3sQUHBbNZSSiO+g1ljnKdjeWvXKYPlxfLMMOE8PpEo7et1exdG+V0bziyp/p/ZP6v8
an6F54QOqKYO4t31Z6+jWeFAFCB0EL/dmvyQLaTqFCLnVWwGSkpLNBoRzOWxVrGl7Sjfgn/Np8an
CaQ+3ueVRzKAFw7EmJG1htWpzIkWXbh0jsiMU/RuCalOTIrM7CAWHDaTAacXEsr8Ay7Osr8k/Asj
bjl4djvImRibce1eNdzqiVyVLGeXA7eGj9/p81b2UBgNwm8J0oFRfRjVFQB2x1Gx1p0xTIbqE4FO
kX3XYOK7x7yUtbSVLHZ7cw8iVxTvAEaKW+fOiPe71JsDF/iRU2OIFh3uaShnIMJP3Cj9rNq0qDRo
vTya6S5eOg2Ec86WwQx1c9rk792ddwK4HkLxohuxBQfSllXm0Y7eGfOuF/rhYXRmhS2YiKlXnUAj
8aNGtC3ijhIqlYhRr2maHLrIjzkfkIAqMuI2kiNVSCd6BCQCz3/DUQWeQWaDsoTFCN6XacJGKnpD
7CGfkUC6lazITTkR6fLVzwlZiyS3HPii3dvEDENDikyWlpXl9mM6zkGjN+mubrzJLsgzF2tY3aMS
Phoyb117/HFA+bUUCJJD4lYS/qSrGOsv75Rl9b6DUKlLOlKXZ6pUnZ4tz7tP07F84P3RoRyKtJeG
R5M3uoxc43lj9Iyr8C1t9Giha0lgh61tTetSqwu5NGDbFTIidEeDMB6Z8VZK/3lhnzrTs0m9Zt+o
fL6WEqg5qExfkSUpYz6DhEnBkoZgIwZl3VeDiUro5z9sEs+o1NqtBUibOX9dCtI1+LHyJN5aDMJa
y5dN495K9m//ho9DeeKsk5HQS7O+1Gqo6g2z+gbfBvsAHWcRnkY6h5HI+QPqyWDym0S+NLJTMcNL
XVbAP0DGfczolRR/5/NLAjlNVgBXsVGzpOHb3r4eX8FlZ1AocRs8SCFzeStOrsjWxGkNYQK5R4c6
TSYFuRq9UMyCdksGbdblDiAHYZeRIf8c21Txkq/r8U4KYrowX9EaG0BiBLmTPxpEjmTpQd431TOM
GYuBj0DRTMGaHiucrsuyqBNmqgnXo6uxsO/yVuRsb6z7DvcPJ7Ye8odIic4Zil0iGlP19PLgPkPG
oO0960Rtnpc8wkQWm0A4AMy/wrEtHvw2NZoDeIKPf/bOx/X+aGoN5YyNgcRVjAGjtwV1qM2Hpo4I
eSLyhgDyI/pST2SGtyK2KM7pdhFgGpNbkoH6xStDOJ0A/A7oDWEdqM3+eBXV4VwmToO4DH1pNIPk
E0KGOtFTqtdM9f58+m7lmO+a3KwDb5ek/V9E2bLwfSe4qZTak93v+lry7WpwrOslUto2EEguhgzw
FxPPdSXkvFq2FxUq24nj9wmGbMjrY5BnGsF9GsedUEW+TWxrJCV5toNz2GEuvBSQ6bW9oNqs3Cbx
TxFrVsqtkcZ7JwRYZf1T9V5aivAilHB1WgS8MAuGpO0m8Mj7OUTLpW+BBxw7OlT+CqvhWwyeQRMr
865OURskQSX+ww9tGQlaGDfU/GmPJWKMgyaSj3Y+zoPtYB/bBJROSIDK2xGErMOzU04mXePq9ojr
WqIcmpfO1d982uymuzS3i3tXXyiQ1Sa1kJO+f6Gp+wa3Sy3eEaJIcKHIy+XBXRAomjE7N8iS8gzb
WqkaEvjU1H5I7dy97tUy3a2Icxf0Wg1WNjpmAmCCvcYLVLKZxH0wDU/9kroqBezDW3bWoEP4/cQo
vCuGw8gpbf4WTDw/gmUwaQycDz8Z6AbGrjqbDIyLjCdYrPXZpEpeNHd3gqSCMidoeIS3d3ZL1RGl
IXz0eazwsk6RmEWNbNUZLrdmrNBKNLwhyGDFyVHXZqYF+jDIG/EUNIHTzgDjzEl+LyEOfdybaiiw
uPvwKRYdpwhXjk2/0wQ3KngCyEZAfrF7ebxEtVlUiGkPk4yf4jvD5gkDPU8RhbnVml2haMMn7z6V
mzl4F53KcyDLOJ3EypXlJ+PoBrT5TTDw6TFNuR5oWN4q7TKlC/YG8EVYYRGXPsMf/Du3ctzRMd8B
e5gPCqwAcy91Fj53poPo6fo5xYzv/eTp+GU9L82DI5HR+uQrV3Y+j4K/PRfQq3FgZC4OTn/qLIdu
8n7jrA0t7C27SXEGcZ/hWWZ3YXYCAcRP7x4GjQQcokpSRVfpQMgrPFLfgQi52UC7XZk0vAEWZGIe
hAPdbwwX5SFU5G2MIc38NrpUQ4bTF0EshdG95igdrW054xJp1MjDGlu1IndIKnij+qP+3mwCYg/1
sy3mxe7Txm76wnduX0Rkr4DSjC6LiRCOaQOiaOW4s4/mabclc5BnqazbZNlGSTQZLx41WPgjPqwN
GU2mFKagFvNdKTp5gm+CQu4X2DACsh85uyOIANAFWldGSs7rOKg9ymA7O7fTg0ItMHByu4zYV0JL
6m9qlAJTxoxjQK1bqjteknxqtIqhmcB1cTdCTRcbu15DlQCiqQ0w8WcmYBuMS0oEDEUvdy4xnY8m
HJXzPCtp8U5Yo7RwOpRJdj++TB1Rm7yutHSGK9y8mjx+TK1d8tNhiT6esRQrCBQCZb80z5RYAbdG
ABgFCF/SsemPijRICRDbrkGfK81RJUcvPBPyzFH5ppnNHepURonuH2wYgZxhWSybvzEwD4sb3a4j
za2jRl8tsMVhbAsl+S83GT3oIt78YbkpZKnuRi9Oa66fcvHCctBPh6QGz3OqQqPXSeV1g09MqXva
i411BiWVXARFC8+lQ7yt07fgNlx0ywkx+afvZdV25ar5Ggptx/iydR4vW7xYfAW7FCuVqNA2+Wwd
99fICR0UQEBaIGJ/Zu7vqrxhI+Ma9f/2e7STBbkOMTuYw69ig99E9wr8Uq4VzoGYWkdiEpPil+yg
17uknvbD2gkYnfkV9xctUsGuPJ/KcpQddQLEW2s/zICGpH55cPjFoPH+LErXDWnqJzPvw2VaZWDh
7dzwyzYR6Zw/6Bc+1slgc6yv+51XD9wp7T+sgWScl8NhHLhqLwqf5VCwZG0qH9A2PNMOuGib8gBA
Q9+7dt/q03nzQ/rymWNOY+/0Ykc9UN8UKT0QmKX/klWmTTQOFwZrkH2crfmeBoUpeebdEIGhuxZI
vw3uvFzWXDrSs8zNbZQjNZ/rAjG8lke+U4jn5m+QTiGsh0eEGPNBJAgHGfCtKqAmTkXTrR/fSbuo
tDQwaE8lAES2R376y3y8TUKEptgy5aOsn5Ssdo3lctsYbZ1J5g7yzGrvUjtG726Uw4tePXqh0Fg3
X8mTufMUfwojTPtal8xXtZSteIhYBipoXzf5MZiHEw5bx4bcgoFO6x6rDpYLl2trPH2qCaK6431V
jxQIobuqBV8d5BwrIFxif5gzVPC4HNQpIIKg6bgy/XFaZL3V6LjTJ8462WtLt7ZQaY0kh9MRILwY
fBPy9IymNkgz1GrHZydpJCZ5LfqUqxw+32GQ6iFGPHF0gjZULzvLUOsDHvzPhDNaH0s46fsIyQpv
spgeSoZY8uPBQes59VNqEUWv2+FvJejRoVLgM6KVzGTpuCYBh1rI7xO9rKUPFMeUGeNrvLEYso9W
uL9G1lX5d1ruwzTF0taNgH3MuIvl5vKUseQHf3zLZtIWYvRC3ijR1Ojjfe8blDiOCzoAOPWZbwSV
a+XMnSqoRbJm9iWDd7PfLrYv25rB6v2/b7Q4YwqSUnjzHwVCgtXH6zvjAmhCwBcdaWKXDeIddaEu
eW2gak4hIWjOg+QsjVm00hIlZNtH0MUHomI+7dad+Os/20an5kIL8dGTtZa6467RKAhp1hlCpXZt
WjrrGuSXwctRHdsP/3A+DQhF3kfnzxrDYKwzROIRBc5AIP11h6s4NSeR1XnenKBlE3udjGqL+pkp
dv1ayQyJ0VweeNKviDf3Pr8eBPoaV4eH4WiFmRbFwGmHsjIR8hz+6c3+A/WIdtWkhSpIFSTt9drB
iL0+YeXbLTBqbxRo0Pr08G1bMiR/tEp1t8eHcx/Dasn2wyIYyoBOBP9oZmAc24OCrNbZeOp/m8zY
jl/siEyjBSK+LMwxRnV1K7kyJBHFdXyRhpLly/k/8uVtYjWVs4zdj/WLvXwRmwgI1DXr5DNfNCN1
gdzxtSgb+P5Az+aNYKEUVX5jh0ZPZnhGfsW31QeDJBkdBUg+8p33tdO5SHKy24sDpJ86w8shNGw3
XoTVmrmTvQQUfh93BHk3W134uPBfC+lH4awIuIBEOEO45hiliQPwW04N3xOCJmQT+zs96btuODMg
n0eaXzpPtxkcAXHlQm6MB2/1g+NgUqUaG70f00WmMNSwJtAB5e4p7cQ6ZiuF275gHb4eBBtJ7RVs
9XIEQcE8oyThCgprHkyp4WQ133d7ht+44Up/EvzECYfqiTMwVhYKDAwaTquKlZtYXKnCe0YePY9R
SrWqt4mTNPdH55mv5rprdyeZwjOjljTl2gmcofZzC0xMgxuRxL7oTw5NQztK0ZW6ZLlPWeKOqXQO
5Jya1KdeYgtshsQJ8XvS7KvlShBW/ZhlimX5jGE7S3Caxtge6qHxtet+x+dzJ35QI1/1njzHwIYs
OcQBM841pmmEwwvOwcjw9SrluLWTxptJUWZhHdW9fsdS2jgxzPlUDtqCiS7v6BZmy8oni9Tli3Qr
/k4hzoqv6Y5uYpY1HyWiTqgvwoMxGFDSRNShroNQPZkrA3u2qxatTBCzcupRn4i/+6Gogcs9Pj7u
IOFctVF+CBj39I8WOxzeMdzvLvN2nMBJQAWN7jgToU6x/dHxKUhpgbxy8PnVUI0KccLVISu5XkBh
AWHknQvOXpYGv6N6RCwuRuWyI1Af7OQ6DdBstMGtmGWZqao8HE+PIwBgSdYgW3rCMqZPfshptTkw
qFK8gwCB2FL1sVjdUXiH/fIEo8QTs7H1Y+/yTaHQA4nkb2aFIO9dmC883614tm7BBaDWPSxKKu9a
TrEPb/N9zQjFWCFBFtW1G4FpFf2p1aBjeNXLInyIR0l2bDfotDAb9V2qD5NAQPM80cOfs94MofqQ
8OfjAy27T4QZRvTTPgok9fV3Gk/IsDgeb881AB+C5gnJ4YuTTC57ZfZgx/O4bTrfvnPHDizb0FWO
q/+QpsY3O6ppHTiRpx1dLcjPUAA4fNhyXTGVCb+VBPf5O12zQiaLiYXBQFOwPK5g4H4zbX+oaH8s
mxvr8ZhSaklErdZjT/nS4c/iYOj768qwRhsuptdn1uF654qkYCNS15/4tSXihbNjQpmZfA6Qg0eu
b/X7uoDgOCM0zl3DiNQSCPLycs23Bd+670Lohwx91oaqN7tU9ltzIfDTUhoZZXT2Rpwc+zGzgtwM
zqTC5UqhywZxhQwTLQoSqNzAs8n9zPAwqEbPgJsfTcMMp/Z7NSV3DyBgMiNkcVPqEof5FbaN9GON
mrW3rWIfCNw3xX2zK4R/VYL+oRv2xVvAgIs9jWhb7N1wEHizknfqoEnKYWFBPBzUXe8K/wk/LWwM
Jok8xHRM8IPtgG+U34U4fy0Gr2Uf8mjP+5jPqOb1nUG78RJY0RuDhSfmX2o4mD7e/IsapM9aUjMs
XTKmTxBH7lgpZcvmxxPrsL5r69rnlJ5lsnssmPKFjgw/dkTKqhdxNiCBNgi2DodfqLPcOEMZo7Cy
Ll63wTSJcP+v8+Vs76xhHJsGlCdQHGEV0ddJarI7YrlUsDGv7Xg6H7EmN1fsEvoiVLZ2agvk+lhD
EiECRFFvJSWJ316J/nbc/qWNLFKE7kLIktb4+qJf5u566Of8N3enudTCpXYg5F+ON8mHiOyw/LPo
nejZIjs2a2ObihllBtGLR+FuYMqRtGo14LozTJn9h+w2xWIAySwtrq/HLSjCOz/WY2M/u9zZmPXM
86SalALwZqNyFxVuPMINdsIkgvYkRV6b8knjh8wUflgDL1HexnYj5MDwdS3a1fWd1ErMjqZlYqmJ
prHiRZY+e5GJob6LnjmDwvxULnbPMqTslJnscc76fbGzKbbUVbglJq+ZO+mDnFbPKlxdXhNbSUuD
AKhcGrsYn4SmVYqJNOVtdBaWUlDsjgQ5IsHspEMJ4Jf0JXbvhBSDgcZYfnMTnCBDNl0oGfLJeOCF
Xp6X/rdz0TNTttpWezmfkXfv3TLHLsPAqXUahgxIoJJXhR23CRgIU1X39hOcuCYQib9Cqy836rJ0
hk989QuSILNfhr6jMSlG3I4ACsq8NphUV0P89jzx4uXVfuLPeVUbWctXRgaJkhXmY72lfL+Uz5WG
CCYc6FEnTlTyOfhOFEWMUNu32DD+IcYPUeTdc9HdN/q2JzJ+xAqsHmBxUfSbbcu1iNPxjV5w6qRf
dgL7PhNsdMwKUHg89tcD3inweVHcU4/5WReRV1CfjJ2qFvPUkFxSZsSGjNrTvVaLwLYYVUUFcapY
kNSKTVCmxMmBNQiouEWmq9Ze7cv+N5lEaJQg1e7Ls690X47UVYBYHFP/1ltnCpbn3nulVluLngh5
21+q4A0G8g1dpbKMmZUJ/OM2BSHBFMyk/6SqUIAWd8of7z+yZn+9+wskGphSQnc6Wa1PxvV0xyhO
Grl6oSYJmy8MG1RSbaamG369cBf0uW/YjKXN40EuLaP9fo6KB780hpspA89lkTRdkCs5h4TAHZ03
A5q5+PDLrhUVWUMSeCM5mqiBOLhnrv7hyRBSudm+7WoOO7Pzx+RDBfqg23rV+DJEIfuDp1dwN8Vh
mmbs1LWVnLYiJo+6dgcKGFAMJDi5ajn/8gwbD9guvKbDWsGxpUYmmqLS7rWfrF4uRTc/jxGs9tY7
YWGBhMfzYzHooXX+YIRo/ufMQQoj1dGFfndrXvrgtfHH2IeRgdgxxrB+7WZ1vNRPYvR0bS0frH6a
MMtExK47npgTZ3WO0A979NcECftjQ0C5ncFxSUZctLnIk8O9rpO+FDEAX/3+5wJ6FOdupYHQqmth
YE7Vsu43SXRK1pu6XEek+D0nQSiSCnh68F4FtO7yCzEqGu3NX7ZktOAzQK5MNI10IBWhVp95BW+0
hWPYR9yS6BTP3kZ6UVTQbnfA9kY3c/i06IomCg8TvIOlZ9SUfxKPgtzbDfTEMZ+qoPB4lcjuIWyr
kgpRjiTDKHADk13+4POAlNJFtr0oDEknpZdAU8v8gYiF4RyUuor+xmvYt4uxPzIZlDBHQyEHPsXG
r9nPtoZdD8zesbRZHRlYekM0OrZD+sPlLhVzsZdzO3snAhjvYeRYIges4fr6LGI8bOBtVz2ourVL
pA2WDWG7Fp+NwkVDi+6C4qMg064pLwvCr9G2rYRlq0klkkkr+qS0DHFZtXL0Gsb8X0SI1z1oH8qf
FvYtjKvv1mU5OSoPiHv0qGkPAavE2tNq0nIO84HnOTzYhvKpbeBXb/VHmCtg6StMGcc7iJDiNf29
NOqvjoVBahT7NEd6biA4DxEVfswXnwgeecH1zNn0ZTGE7BOJ8206Hsj7MngHVmj94gzoxg8W3qTH
dwnbx0i/XyzGUgc656PdTC89U+9dssy27XmhoWKlfkQs1DSu3pNFNvYJwtLWsWIGT67VmpUEG8+O
jgGPkqJJbyL5U+EcD4l2z8xoaoyr39/WbT953begHZiQd31qBQlxXHnvyqfwOsfYtwpCLoKqvKmt
zp7D4DQeGy+sk768fxtdyHY5kk2U9k8FAzx69SxFnKUU/ytP3NyNFOWa2ujBnzy8v9s+s20FtdXy
UthmfFEzmZh9zYnqO1wSd6sIoPjZkLznKhivFDj8xNnslTPt/8JXqlqonZdXCzCHNWN8TT3jlOS8
Fum4U3Dn9n4ETBLWDJb4PvorJemccB3hVRbUUJIMAtV/ivYlPaDY4+Qatz9OlPqfTtTny9Vxfbq7
0tycOIPQEcWnn63TSEONPrsrbuww5z30nshxEj030JU+PSkHkoCaPj8A6ouJ+GT2D1ktKI/aF4Ie
fbqxf7W59Yar2/pqo4MxeTalk9ADkjtKBANURRclQWokLRLI4RzK6OHfD3O0iUoPU17bt3Lxo6Cj
UVbZqhpxEzLyvMHBPkhWbH9YGpgKdb2Jb4kYhnhwlgFOShzISlpcSHKcdmrpmfFZr77Z2TA8Re/M
WmEDP65b0l3egiDZptLVHAF4TlpV4gVF+QuNzWPxWZ3leSEkUY6Hj2MpzQtGL05rYYyUBsvDYlny
SbaZdOA+Gy56TRmNPFCndJmnmuKR7g5QDM6rdMRChU495Y5LKEorrVDVISEFQ6f1Byd+CN74bwuB
NWG+F2w588vI4srL3WElFmksMwknL1e8zRtbWHRG/Y1JEQmU17nHVTj68SceCWJNjw5gKg6hIGBP
8tZFHS1tjxIIVBfOe6O3iEcqrPIyDyYSb6y3vNjRLxLqe4rpKjxbtIveN8NqV5m79J6DN3zoOJbP
6z4I6exnYKTwpXIFjtIuHOmiLGvxFs5Fg4j8QdC1og7GEWKbb5PnKLj36n6cpfArHSkrgFF7NOiO
JKLzpoisIKNl54o3dKr6+zm33042SP/gcj5iKEAD1ABjHmo9CKTbQh0aBZ5o8DpnLlwg9rGQrbYd
HGcpyFAp3y1ONZjTkHjI3WZuPisHSks1o3ivkL2/zifYyjtudpc4Qab3Tr0/kGavCKRwusawavFt
9sgqRuC2Iankp5vEFj7H35rBFdJVrNv9e5ywrycU6u480+EVZ4K+Y5fSxKOkQTJnJ6WBa3EZZVz7
NafVSPB4OF2/ERYbDeCqZ4/K4v+U7qgZUJ9Fs8prZj1xsRQbZkPLuTVD27wJnCsFncHEFfnQEJTN
Y9JedjCatdMu4hkL34Vi98FPTaRFi2IX9ZPmpCvVJ7wE2/ZcWCEx1ErD6/QJLh9/P0pZaR1XpvCy
3BwBBsNhQThggaq2IUITusbKWyc792VD8RfnT6VFwgJHMxTyCBBHX+6vnKW/eJ3EdPFhFxeUnqIb
RKtIHD1GnWNvZY9awMi1O4cN2hArUariZ6fEFVZr87MY96slm4IKVnSTOCJrHCpD1wPag+KAajH8
Y2E1MZGskXvPqI2Ednare2bWK5hGWIJYe23DlfWQBzi0rWbNQcwXQLG2+pH8f7ZeWiw7lzNVPrIB
N1YTBMNcYFD6poZ56RVDIpTQW7DRSZ2vURGKaKx2DQ0v/cLMy3eXsA8OUjvLhtHhjHn//M0MCnQd
Owj5YxvoZ1hor6TScYU+jmuTMGOLQalWQJNWnJpyNHXEAL76eoBxhwCYJHecSuljDDMIGIoS925z
4p+8y/TsnSdx5pqH9yHJ9BiUDasBw5tH2v3UR/47Cli88AMmNasiJ8QUrdSk2Efgmp5kX4w3kLuG
JbwfsFfUGX+4EHudTu6tqhIYzffmei66D0pI6+Wpr9pslz0es0ChRGXuqlshs4ssLyqutBT0RLmH
mZ9LuvTGq3kiTtlCC55tgFHKntUJAY6PG0pVH6xflPwS5WWZanTxOH8iOBzAyfzAN7py9PZY4P/a
EGluS0HIC+EU8uP5L8vYfAlUiMcq8xdcJetFDx01tPicqF5/pRU6609wjpWp7YW3GgZtj6fkSaNx
akD200zZbrmvJk/beRIRxHQSFkyWuTVZ24y2tJ8Nh33+Di7x2+5tFB2ql0DpK/0x2i234TJ4gYz9
q//LTQkqjqc+bxeXFHpY1XC1fZox4x+RFIOOhAjwCBtRQ6/5+yCe2KOA7uCGH17cxAoWkBXU4PUj
1kaiFRVWBHzKLUTm5MSZPOjQ8iv0vqVNj8zUhD3wnuWRvJhBQdwEYJ06lGLgievXQzzeIXMLHMgt
5ONxBgyj0C7t/fVW5MxrE1IUgFZxA/ikLSUv1yhNutyk4b1/AUZkwBo0ct5pQm20KvRMbp18LteE
Oke4AaQFoPv13IuWT5bD4nQVkoxWfLYBHbfnGuhY1jbRokEOqbvhB1iNBoLObnDyA4Y0TWnlIk7+
/DM60aI4xf4s2i7Ko2MN2Vy+pXr2YNUnQfjbVHDREnMNThGQDPQZb2ifhmt06srv9CtSceHiPy2I
U0Bkb9YquoHGPsEDPWUOufqLQN0A0wkXeBbUaSJDwgKuJuG+1lsenZP08HfQpupoQSxBWwvRpprX
hTVS3QynTw3szP0pNhwpPgAUrMtYl8eZjVDHzV0jPcQ+s0VCyjQbrZU96D2UMdeGRVcyOAjRBn1J
/W6GOBAGv6SWEJoqjHrXsSwpSmrYW+y8Gqy3t6ytN2ZQ+PWyykUBKbXLYVnsJnUtOcvID4/rsqgr
EDOSGeJcj+aq4IaoSTuIRr9+4kOK/CIhtvj+2j+bLwqNLokBRIVsJbOAty9w6LCCAXsGLH1OSsx9
hfRdAeNbxT/Wx5Oqs2DKEx6mTy8D+xzMEGJqOk2JwAEVodOaR2u4pTKvsP71UO0yWDOef+XWOtVv
c7s4+2DLnDidanbb2G2PyUxTUoL9OPKpW2LSbtT97cdxPcou0iAVdpbY4YSnqqV0NREcndhcYGmB
buhq/UlFGGZmYVnlKXwqWoRWD25ij3E9t/Qc8UMIZKjeTm2VpR+c9MIJYlQhPqBPu/jKy/LKL/9f
HxCFX8g2m/RnZo1e8aIKIRyyLaBdL3hNDW67nfZkcPM1gzx2KRlqjnW15w7dR8DwW+esF9VTkKTH
n2d/6CmoMbsSLbOa9V8vtmnuuz8brhzBDVqOC/RR1yqMiW5vV4/9a3dhDBEbKW3S9yD3YBbqxqjP
pnykkpIPQgbThBxULIC0UwsAT02jK7YulTSjT1WRvymsi6Rpks9aALDWDTnoY4qawNv5UWNWQb9+
bFza1Ri547nTUpSd07mrbKjOBHY9sp71GoSQTiQa2CasU6ZL2AdeHji1B4FQD6VW7/roPxiAqAyF
sgS41vIckRnMYRJ4MHcvjS79tkYcH4EtfD+iAcm4Qmjswk9F1R4QACkxzNZ23722aCFjP3Nkxe1q
KipZs4/QlBWzsrlpckZuY1Qe4V6I/pzlK1QuZRmmeVOoDabVD56t0k8He8/ZkSAh2woXLOi49n0q
fXB2g+77A1RD4qP3XBs2aVKuLG4G+UArDB/uF7LNYSeDVB+z03QSLCDiWyoj42kNJWPpfg7o2vrH
uNd1prjr+bpmVzSaIcI/watVGSC6ffrbVQZl8EaNVQOB3CqjxtP0F+k65VobsnAfgNhPl78QdcDW
58kwOT5mBUfGI1BaKPtrUv44FxDqP7gj4/2c02SdszblEkivxZuaCHMJCVMMybCYk8nQ+Nujw1s1
dbcIn029WFbuBuU0SfjC5HjjkLuoCDnElaiQZbiMIbVr9FQxlDwK3dFjkGP8kObmXoyb9329qF81
2fRBVfFWDzhQG+4FP5ENjlavmsJrXGwultEbiOwIomv/jjVREinqjxwfhKpBj4neXrFuU6XzYuR8
sb3428O5VZqHN/KIw7dpUtMtBvkvT6jr7iF6rfPXVdEOGA/x7Bo0qAItL79EOAJmbsSUwswTmxw6
PQCN9PUATHiK1R97auwWQNjpDOzLGicO5BpyNrpBHOczittr1ms4EVStg2s7NilBvE6llYkJWuiM
Kvt8SRkLYsVjXtOYS4A3Bk8B+IgBNdpPCa9CP9KXsWfARPgh6O1vZ6yIo171iBX7tHOnf6NzCpZS
jIBj6dMqoxjHAqFh522cTZkCsDeWGGo3oB4wGddWxfkx/BzHdsZIEgbZrJ5UATN325WIo3rLjH3d
9cr4PwDrIbekPsYbUcD7ylqCNN0qys095c7KM1hqaZMDq/xsPhAsZwvKeJ5ToyVCXOTWVPvOEsz0
2+0MUMhHQlw8E+8RlXBI+L2FL4H+MYwvuvIz7SniU7N6QoE8vcVtKg0oGJhdzm27C8MbXPPvw2dY
pUeBqMtT7D56yENgRhr6vQ30zQZqmCXVDUoCrBxuf0PG152M9Xbqvl8hJE294XHgBA3eRxbxCtNj
1GxJ7Y1b+rZAm3qpomGxGuxGdsjbABpNVNM6YF5TmG7sI115b6yDt+JOynK8+XA2y1b/VkYxVFhI
LBDrsh4c5gRAsWI0aMK3yi2fn4xigmhXWNpd/6RmRdzo0acSgQKxWF+tIprv646bm72I2q0uf6pV
Mz0sJ9Cz2hTWpHv21IL/HNXpfCK0CGNmFZrpUPJHEW0EbqXupjzyF+piADnjCfCq2iF5fJRSqQrL
rJSOEQ7m6JGwQM/CRzaWtTMdwP2Djz4DHIxiLHjadvIPR7N+ArATGxad1F/zL6+RLBKvBZYVHu71
IAEZcE+XUoZsdfNlWpunBO9zoDOBMTAi+Vs1XXaOYnnE27DZUNgJGa6q8BY+rcW72J/W3twVHLH8
iCg7JKWb9bPaeF0W3wB4T4HBER4HqhrFK4S4MJ+hoXDxddnAWmSj6iX+h157b7yAucxrbhmGCtT+
Ut890NYJPrLWj+ruA2jN/7UT35HSZXMNEkqe7AdJu8pwGEfmD9lvAIrkLEIvX6c0zKIvksLdafxh
jLdi6P5lKcvCQoMSJpWV/h5O7GF1vhqt4xexXV4xWwJdwlwQi2rt0YG9FBnsXCZfnTZKLwiwAJJl
E6TH2HLQl4vqzIRftnWQz2Jg5BHf+C+TuzbDW/zC8uyYsGdOFQYHFalQAtKndwVWoQi38ZdwZxUR
NUj1k3yhpxqlXtpx21YHySj91q0kBPX4AgXH2DtObR4Di6tfbwkwx9x7k2hAdQkCalOBpb4HED5B
N71cLaZvDfSYKWIBEEahAPMFLfh+xyp29aNNURgCDW2toXV4RfaTU611wqi+nXNDNH1QXYjsD7x/
U6JLFHw6JRQ+FU6u1sJmoxAuFtNY6Ttnq17xCcl76KLap5TVdApI1scUP83TkRRlsGMzUhi+f+01
Y+XE4LJ7XjrFMt/+T3Xl5BxUZD23ffHAS99WxT7UX1JaMINRyR1gxYdgrPnBj2GQhuHoQ1lHmzxi
tk4x8xs3YjhFznKf946X37l6+PpMA6AQnZgIv82HBKCe9sKb8ysPUYvEAdRQMn7eWoVjv/FFT6XY
qP7s/VDO2ufVfLhP8/jJC6JnnTKeQl+OA2oFcbdvr7yK2ywV79bQ1+Lny9CmAegIo9Qz5qgnUnnG
zrLslr0U0cCs8Qp3VAsMAyl0OouVP0Bit/+d4bYScRU5WmKAXVj0Esg3QQ87MkWeq5G3u4EwZ16t
L2+Dn1qhU+HsEsYdnUorKOTeU4oH6IRD4lKjKQg+Yk7COGiutmCyExcULr37oxyoyUido09jo4NP
RJFepue6TY5IXWQE9n8vXxL7pIWqlJhb915b41GnO179VYdABQ3Z+EYOqEmIMugxsq6SXAf0UYzr
FHBOCGK/kLEaiL25+RNAex7zoi43oEy2hkijP2e/7iT6hAPNPP6wNbp5alzTubRGuH231Mh43jax
ELsuTqijs8uEG6Zwey6+yrSn0/IfL5Z4sW8QER1zXYu8MqjD3eKiRSo2zPT5FnyUE+0bxMfZec0P
0WG8EcA0Gmc+GeLLgHJskRaMQMu9K75YaRQYnzRIpS1oUaICtZe0sIxFpoVc5Rs54829oYYl201K
x6Mq36scf76tJAN1aMbmrsmsNGYtUTv2ZLCpvO8XpPFnrn/5P9ahQ5Z3tlh60pV7tm7MAAYyuhzv
1Hqfg/shC9lXipQbOUq8ncc13KTZWr6uYNp5vdc+66x7h6p1urwH0NowIZRVQBnsvEbuGaPb5uGw
3PzHn8fR912zfNOjw4ZW/QQ0+c7MwyMiKj/Y3fwKjM//p+lIcSMKocmzEWxkWpUK4NWT9FvDtWT9
ecuu1DcPtH3oKZQCfOs84aSmEcsqPb+KLnRwTJrBX9FDLXkD+Z4xgqFXS5M3TjDTU5n6h76GodzL
xK+t/iW91qa0lOe9fYH1PqCl9FbuzaIqZFIsbAMPPazzbdeQhcaI9lVyzVuNeP8TBgIfafIegalh
yKt/ue4cK08MYcjCHr3Im4+aHq169FJ68DKygei8xZ6aO+rk0/tLofyx51gdLtL46k9sD9nWLMF7
VOROoOp7pwOsmT8EQekHvUZbL8pZQr3dACMg8OkgCfWU1rgrJpKZpnh5s3EwBFx2PjY1IJikYg6r
FBfRDw9TXAPzBZy3kEnXhE8tuLFvA8o/LP6/eoCq4HZLwGYj2+fzH3/ixb3Jb4py080Ii4OjVsEE
lxiiDJ56o/D/M+nmxDy64es5yMhxK5ErirpWgbbSsWypTrmUjH8MMK0gVIVTUg5sfVjxojasjv6S
3Oocm5lyjH+0pZOR5lxhqUe+pnReb6ioFRg1oKFljh4/tLzJOWdlY/kAutljnaPUSYlhV6HhgjOx
dmmC2JnDM/fQffSqJlCqHXZ7k5VSFQi8C/z2HRVpK4g3pKdMpV1aFUXSJ4CVUpjKVNInPXSych75
EsynaFjjBmYYiiCAmqsntk8oI02KugIJYvBDFiYjDvRuLUeA/BJ+CFFOIggEdauzPxcCf+JZklF4
9KpzA1iWJzCEbSgyUC4gLBNo0YKt5Kxw3AJW2F6Jfr+PQR/FFazqzhAQPPYnoSxuBMJ+Szmbtqed
MIcTy/AcCBbk7r7omcbGuFGxZWP01lK6avy5Hu8r2R/FAy9g/rUS2okm91/WmYmBOVoZrxSlrFrC
UNQye6pBfnQBLWE/EZQJNi27Js8T47frX1L7i2ElcunlPwMWZe0MmU/E3eOeBT5h/X8EKz7/gyCo
mgyG54pdxQOdrnHEI/wz5lNRVfo+mKPTyaJMwuLhoSZh3oUUK3kffJ5dg8QcgFt6QvvGTP0y6z+m
2gNSslt0LVcoKgEQ+9waXBU7QAJG0470z6OOgzJIq0/qbf7y+zDM9G8eNPDu2uW8ensrman2IdUE
Z1kkQwux2aXgjaOCXP5OwfV9ysWUjThjdKdea1L9DlVmamDHzhsyZyRYOyG4SbZjoX4iCNNGlIgT
UMp2VJbkCbZEE8SqWzNmdSAJGMBzcx9/mSgR/uW1KcWxa8t8ka55nCQ4S3jI92eMcz39hcBv/QaC
Jpm4vhpUksRMp8w6Z19v8BOlCCxh/UCNXCXixMnAZfmPkXiPW8LDHqgMIfwl0id5Fh3pbcP/0p41
g24dDBzXkYxjXm9Ys/RI00XtYiaRdIBJ1H5C6FaWOaAGQPB3ACMvi6LT+d6EU8B3pfyiKx6G6J+t
dOXFGrAtu5nrWtDwdt++784zcYUf9clokiSTSFgvg9PFkm4+JIyehmAx3nuhi8FXF0grfLHP3mrI
ntTgm4UP2ISTjzvJzo5MjLlLjmiuNueCoTyXZMlhWNWv9ftw9eO0z99C+cZ9SpvFQoLZoO6e7w1N
VX8Yr49zg7XSVY7M8CEzUd0zMbtYwavwealxxZ9uoeWvjQeKKPguosUVDypYkg/lJ3/0kesRkbVX
EMXZbCEVEhgkcYbw7rFCtv3KC60zyCjPRhP6Y7c7asoGOOUL+JC66uqzD2zpnJxrIABVH0zBAaU8
cToaPP3rAwPSPb6H0uU9eKS4mRC+JT3hqJ0eh2b5LOurwNS40U1OvrRmJlDh4WwDx9YrV8G9AsA0
rKuIOkm5R1Au9FwYoJ9zDw+Ph9fKBSpf42dvfTUKlCghT7X9GX3cYs8bjGV9ictNh+LkxOeP/i49
VWiUKSE7SF++6Xu3TTxT2rExmGE9WlYj6lO5tLxQvFp2JV1c4ssnJLRUZORSe9DJPW4RETcvOKR/
oxPtIP8BF21ozGmsugwbOrd6AbsZj8apDVdjR+9axoPFpv3d5T1hA+c0OIDHKLJOMzTGKDShj2R4
do+4mJBDQDa+dOS+70dERbgVvqQ2GhYaAGOoIJm2C0h2WvElKBYi3adSVQn/6o3ZIRqZ5sDZY7xk
JmQ1zGCHVGc4UyDVDiRvGzMF0mT2HbTFfZgFGRje1v2aFbtc62R5O+70pB+hZfR4hrLWpQu3MO5R
ALO6sggAGtWhFF4N9p/rKqYDPutrB0k1ThP/fY6G9INUY8TsyNRH+jFKAOGtieqT+9kwVzhckdnW
1qmJxptFAmfab2g8eLM2beVdCuQqVuied4n1OCD0jWm7mCx+B40wAAmYERV+Mmrh2vAXCkKLJxP6
Ufs1OKyQIDRuiuFCUDKLIU8OaxAqYcwyekA7MptKda9TAsFP46TGG0eAN6keTV98KUn4IkPlCZZ+
lRsB/VJGU8QS7s+qf4w7IjRpRUxR+mqwV5lyvnC+jkD1voHDejPwwfBTkPK67pRqJ9euazdEHIuR
fAQ+56s1pbnyKBQYxamxLBSqOkqQcrx+ZLV96EPHNEYEYKY28vQGZwJn2VheX3V96D8kuwZbFWah
JrCnWvjdBh0jgEpg23Q8alc3YL5ymvWc8a6EB0qV/XpCwK2f+ZzFG8ep66fSLYa5phfFCtgiyDZI
2d6xbbT84k3JXk+1X0vF2WBkhlgdUnjF3X++BduaBaXU2S7QPMrQbM+pGLdlKmbwrnU6H0/jl2Du
hWGSgW8CvRbipAHwG+yT0LlUyRpZPycD/kymdJI6r80s1ZKiWZ8Rtm6am4KHDvUAobwRCmP0G/sJ
0/OwHhZ59GCvh0fWSGWLktsalNzvN/p8XeGLtdbHYFxALIym5fHPZsgxNoF0kxmdlf0JbfBsPDEI
JXvN9gHVQXUxPiiPbDx/1O3uF11O0N4wGqgzr0gZFqiASMPWrIZbU1RUzOvCFxd9jr0KdcW5g4Ca
z2X8fSuCvAtVfmtrlWYKzS1MIhScWOt7QUhUXS4759YM8S/XgUiNn9y4yIRfVj5/mwnz6IjYL+W/
WLypn8e0Pvn65gFmNqHPQ41mNPiAe7FytlRAPmpA0uxsdsj3NhYALfKJIo8AxfDGa2DFBy9kRpP0
rNQuZTk/rd+XLE0Jit74USr32oKEkEf6qvsukY1asnKYevo03TzAPofarj74ONCXC5pin5g5XiFq
VSBP/5TcQSotzZ7iqbNRnHDFxL2400INj85banEVxOqAQW4aixji55Pv56zR9/XS8PjsmWGY8Ryz
4z+N68UsvMN5vUlbR6yIjyT99TTvkRicLH2MYxbq5lFaYYG6ue+e7fWmUJZ7rse4A1urLXhZiC6J
+cZIsunjXOHG6SlBcQFSRDpLldQIZYE2THD8rMS11tlHZ8p8yzbG5G/pVSHd/20vAHNhxoYvRHVy
CjCvW5NsM3ZmKODMgDs2Q69yZRH2+HgHf6PfjHMUBa4pfzl//H61d1JL3rLfdaE+eWZUiQ/bh25c
KhcBaHIbJJLnq6xwnRi9cKZW1TN4p5nRJOLg+xHKDRAboIawK5sFOElKTFLMZiAMap12uNlBwbUL
5/DdecepBW9XRv96ohbsJb72EHxQwY40w3wqo8jzxW9PxMZzvDAGAfs4DGy6TDoc3y6RiDPMZqx9
y5FKcy1e8gb3fvpaZO0yPa2eAozOspA4gFSQ/VQW/jlq4lpgYTUvk1nsZGdkgBrzFPVOlolwYveA
rdUv+9xBMiidz/oSAeFBWyc+ulfKm+wiRBX5QDpm17n7zC1OWSXph4FrwuZV8lp6wXuJy7V79CpO
Ch0iRR68UPqNUhrhpzphph5INWH+CkqrmblTIi77xUISgzbi3Qq6l0MHIlV/FwmeT6ye+BKalr4k
4/d40PYsFlLgHkQ3qy41n3gJbnM6jWw4fmbXxrKMLynMPY2nsxfLpECSb6CzzoIMobOfVWW//fDq
mNMbS6jKgDUVWGDRQ6fG38poP469g3GWYlrbNbpL5haAEXMS17oqhR/xXltVt4MG+0MGlIfs2hq/
FNZHZf01pys6fRVuvffdvPuTNXz/XJP7iwJUtS+LRuIXylRuwWBCbsh92f/cQgaDHGdtSW2We71q
IyV2p89hZhU5HmMUGguMJCAOS0riVQKdHkCoeXOLkHMAofUpgy19/1ahtKhjgS+lmiIraS/bgzjr
hKeK9dieV1FEM9+7kZoN6sLxUbXN7Wa7HEobmy1Ooe2YDsvq624Sy5SVUq9NjQxthcqpVBXcmj6Z
UqYZmjUpiX8PNtWhYcgLbpX3YoJEwYzaRXQcA6fF/zjN1QiHblpeVIDIYA3SqRKW0iwtiwmbiHkB
LmOOOt9tQGqRvesUV5/OoiZyMef3Z8ceWtRg5Gj+EzlGtsQn+IufVZ+NhGLAXmZ7MVtURmTves/w
LVr4UhyLu5yRduNFbrGUFDymZibCHb+iA2tL1AWQ9yV/izQNCK8516TPdhOvajuvFAX/SS/AR+ce
HR6QNkhqktZ+Q93+pzQe/J4kc7wLl+zePtwc0YEUhLg7flIBINo0f3p50mH4rqia6VsiCD0Hk9Rw
6oeVLa862UWvc3NZdBvFT/E7OqoIXe083Zj+9JHdBEvjkgz+F9HeEKIAJGHACHj6TaySOuq3xShT
Kn0qATimuYsfU5d5nm/nxI0NsRiM4UkBurHrc1X7WDNtNF671Ak2M/4YMdxduva+XhWuVAM/QFRd
tm0XtHpPz8fn7Ot+yivlH2fpmqw1egA8CSRQzw2B2/Le2QwbpbixJUJaiMa5ljVaa2Fj/h54q4sg
tYdhBsQXB73U/85r5KZZRLAsKDXUErX4iUXg/3oGBUxw9OZi8kQvggtYcFG/Zgu+XA5LzheOXnVJ
3K/H+doV27matDmhYhPimTVxx1+KohISciU9tRRwmvv7XdeqPFZYKl/MDGV/dPId35KNdmo73UWV
S/8Pecv6CcqE+8CW4lu5p+GI0dY5nM3DFXrn8nW5lbk6DGBZEr7ilyck/suwXEd9l2bBSzP3eGa3
nD5rtSq8PQgXRqCBLuFFd3FOyYE8DFUnhCUhZzZfZ+ldtVi57oH13R/1mUTSneVvMnUV+N/dL9JB
J9+3eSyutB1EYOCjJs6LIVd8xvV/okb3D9925hZe4TXc5OOnCrR04q62a8RgwtlVqmNsU4ip1cFF
54Dh+Z1Gc2PVOzxpusxAGQbWYrZXUGGGTopLVPrKhcVlkPX3pKch9DOV1NSKVCqwY/3NFdyVDUqa
DH7LPN9EWshQlngygtEDbQd4W5n1vG+nxT2kDVhr152tBpbsyb3fsL2kRQr82Rz8ZPCtq+WcBBQY
ziOl3nmsoa5uFAK9GhdbQrwVCc3i8lIvZiNG9o7/RR9BUih+7HY1b57BPnYL+Dc3v6GPvPbiBpqY
DvuOQjBuqph8H9MBSzZ2Xmy54Wr1EFX4X8ZYblFE28XCTF72U3wgTEkoNuHC+42rVztNMnEYOAU/
+SaP1Pw4JzDG/DiC4cE4UjL2TPGY7e1aUC6VyUmepMafv5NRciWtskUFuTd99gaPKSfMJIajRdlV
1T7cb53YhFQwpAXlff3Mx6KpySaOwfpQ4lwXOvWORZdEiD2tOd2DU0j6Lsz8JXh3h426HHSKHFNM
LwYH/WEwlPXQedknOt/c9gUG+XKjClkhRwC6YUbv/kwSl0AspqXpSrpsMrgjEtqekH6cyUIMgfHX
975zgM1U3+OpYJ0upG6qx8hcUJxgMdAoDfYeAJhIrHonZ+GOVqRixXLqPbt+bd4kZZsWJk4tizYX
gPALFPWTuJMNaOGvTnUvQi97nRGBCCFTKlDYY5wKodr1qNkSiqO5QfiIoPEf+p8qFrCgjYB9Sklj
upReiDxkEq4y5gpI278DFaue/LC+y6Mx0KG97UUKptTf9Umto6QsfL5a+vsL3Jz4eBSThVGuV48A
hf2Wt8tj82zhzAP+kKJnU6Cgx2vkhHhT0Mikx+ZlaiP1m1aiiJYS0FWv/Rm58Pgknh8po+/eIFPY
FL8IuvGGabtpjUgE3MCzmnDmXccEaWFPuvvMbNsKaerg3ued6ospHUeQSq0oty/1q6k/tJ+dedj9
XHR3xIcSNqod2y3V+35oFpgMwG0MfbIK210Kw1TKPAZkzajSQwsQl4cgJAsK332Afcr8KEs0/ArW
JqQzlyKtEw4RuZdZlt3uRSEIj5j2XlVLAfutTrRnL/Z3//vEdITWvZru1CrAQaAbrqQOi3dB8GtT
ec43GPUIfWV5f7jYb7wwLBWwfPuvvCDcCzQQQr0FB3oddEMmT7ZwdhUbX2mqEBSxfuVRaoGAYPUK
72vEC+UxhqyXAfbMKs4FQHhF1434x+gUQKvrhJrgY2q9pxBEThfMW84BhZF11njoZsSRvTuxXtqO
kcykz6P34VYWaPTYolcVYgkmP2XJG7bsCHwydrH3VXrkYmLr4M+IiUiRkohpfzc3F6K8v8utX93Q
2mvvTbLDJRIp6XaIdx2pUQO04SpNWDTvank1ctapdb6VRb6FbL2XkLz3atcAKedoh+v2a5p2c4fn
AEVjxpE/qgqIZumrr7qrlYG00PD3vFEN4DH5bq6JoYSGSr8+4RUYICbqcXdWURXkpRCoKqWpGSfw
M0lL9tkTDi5wbV0xp1mIWEcRZnzFwpnkk9SO7Gun6BBaR3CbhOaBJYzJryOR0Er5bxp3k8CHownQ
oXb7JZvCgRwQtnMvkHDd0f04We1DbguARhS7POsd3H/oBMfCtQkw1eWSss0RQOO1Az3Lxf7dPxOu
CJ1SxafljKQg9KsdgDPuGeylwoSeLBYUMt5jAkch1bJcOEKnQo7VoFkDZvJUemz8OpCBhKneFDoI
Bg53EsmuMv9W+Q+Aw2oo8sxAfLHXxLZrZr6fUS+BWq91g2Pzo3FR2dQheNbfAe36k3DLSsAhmXR5
9TX9Vg+RuxMnkqFmbmkemC9oLVLDV1GjrXKtBO2+mjVgrm3dCXExHqgW/3Ec13m+RfkJg3umRmxs
q1FFKLLcRa2TROqP0IiPhGzEOqB4NwlIPg230EIPqWAJC8CyfLYO6DxWbn/BNnKwTXG2Cwri+jRd
UwqIDFWU1Cl9KwELnr7u6tRU75KP2NiyY6DKPFyiiHscRgzYGS4xNY3lw1wGkc66j2Gu+cbsDbdQ
J4A01y2S+wQ3CuWbeH0P2nayey+eKHhii11V7JXcznv+VxhS8mi5GfmxPYa0QKMvZ9gsh6hYjm8y
/CxeAiL4eIi0LAOdil92v3ZTzxNfoIgImD1tVC2YepxxdfY1PWKdRcAqGZwl0UHWZm7O+8qU+ugj
d4mn0ikGyE1SkdpuTG1HjIdrlqL0W8LBN6IJ36+RTjONX/ffbNj2oUxl2nViwor6lHrBkEgYGZ+y
h7S5BlgBBb1n7XUfSJXWvgvNzBLbrp9ad98b/o4rGobTwTthQEf2o2QPuV6JGUUrx73Tm/wUbWlA
olx2mR9bL1MLF4OO0VCXZHpGc6sV6Ii2v3X406ACkQrBnbhUSmHwDpgqf7LNUbEIwfcIs3FVt8AC
y8nBNqZYmhWapkeqNNZeWztVly1fELuaklJgfT57j4GZ+/8NoUMEA5iu47tdFClH2ZMYYQtU8gsv
UNb/4bzKW99oU6oFUb5Sx8uWjiaU32RK2wPi1kh4+2flxqLj8DtNr8E8zjA9U1KZEZfmBWIq+m6P
s5/AxcWwalcMwuEQ3O8mK2l7b1YkS8//8DmxMHYK/1XmcZ9Wb8hB/y0sDrL3o01PIkCOO8JGianj
9+zt551SnCRsHSXMROoZwPhvSK9JNezWe5OUEYGPOubmrHzrAbaPV7hScumYr6YN7X3qWteX2gmh
4cH9wNpl3HEdKoMelCfA5PuTCu+spQWkVkj/SJ7bUEKLViecVUbWkBBJmpKTTuKewSSPvjjsy9qt
U+pradfEjVgKQmfcQev/iZjogr53QJHAsX4OZWQlgKo41DiPBXRJbwp8ppu8TLbSVl2wBA/S2nxD
O4pqiPWISVGn7eqa6A1uSQ2fjIoiHJDvIZ+y3f5IZqkv7RpD+eGiz/87cbuiLlkCHlp1eFNmO/Ok
N4Fw/0P07fRvbEp4HiY9QvG0Qk7lzP0uuxDBxbss6NWtE+xubJKryRqKPOrIkEmPvwRxvP7TxB6b
jv8bFdOumqRnS+03By6N1IoDI67GBpeDBxLTDMmwkgRxtzBXQY6t9PMSngnYE1RKFrjOsVK1pC8d
6gkIBr3T88siMMBB4BZ2gSrGYn0GpW7B9U1QRtkLupsvR5L6TfFhvodFL9yGyYTP2bx5sB/zv8hM
K2EeirBBBwx+DpG+/O5WW8Oav9GrZzGrfISg8e6xJwh0Cpqk8xpHXWob1XgLTppzsZqugKHvnMZC
c1oTDWBXTXovF+hXljvi102XNe454MJcKvp3wlu2b1eivB/DHN3SBiwYxsUHsqV0CYlY9DaZE3z3
twsFtax+p/3ItWfl2dCF/PLbJk1nXH5n5MGkY0ukcNiuMoYK3dv1FnaJJi+v4yS0E2WNkyNTCo1Z
4a8M6Y0mzDN5Vqs8WuoKPlcjv7/1noipjsaBfd0DMGh9b3TCSZA52o04R0z+2qeqTU6/JehsakPv
4Zve/Zop1qc8V5ydcJUXOhjY8mddqGjT2CEtqznpCp30E7pu/reLmaHCxi8axMNFWJjFk7dYxO7r
muF4U/AoAlehqg4XBmkg5p4B2fh8B4EnZZUp0SNrgHm3GB5WJRU/a0o8HNlgmv5vQX9oYTXCQ9t7
DkkqnjAFhNU08md1d/Fl6zUqpyTxuP9Jp/ndxmHahqOLevuG8RiJCypSoK3ltmmPj3jBu8e6gkOo
kYDUhEBuDl195mm/Z87cN6axtJqKe7nCfO5LisIiQUMCQrcB0X/iaRkBhAUjGV2MtXCqIFrWyW6o
7v6qH0i32Gg+vxKwyzBs/9dvIq9/zJS0CirYKSyh2sQXNx2dAECcXqFhgmF44bZaB2GmPC8rusZ+
KfT9zR6lbZ62Zrrfp1m6gJdqKAxnaAHwUYffLD6Pds/0McSv7j+ovVwDsYGhWmN8vK5ExbztqHpk
EvDcChDjetx5O0FcFg+wBUw4O32Iw1OePUVwdTgpBcYqrHPQCK+tmEDa9QiIgUKASGldhf0d6N62
KVh56S7LQArvAT9rNRaEnOdL9kVvCxPvej+gkV/pDVsVvK68CNl8lhRUJl/fXOzb8awDfvnhAS1d
QtMnt7cJ4EwMITi8AF68iX3OUBkuVNtjXQdm2f377d+uaBGAYupmwnHvq/wkg3H5JHEFMmRsAeIY
/QYo+HM12kDHGHDF/ZUlN9JQBtIxlWbmI5GyTMpfrHMlsT78HPWrGiB/JCmFaiQfJMi3/S0151vq
k/0p6Qsqngb//t/cpRvbk3qMnCugEjNX7dTjdYhTqnzFRcLHuewn8QMiTXBjXkwdhVcfSVC/BtCO
G5bO0hiumgSvtVLGa7AtzNAi+Mkl3R+DXIvqlbNS7LDgsmRrS8h/kYiB6gTo+ObXf0s3wSkEafOB
6CDLyV0v0ZNZga2z9mphL1iBVQNFSsAl/6z3yMtK89gEu0Ftg+WDL2DB/x0uI3Mof9GO1yZ3YKG7
ODGZIEWM3B+RLZrnd+/gW+80c1JCyaSCs70kJEyq/4pfZe0hKeA7sFZ1BJypd+jNqlKHeieIbxMs
bsanaBW89VKSiLbbQCp6ZnBCHxoyymCgGPFH7FgdlnEYW1EEc1hJ4vKKdQaTF+4nLUij/hPyaw3P
6Jr3hE+Kcx/k6xoOzVewQQ4/l1NbOdb/4YvEIgae8ZO/SgP5/ElXqh3+GwCKMs/v6w3hUwrFLf1B
0u/bS2W5AJb+Qu8Is3Wv4xPTIvLRdKgylFP25dVQlu50r4cPXdMcxylIWhnyrOL8jb+j5RfJOK6F
Iv52JFPg5fpHj1fI64WGidvLFkYWAq0NAN9eRbKTsV5eU4KusANL0OgXHrI+1E6N+fBRBi9w7CMG
zEtQriCexu0n7Arh0kxAOOqFWB+bN5dSL4dB8G5H223H5Z8qdhVxclyuYJxyrJOVH+LOIjOOzECe
axSfqHwa2GvYSg5GBLgz+798lJ7s31Aa94QfghEgEzLXhqhy3Sj5l5qkajqWCFMrAwXN3uY78Npx
Z8RAwxRkxr7gqcBNypVQJnrbY6eMePajsjKfatZ474SNIyWA3I/arsc1gF7TtzwbLYewbC2uW6H9
21UoCaF/nZavwtJt4AvDN4qAPl0NVgxp0R6HYiTsQ27e57xeSEemnm0NhucySu3ZD/1OcF7BfHwI
13tcWAMdivcgWj3wGMUKgWAt4NOKIwryBiFiXTyGx+hQ+NZvFjiD0vy7gMq7VpqCZkBzHEbYEgPO
ztvGdbHEGG/+or2kcKITdRgaB/++g1Zd8FMYYqrkGgF8/QxbdVo0xL6Qk9Qbs5pfI2RKHAEO2kfI
p5hLfTVxvBCpy0hx95MX/fMA5mcP6fzjzL/Le3WZM9hLx0xXBN4ymwBbSWgcm4eDMPqDmgYl6soZ
7SUW8P2mHeqvFmGOr3X2uHndy/GyETs9hrWA2XPR7rekosUCdBqPZ2PBAB+QJKqd2xT7y8vd1O/w
H+FPqm2ACIIqjyGjDl/lAdM+YaiijmWyewNgAQC7a4SWunfckIp0Mwg0pjw1UVKtPYrje4wDs8Km
lIjq58x7i8UYW4dp9d/Xn6uMXif0/fYjTCHIcoNpNcXodMxn2GZFoVwlwNktu/9fcFLR5JedDts9
la6doxUk3DOFnDabLswhwnMyWvUV0fudqsf8TdChfGv6so0zvqpIK5Hgi9k8zVnL4MtfrA68BVzf
s69eUGtYU3HKVldTkRio8t3SrL2uGEf3CQcf5yRaj0lqOn0Qa881txgw1CqLUUN0/8pNHO2rQA+i
7d3SVMJu/PuSMNj2kZYNnwhcaU5klBzknxUijsYVhuGKqIm8uCkdeiPJJRn1Z+wd0xVB5kSbZMwi
bXkzuGv2XtEmyxyyZpcSTRgBsKNJll1ulQyNxu6L3vTa17iAJ2le+SOGoJjp83YHSbqZuwLJ5g6b
2l5PL0QeBIpInkVF3f0are+Rnvisl6Azdj7aSStcA4uAW460lWy6KXJ6MhFMFN34DzZWAN43YvVl
mIN2xmu+VmvIbTQbG6kwgcIX9+Qpv08PAUbNRc3MBVbpSennzP+zkkOeI+20L5baJiRQ2I9sXnpl
zOEIqJYL2bU4LH1ly+UL+dW70bUcaMAEA7vLYEWGQqBaratoXODmkQZHTYLm8wdO3gJddDEjDPzv
ShZA73EVZIIghD+5hn40rRGzdcPIYoeDS6oIQk3WdkAuroVG+XWJ0FLnrU1D/ouGOa+13Xym2pYx
k9AbDwb5Nd2tzBm21weuzI0/3okBpZQtEYDWr1zDTQbUOOqXu3mRnygTZl48GHzOIuhaM2a1mZeS
nd5KSFmZf7M1rGeXxKa93WSWqjvNQjxLz2xwzXonSGbVRn6lZW9ONMRT3y1TTy2FTZ7WxdzJidU8
Y4nSyVTiah3DGbn1dHgAQxLdrrPZlZMg+qdei+DCTQUea+tQV1wf5XRg+NPoaSfxB13BBHE6iHDe
CuJQ36L35ET14e/9VMQ4OJkV6XtUOd61hURPUPrdZsHZEx5+WZFLrAxUkL+u9DPAy4e1vP1fbmZU
21hXouOf01IGqomhIizEqYq6z/wy0d4hPL2N2BhjlXY/TrOSy52fclQzNvGUullayn+K86PLSjH7
65nuGZbaFhY5Y4bhh+OanDoMAY+zjaYFKaH9l9rwaGLOp4KsTW3BBuERfffG/7+9gLt275u26wlh
FdBaeiIjUrbNMEDw2TdLoGbXSi7MTfJ0DLm0KXggSC+qjpd6hmdiXkWoEA7Z+LZZHzvPCj8Jui6L
B2Oje9D7JpucCD/yD+IqerypxZccznBdUZlKrdsmb8kkCXSoQjb7yBdWUv4u3RHSqay4ATRQeFXT
5Do3weQH0ka0SINT7x3bHZZ44uNKUKOfzrw7AeUsC0o9sIhMFEAZu3HwLgJHFBtgalPPVlB8uCJA
6+cWqQHI+ieOYFlKlLANhwsP7ZChxgRESFh9OWphzTEC1ZLW116Z7ot8rlioN8LBNjaP4DTBjqqY
Uchto9tThmU8ssITMAyZxAchnMv6WVvbgLdT4Z2pHskaiK7yqy+On3h8Cttm5BcBIPuuvsCrXFgR
oYiLAh9kJJSH5LNIv2NkHtoRb9JbtmH2iUj3zwl3VtakEX0dqh3TT9mbSA9xItbUCIohuh6RM0en
olUqrphAMaGIzIxxqdj/sGNgTcDRiAF8XQyq9mcb1EUy0uMNCLslZdOEJ4ldWeAWjNS8h5q3KoCC
12l7znZULAfqqFeNB/U/l2Cti32BoVpFLU8cRvaHHw1waUP7efVAXlYJxm18FKe+AiD6F+7R7D2O
U0Riwb7pId+/2lcDUfCjaenwmi8J95v3uQfcWmO9QKkg9rS2ppxJpmdnDCpi2P0V1X0vZ7hLJShu
QjABUGyPh7zu6lGL4kUHEkjZC+tfhiXoO+5mjqdPIBneAykc4jsmJ9UmdHql+caT0SQVh6MsttCn
h7sku1p3XQyxkOoDkGU3jjokpeArHZa6+NF+nmwOcJmva7Zw2fE9B1APqZPrVRUWsO9qyXUeBiSO
t6HkFoZ31KkOCdzLSJLIN5BJahvj5Y8IEi3mND3QIH0MJ4E6MvU9RiBYfx5zM5m65HfcoiAQL5US
CzPw0b+DFpZp1twyEa2xlun5Jz63kC8v0mmcXMfvEAzShq5GyREAbLFdW5usnUltwbypR4PeIo+P
kwWPLEA/BVIJQL89FnWEhm7Dqotx/IGnX7b6JjH9mRNmYJjDFcFEjnHRrxkPwT+pNtvwI/L1u7BN
T4wH6ZXxa2rmeyHwkbFXUUr11SCNKJougYn1wIHO/hWOHMXOUli8DXlk7sbLnYgE8kks9AyXSLFI
oavlvT0Itv87GaF+zEsSr4cr9YsmBbmSOxejDCaDUCJZ5T9we865TRzcEX9ZIFVFfWfti5qvTPVY
lbIhzMuL1U6Nt1PoNYfaltTbR1pvwO3wMVrxLEx9J7hxQ7aESu5kDRXYo843so9jLdxCxXWY1Vce
zI4Pft0kJ6xFeLxZbFRDq1Y6ZN1jZ7nx6ZUJMkmDsrxTsx6MtTQ5UP0up4OZ3jA3F5btpZQvKoaF
MDrmGLgZs6UO/0G5oUGoXnb7ArkoaBmMJ5PpsoFfAQlsWgVkF6hQLxgOiIO/1jw122PXW9d3Vb1P
Q/Tpz6UmgtgTYUN4i/vzwZHh4Y623s0eM7xFXjeReYuSbEM2E98WPFGrorMq9bqqiZPDs2CmzSVW
HBcM8N70OxJnL7fWltVaIkwcKLRbqfja5g9nAXeCWvpk42CTtiMNSarzXHZ0udsH3feqRA1WXLwK
KEGeDPoTpb5lUKmMwuQNOYHsN+uO6yMEgz9Y0lSf2Tgg4QOPTmj4ovY8b8QXivQDJZsYRG2c0vaa
5vTQbeIG0vuuDLUCpYFw9+UPo+6J8Ys4Fbk67oBpgeUuTzcpCqq1z4ZaS1B37M8FOzOQXh+0IyKi
a35Of9RUVW3wd+jLdjJsT6VYZh8hzhHjCoLKVdKWoxmycVzexNs1gj7usG2CpOc8Zs3GBQh521oB
bWH+mjOs3wH4SbrJzJ7ZK9F7ufUyLSCafHC51kJFCqwctMKZW0PuyACLAnKDQ0h10dqvSI8LshfF
zUldgmLpRerW8voNpmqGluo/LA5ZUyR+uPGeNFFjYX5o/4fHHarlF5KgcVo08E7HH0ltNSGdfcpP
qvw31yYUA8K7SJNAc4BrJw66XdSzuJU2cIpwGStpm+jFipkCbNP27M0+Hq7L2UrsyYKlZa+vKRPh
F92kRza/stUGHD82p0ERpG3fAd0tsza03SGCpQRl3r1Ur1GR1kt2YwG7TgW09JmKZDbV/kClOhVS
sQMTXvB2Ofdg3aQjU6Q1rFl4Vs6pT6/iQCc808X6VGW7vb3QdH6dnyji6gaXdUqwVrJ0i5vaAUHX
S3PHYY+6ahSqUSqyKBViTuFMB7qK4rwZ2Ne2b7bKL0tHuivNIF1MIJnkRtsjWh6ILdMCbwJCSdjC
ZnKC+Ztu62bteMW/+zblUsRCGt0jn81/AIdsCLpV2jwsx/MnZXlNflBq8ZQLQq3QnUuHIukKYP+t
Ea/xwawXnwK0/K1t0rDBz33mz7A4aDbhQcrAYxX9WCTJCbEvYJc9x68QNODiQuKRP9dme0TrQi5Q
QAjWVTMXhFChzLshy4IW10HaNdBOkxFKjRWRlwA4KRboXGBV20DbfWAbOHU8I45agTikxf3c69Cn
9pgwX3O8IdNjD6ojmySlzxD5hnImKpsKvpWbqdnP5vdM5JD6Gxaoz3fN2XspCxy7ALyGkphEIMlU
+jnJxXtScDrP6uN1I0GpEhB+2HVaVUohBvKCRubaA9uWPXfmPFe2DLeh8V7BGma29KhIcg7z5M+d
UwWKqsFBDVvpCsgszwYNIZNB/EMwkipbwXlToxBi6wMfJw/IbxL/StHbJFDEtUc26VngKZrxplyI
i8mDKk8j4aOilzYwJWpxnhGd+HFu9DP8fxEjp9SW7yWdyuzuxe08cyjOXm7vK1X02HWt8/vKgoTQ
9bqFVfVr8L9/IE0nMrvzbcubD/x7Hj4120iRqE3W93jkGxPlpa9V+cJoq74i8T47CELhbAR0fT8p
/yvaQ/ma9ZoECKmF/R23AIzFBEtpULlhKNLApb2ADpjToXihLlFCWh1u5ESoyqob4YWSjlQi/WyI
BIx4o2FXPvaCwU0pfaclqfSXOUnnPgIvsvilOJ17r9iGdsaUTq/xiQ6bB/19BK8wfcfmgZXKjoZh
SjDRE5SVZVw5UtP8aEjWAReGeBxInUQ4p5j9p1v4SAWrS0YHzYMsAYQ5xqZFHplxcyl522FeWfee
z3/db5O947qv1jpkDWC9eI8o98SiZ/UuvUWUZ0YAkMg5TKzj1ZPeVq9xIZlI/ax/Ukwmgl3lPUGS
zTzcXfZVKxhqRgkKLr/ltH8F7ShJJ3a9yyNXHDp7hrhVJ6FzllBz4nKE3Ijt8+ob8ADyqq1dBaUb
9S1l17oBz07b43Si5ZaogDHn/BXAYUe9AKmi18UCuGu5p9gd3uMb70u35QZTUl/oh19JG5sjE/tC
0IaGaCFDg3mWCM4TDUKnUuWKaabVDxi8ucwGBQE/l/5VD8ZGIy5fJJBRlHXGUxH1CgHES+CyHtUO
rD1l7u7QpJAxiXpy3eBMeOoXN9z46zSWO08cgRCrMcl8n2VvgnyFDf/eXqnoe/ffQUCEfWGCQzPe
5ZsVkUb+le/A9s4S7Yoq7cCBM1fMmr8DtciZFQbZdS5kNVAf9lyxnWvsuJPwY7xflxTer83gnz/i
rNpVB3OIbLIR4XZj7msY9p0m5bcyeMbH1Cq63LUPFqhw4kZugYwTWlyua1ObxKwZwl6S59ODRESh
HEK6pd3jIdLnhPBdGwRNY33dOSOsrIScgaklu++hZaWVkYdFlKn1QGPD4B0a6updPY8cI96c+SOS
t0KgBq71pd3n5aD+qx0D9kQjGcgk5leczuM3k915DceYFP4YxWIpxJwivKVcwqsmkoTMEtXa2pFh
7hLzTkE5VjYfuqMKTWblPhdA5GyuZ4HJ6lngIdVhrAiuL7bJKy+RQsC6eT4EM9KPNDoW38+xJIa/
bPDF+/gjm0trQKsjEsfEyWYnPpp7FEVgRWFywXmcA3zZVOLBYASO/yD4Sa3sF2ydoXLgvtkgBwr9
nWfFWarIXTO2qrIoutza0C4E7AkIEcC7ODV0YgipgYxiXwUIHsTXPaYMFcjzQARhvKrpkey6vtQa
twwgR0hTfa0IsFMYSLh9v6qZCh5KHkrfZDFHHdMeasxIhwhQAm0stUFPK7iqfuWurNvODIVNbfkw
lZ2S2q+mhDe85G1MW01X9y5Tv2Yh6rUJmB73SE8ER8nHvKn5Wz0NXjIEssfeEHQr4W54cI6JS92X
JczY47ICDMm/91MATDOOrfOPUuquZbO5gxhfmbW9gXPw0e7GKf8rjR16hfuxlXFP37KfSKwVAHtq
YcjuoyhbjkNT8+PPipQXgx1M86WP8I71qkB/pn5sPxHu1WedrIvcXJ/OMiyHou7hnTTEwfAW6m5F
UX3FHAnJI261jGLl01u8QViA3mIe5hdYttyVo/1xR1HPD+bxP9d/WRhkDrrTkgsiTtNkFqqV0Aat
nR9icwNLc4oe9yU+DhPMxgmr5fRQ3M896U1ODesYNbexE6ekogl1FthSDuJ2j4VSZUB4qSctM78u
XEMea7h2MAh+OwIYV5uDmScHY2eqB2smby1Wwa4PobQXCJRbmQVJRk/10LzVQUWFu7B8eRG2Qipv
42GS5HzVvvt2YVO3sEK+ab0GsRJ0VXCYzDO9Ow/hc3XHIQvjuPAMe5J7SrlFfmeLEKNsX57oFQ2p
/VH2Pe7JaafLdcB1BSmOoTNnMa+L5GSHiJv+gzlTJqOZKHFvFkJeDqIeb4CxF21sSb7s46XiyS5Z
xMUc+yU46JrqqPXRvFgVNQnwn3ozWHIKo73WSUCZuFt10BWjsYkZpJLuNg/4KWKxzjgNgXP/7yYN
WpZTiJZpMmnafTU/BfRnMxpWSoVjwlwF8QUftkUQjw7tBCcGMJmQP0uE9JcwLzqpJL2anSPL0Ff0
6aLREuQur+Xv1P5o6y25L+MLKSU6OklGwOJZHHfYG9Kzf9JLc0MRpgAX3zT9kbqKgkAMPvK2UToG
hEWP9fqG5+DlzKgZH2HfA2zteQNGsbx5gKJssB8jeAIIBSTVEFsLyGt9BLtxjxNMEGBXGjKPTNO5
smmf5+bW23JrFqZxjMC1IE8DMOezEJruEbtwWnhLVDWsNnFKQoIC/LDgsXOJwv5pfmH54h2vI4Ng
DmtbRBkKmbCKDkR7vJ74dxRLPu2KAuju4CtkyQnRLKiaRk2gflCpk232n4WepDrZemoQqQzr0iYT
nwCzgBxw2IMpmQFfG9BQ6a3r3VewVCzS3+9XmilRxVz5AHgu3On5sKiraKn6c32O4eWNE3gO0YIY
B9/MXrLdohfY35DxDjsz3dSsXu/JjjOivcWlRLf1hi2damIABzb1bGB1K21C73MMzLJu0EyYolyB
S2hOLvenXFNgqZc9KD01R/5iO1CIMNXVsjCT/gSarHTncvi1J9v7NRp29tyYaEA1ExjDGj9Mndm2
2/136wX4jPcOmU1T2Fk3V94LDQBvPCsAsZlxbI1HopKKzMfJYkKGL2xYUIVuXcM9ey3H+Y1746kE
X1SKtIdYbEj7Hj6E8bY0iwtT/V6BDhmQAVU4JUQ+z+FFQsMPJz4MI4m1c/Bg3b44T7BQG67mHNig
yHQS35p2Fzbk659+aZRqGMi54K+hJeEeymEsgY1FV/Z4PpeOjR5JJFcTKzWhy5NHzEzIIKr0T+ma
8gi+d2y8ce0EE+u2mr4hfH19d7zjMdqxwPcx+cdnDTw+NbsOzZviGwJOtlxYLseB3ikH/ejvxI5x
74GetuAiua1846p6hh5zPvY7RXRceSwllinh38v+sTh+SfZ7xjHuHT4wO/5PnTAs6Hg8Y0LSIPGv
pdzUVKJbiYXTBhp9m1CiN2G7Gz4VALTPFVYqMyZ/204/93GC9km2mfPfMFJ6RwSBQJBuRr37VeT+
nIPs41Ghm+3qAC7pcqpYmEoPuX2PYqe1cxDITBLpIlJhmMdgT8D7SjJ6RAP33HvmieFtYoGNItex
KHc7a7xDbDwtyhdM3mFD2Y65F5XEq5yw0dlq3xS/EYr3hwh9XcfeQy4D8lpEV73Pd/aiknS7TfxU
XIheZnOv2Oz/7LCSMPMzJ8IsePLzNc55rc1GwSjtiyVq4J9EUJet6g6UJ8gkIiarE7y4zRA+xwIg
KIgfz0WJ0aqjwzsp95lOs8stHn4NoFujvIu4m7MVYlXPhPwfLejXGplwI6eFAI+wx4EvoYDYFMZg
NEE3ohWf9k2OhmA2SBDc4RppmnGB4BavkSuLE2XKrsqY+DVgQ+rO8j3Ikn/wKQUfIuiKOSN07eSj
Dpje0Fx8ErWkRSm7n+0O0VIJEjI4x/DweAcgXmooTU3dacV4LibHBlg93zryC8t/+Hc8TgXwDwND
XZswdJ6tmtBulevs+zf4YQvdanWf636c7+Kbkx1FnyjWQkAwRvUofGdTqXAA+tU/7jsftCPgt85e
iHXtfimrn6pCU14n0U29rINdUt9526McR8EllHQG0UVZJ4yUX/ouKOmQ7VBg4N4sinVsieFflEm0
GhbNjEpZR5QUufRz2+g4ucHPZnfGYUEzeTLrhavBjWV6lGrzsFuMDajVch3+hn6qhJ8yVX+lnMSX
oi2YVg9Bt0u4TcVYEh+I+9RkkGi5WbyAw5Quda9YxKtNi8+xM/IvyJ+z9JJZ60r1yeGSjp8qsOrs
5YvFCcaj40Z5wwcUBvEY45bp0wRq/WgrEI8jcMnC21jR8+HLG1MxymWKAAg6PTySmSqck7pNqb0a
sE+to441k3MESXORLYvyxWcP1H0SDYoP371rUrmTgyuh8m2H9tFt6EyyGyRjNC1yO4hTc3+t/eiN
AtO7JPqreC9hcW4M1KelbfD0X6twVBmoa+JiknrqHGAN16zQX9WzDNdzXIs0ufnV3k02aCaoSJog
wlmutjnZeu/pj0BCN/JRARmtvbih5g14Y7fYt54XrU2FJiMB7J0v8tpmQRJVWvJEl/o8BrKAx1cA
9uOsbUdSMqRAvt3kIZDkq5zOhcXeKIL/AhXloDYUk8T/2Uz/f99De+EhR4Jj+ioHGfHLNlk4CHaL
l+O0k4NDu4MnW6mjN9Y6eSGVWNQpOqkJVZUdt9FuuCDUkOQ4kfZvIIm1TfqglpEvwqOqe/HB61RY
SKSqUKa2DXwaPPh1u23s8YLWzW4dlY9gXhhVUUDULDpxlAl+ZNrtZ6xadVoM70Y5mgp2Yj4Ce8rr
h0QvVmfTZRQTc36c6tsID8F5GwRxVQv/XwRjotkFtlyWLdVRnOGMGiqX6gk+vF2LvurqM89CWrcS
eP10LUh2N+oWAwFPVnMVewucDwztzVAeH+pivYk5jUXatrAPmGxF86rNxVIr91O8ym1tiQEEfnNG
ifhSIUnssgiNs3S89QVLibH2qyDUlXKZEjdIXVbuEvPz0ScITcj98aUey3BbjFt4GAldX78zp1Ts
LDSnvgIhBT7ybFAahEBUiOnMvYBDSSO642EiEQckotdpy4NifhWmPUAOdgDLOYQ39CW3DBo7euru
8lZqNS9RcvhuW/VmkyTBnctlTU6pPSk8comeCG/ll+xCqbI6wlDRMiXAGW9TmlV6HuygTwpeGD5H
XnjgP1DaKDtOiMVkz0P2Xd988MSgtVnY4PtTO+JLXhc4QHCewi1bD86IbOJxLPfTWY2zC6Pmyjoh
+NKTthJETcV4lvbXe/WCkKZlvYnU4DuvI9QpBrhiHZ2t5cr61ROb9UAS5uGEm8OWuu15gYrzPfme
SIvsIlwoRZqq5qfGPpisOfIJYeMwI3NuLTA5QIvr7a4AUYeKjeG5bL8XvurVMbt0zbxssCmFvwAj
UHc86ms04W3tx7aC5pDLJ2yfgEwR1+xxQwDW37jB2+zNtjBZRljQN4WWx8O4lcB8rLq5hJjPedKk
5DRyMJH/oXKSMTj9OdZfeGjLCIfFJc3k2IoA80ehLwWft9e/HismTA9dMqc9dacobsAyGSmUr122
c/Ze1zx6lTRqTsR3Mhw6M624rpgzdABRZbhQ358fzStYtiS6/bDRO5Wd9kjDbWgnvjlqpe4+4m3V
yY2tVHGMuCgdKJvtEe3NbNxTvboqDAkzeCUvrLgHMSjGNmVO19vQ2evDXCH2348BO9LLzIywks4E
znQ/LGGQrbFgLO0sKpxLYkbVdAvezgnwEGuH5hNd7OhMxjGxWhhZobrok4WOMqjssh6Ps7T09c/j
c3e/4pkSHiYlPqyFMfMNjggQRgxyEz80cSg5vwN3VF4sbTy3om4oHHbka87Nvq6vGcFq28+hD15m
w3AQspy0h6iu928zHb373OLF+/vJW76L4JeKaS+nsnQYAeRf0sCX92v5Ko8vF/TtvF8rwi2VmaZ4
rNftUvyyYo7kkyBnY0M69Hz7TOuNHmzvEpsbwdGrxaqpnqbHN4F/w+gEEQ/h12YsdmVtSM01sj7Q
PnsWDm89mEXz+LxWN8SLn1LiJeyCDGn0YKn4EKw1LkqWoNcE5t9rqDGITiEeIoE9+KDmThV4CAej
ZIeaVnkTiYznuvhqanTtH3rpzNCpntcIGeLabHsVUyja3B+PRfNSe3R+quzwTaDYGh3/o4pNACLl
OVA+taK/V/WU25OVtRzb61/pYsnq21O4lfu11aNL6N5xP4Lnt7JJlMJa2xSrfIQZY1exXidNSYKU
ZaVlc1Kb1MDyPI+mz5LepkPki4ccgPgsu6jIVTN2t0wJc5Mk2jFPvA1l8Nw94GW7eXuD2DeVo8FR
uO76KLtT5EcGTYfYHmQSnX/z+o9sCH/hnhal2ZRCQTwPmMZh8ZOjN0rAtXB3sRlbpCve2Sv36L97
UreO1zQbxU4IfZYXfV4WnSKfFGFJPQLNx/DU37XW+WG0Mw2pDoKtyacFrWjiHZ4THAfZkMwF3P+V
371xFB9lRlO4lCD/OtNnQJ9iNZ2iTwNTs2lV3sAW0Gxfkm1v9WKbC4sLe3VZbRLYdppTtDanav0w
6TLBuho1pKwyjqqTYtc16UReXFv0jDGoSb0HOo6rUOZ8YjEcKvOfx9uzqh4iIRHA2YbH6qLeoI22
PPtgE5mo/OSJjLHbQcIwbQpnv28xLzbgfsqpyFvY3kscrZEz52vu13ifVNzxk8OlavPRvBY+myRn
hTqtRgnJhB2keh0kkQSxFxOyQSvXhCWqdKihlaElOTWK6Szc5grdwxtL2E8pnfZWL8vUlljBazo+
QZjRe5Gf+3B/Kx7EubPojWgZmp2SsDbZnDXjWbe+mX2UEe62BE6p81AwvMuvYzANbW3LrTKyxold
Z5tZGi1kYa9Dj5oaA9LyO7yOuzeOHwkOhg4ynFzHyZkH35VW0GaUHJYcBgvi4oBPMGL1qXIZn639
glicnZdGP5JZ90LnDBotPpwWxNRlci7+CM5opRdb+X72jAjBtQaWSev920nAUS+aEB+4rgcrjlDF
bXARPSY0/DbWz4KDNN+jOhql90+BPJ9VvxRrxkZ6l6XosEP7h47VbZybvIe2irT740o+F/J9l905
H69byy2KpF0VOC+7SidSf8R0D5k8wzVzwQ0PPEB7TmceBo5uGNN0uhgGxg4L9G9c22Cv4tY8pjhH
Onv17bpWiAYvR8yVmCQ/BLML5lVJdco9l/wlgccYx1Yla6dosapIVe0EUJOT4w946S6JdxddN75Z
FqDDAzLyhl3fgKV69dqc7GCa2imMmxKzkcqRo749YNAOi7NndNdXRstbfoZKfTWD2Q/X1xRaXeI6
dhjnFOhp3sLBMgCZeEvBgXILzATmu149KAkJb0/ggDbzA1ckygtcctNUj9Tv7bgk7clwudmyUnrA
jBl6lPpHDPccvdgt8MaMp7WWRjsm9oVWGJIvFZ0hCpHTLCJnnHgwFIyI/ZBfhhdi3qlvavEmiygg
IHINTwZKS9isNoGi4IgU4X50kXjKPCE2zN4iBVlSyb2AfZrJOz7RbWPh7t7hUY6/w+uZe9DE34Vj
lI6kGlPUgdmoaj6YOwLSLBjhZYYRIW8Xb0U7Q7T7GCrpp4mYsfPObhrNEy/pWnOZS00pKockFMLI
zFnKnLEo26qGNlhiB/ZJshb24JPVWYwzIreciOli8LQSB0uxmupeVEFnWbspKtwE861DqwmG9VaE
V3HGqQ4ZhSey4cqri8qk2ZTMq+qepkQPiiWhXbnskIwjIiRaR8nK4dVfX5kfREqJvuJE1CBtx1uu
4H1z+Epy2GjiyKvaMMHMIwWO+193HqaeMDnu8pECpZ+dezY7HVeI5EOOXbJ4+bhHL3ZJ3KMU3R0I
99aoenL6/W4wvnW7hso3S+FEpCJTBRjZnr7cmVm9RPm8PqbAsKHQ3XNNb3yrxnWnb2+FvKWRFLsj
meK/2yL0hG6TGLlRX2xG+O2gyXpH7+2ov01S9fLkr+jE1XKkl3Urv79SnPc+yF61JY9e7nNakUh1
YB8aySRjKVteuQrjzCtroewkt5piRJkOw4DJvMqhZLwkhz/xh9jjxgHs6sZ4Mqa8kHrU6Sg2EAuY
c2CD6MZgHeYXwkW6XFzg+7Jrk9fgoJWyNRsnrxj6lZgiSjOhjcNchUqKHtAXTTOMJJLPvkxhgvqf
maoAVMcP3kYONUc7XzKFWkcAACLJee8uBhrXVrgniB51u/xOqQYATtRiGkewixuBgvhofl/t3i5c
MQYLeZY+MHnHDw6HckqtlehhsOr1YSHwnA/j6oelgQ7+ndZ64U8SiQ5lmWMrtzlxuGtetYBIJPAJ
EQxBYjuH5vUcLIMRi/LB49+cdCFD1csSMgTyVwTsZXP9XnCwOXzJrTb3GAiYz32HYkDLGBZxlP3E
77XsDvmRP2ig+l88NWZQU3q1rjyq4WhjDbX9K+suBTBAWb7SKqf86RW6UKKfdqW5wpznz8fP6a3W
DFGKaoOVJ3poTUdkT0vFinU5flQnZ3OqTXZDdj/laWxyPFoGcdwmnhmBMIA9O0L1P63spdl/Q7W1
GS8a0eKQQCR/Y9bDlvxD+U0toPlhRNiF5tEMab9pn0VwzRwymActg8vJYLigYqbliM/Oz9Rc3Pa6
2qqfDAOouJVZjZ2XGshOiFA6LzScIAO1VIHS45khjZQe1gaW7LAtA0jAhoU2IC56kqvK7/gr3c5N
WtsuYk9b0Gw8ZLmQIftLrFslSW+0d7sYFPdT35Wv4oWekPX2cFKICyLuCjRbim1IXdrm95WK+oOF
L1BUnAJ1AX8yJ8JUbQGKcwsJCUuLjqoJ0dqQiRcVYwBKgjuCj18HRsdNVpsTS1wk+j8QpBp2/RiN
PDM86EmKzMRqfg5tQNhh1QALDbwPGzK2S86JrK8rJ4JHXU8AOlpfgKcFn40RLzciRbeXuwvQSWlO
LguJQ+Ekk3wa/utpM732eVbtwv9iBoUGG90QO0rILPgxWplGvzYwtpK/omgmjHgAi+bYvBpUNQFn
5/ercaffrfFtJUb/VMfBKBwpKdBcLxP3ky9XjP8z8hZk7vEO95F+9oURxKbesKn52ZCDBINqYljY
F7MqO1AR8KAO6mbHLoCvwwBlervadVYR1ebWw9YwI71uBTA843llDqnsEKxrM7hF8TeGNnXKkAav
I6KVAixePgrXWb5jC+H2d7c+s/JVRUs8BloAJKcdRRI1W6onxXC8c/qC4Tu7jgHbtXUzf16Q7QWm
7ADvWx/qe/zfAIZgaB/UTFTEPTuYuuC1KTDW0Kl6gv17ruy3cyzDBbnVNHC2hUhiWggKdr9Z2jt5
YOTFAll85sk/wqz6oCU+K/rveEtHKMr/cB3/nEWlfT0BROMooZFVpiEBb1KG9xRhpReWh8RSY0YM
jMP9y7dNn9Hg+oG+n9yJuMF6y9gTrBM9cU8mP7h4ZVye8VwrRyX0yEXY5TOv7wfWLWmnsln69XiO
s8aXRzTKyoiUSmSr93CcxFyF6m2Y/8+gj/1BOfGhnOVEhaCt4IK+BxMywFDwwyrnYd3DVSbx+bAd
43EeYVZA4NlO5431QsglIT3hWmLQxCVyvKnVrWP8Rp/aPFZzV7fmP18XZSKsZP4DXd5Ix4CG1M7y
K/t7coz6ybHXYDV22fvj9CW7k7zf63DTmz8Ctb13x00vDJ8ssZJA0jezcE14YcyhdbaFmNv2Kze9
OdMP+RyjGk3rmKQoE+J4PcTn26HFTh8IFNZbyLryDy0Kfn0JUT8iqvYO3eqaYZRDLFQi7P5x/F8i
x2pA1xSDIIKy9ES12Zf2bkoF/whHqnvhVqVj4eOAy5+2+91x7BEnimJEwJ+jNmnOD+Wu1NuvYyTv
WesWoPmE+/FS/dRFPCyA6/3tem2d/tkDW5hJktuvlYLvVdJO5cwPy9VJz72lAyKw6x4ObC56mnIv
401gIllVVsLKgo2Dhr6ThKcYrQ35sfvAkzU+In3iFX9nom/NHJXaoZNS8MrIkNV53WwTJNWRbSSa
tOMaA+kG/V9fKP7lHldvm0KMCEYvpLmJWgAXTqPrtyyAfQaKDj9YKLD8YLOZMkzFRxTMrsutiMCE
1yLEqcG8GNfnHbtsfsF9KRFV+VpPV1iIdpL3Od1QchFTGrs/nVvt58eQmcunNID/RbbYDnULH40Y
Z4yK5mpUJGp1+ebLeoiPwOYv84pN0Cl10SI+P343/MXk+lRsqEkvgqNtGvu0CvF3Uqe9LKX4DuXG
EUEVxD6BQqSmuvwWRe0fB8/nR+wmG7RzO58+bBRAMolZvftKry9dBNw5035bm71/4IXJQjqa6UxW
zSTYUnJC4TPAUo/ksr0YcKLaw7wn64bNFH7HcMFMOyAwQh8w+2K0CHf6ZAK4J+gQbIZfuq2i4Wbq
kH9wlMTZ5E0Y7qh/EKrxdQP2xnAIaxHji8+bMsnweWfBdv5kD4E2GbtOQMdQmclaHs/IIJciV1+h
yyO8eyL7zXiYSI6DCVJgApK/RPX/T7BA+ufTzAQWDflh1uOuiU3CmEe1mtGRLIHIZmZmVPN7ML5D
0yZToOnC9r0FymZGESyyLZsPnxqNekQSAuG82qQSohwIbxXeI2vY1XyCrr84nGYjVKFjmLMhgRBX
NdYVKU8Y88E1kKBl18Od79iloQMJuE9nf1OSek+x+tDvuLC8j0amlut+RuWzz1hheM4TFWqfb58g
BIlpBRKw/CCQ3iJbsd3uMdP/hbvXvEj82vViVX4kVaSuc2Ta2vpwuJDyah3YVM9KLRKXsou8qI9k
fvcaU/R4VygcMhHdKG9twwETIA0pF3q/nFeq3z/2Usw2tjPXRPa5UTLfkUpiSERlYvpO4Hj/1dBH
aYBZaYLcbGPD/ITyHbVAOt6R+aPw1k4BW2XSzaPOTqEmYi/vYB+wyqgt80vUCxEezmh2LKxr+Et2
ULTE4n96zPLu8Ospy8o7VEEexnOzqREAFwPlCi0KIaoCL6jCpQ4p4RlKR9ZfCd11neuHoCqQVZGy
WgCAN3s0VS3Lf1BkYy8gnd6FZdpAD5glhJjl59AUHYSJNP+73uePyi26r2be+xZdo3zp6e10dkTG
DjTCxJN75ilhz6UyD311/E2kHYPC73OBID2NsiF9LQ06IQKikqRIOfVPcAB0W10XwTaiCptmt+u7
L6LONWzY+WYUmTt3mymJZF4BG0qi0jmpWS9PlHMqfqDq7lsao6a+5x1xcIoAmNZ0LZCuOKC3rayU
iVMORN9n4lSFTtyaHA2lCaCmW57Rdvd0be+1kSveSu7hLDxGOM3sj79SMcJItEvAMBFO2OZmzdDu
1OQi0aVfOHGkhnqzsObDk7mJbl7f305RYR5n5MFO1p6Fd2Yt+5IKryK4aWaa3Zw/L9bH1krQCtPF
+AzloTwfXUS6sCsOaF0wxYjJhjn+lCcrBrr8epBv2ttHHtw4+3b5eb4NwgLkagDOZxreGzxEABxg
r5c7TnKn/cO000xlDO2Qxan44wm3rqqkHGQUHRBrBXKCno1Ccmob1PsBgR144n6Rr7QW2Y6gFOzI
gW525ky+EVoFlMsrwb1WyespgyX5oEM9p1OkWy0FHSYNtsCYBgVc3mzL91Q2EqraDPzyTOP+2YRY
Twn7z8iMvSd6YQn4AlQIVYpvyj3c1W3O0MvRCjbiNQmWIGY3e5hlyXfJ8mWQ4PUSwpULgEuIHM08
OWOSOkX87BVuhbmAN9a4UB0xJbsahSGY+hoBPk7xjUZB+u2D1bbdzXTCSp/MjoxEfSHHa4LBgxpU
pG6WdEuvInjrhd+xrPRB1Cuyrk+dyHPBji/1nRlfS2U8a/Q3+6fHeN316nNvN+rLzYfkMPn7N0Ig
2AiM41D0QzWwfAOlh/3vUTQAnJr0YJtYsUo6v1aOAKM0RUYGoSYvakP09tu4NYRF3YCKB+5oYJf+
LPPxFOoThNJH1J+jou+maZgdHrlhnEaP5hURxvjGvueVVbe4+fLoBTuZgo4rIcxOhrFd6AF0PLxf
yFuWnCPJKmxzCWIgUlk+n6nk+ZTWVmQZv66GygdiBBZ/eCL3uCiVrPgF+pFJnzFGJM2pLQ9HUtuh
+7vQGwdSLeglc272k/TdlVMS3CQJd97ga90+f3IuwBjzDFsHZPeLC/vKu6fN7i4feRA1OV4Dqary
uCgNgQ32tu+EdAiyQaC0EXaCKUZCNtT4n9ZAmJk1IqYsMvlBnKrG8MIWmugZ4Y+XEJfN55IGsUm3
FgVU8lNWSQQ4T3hqDMu/OKCz613ZXnA4o3bgpvkOBEIdHbg7LH5iTTEdlomdRdogsFMHtzPR0RJP
unl+Oz2OpH/nuViCZ1PrAFG5mt0IANoQI+F6OIeO9uBrQfledYHkKxTHQc8T7KolgFlzSCfBIv81
k1+/5+mLTh1Mq5fRF/qqkLmJZVg1jtiMFB60qDegzO70UOCDXOB2jlGzwk685rfGUvSRruqDG672
GdJq3Wj4w4aUvXaYIGk+2htrnCAOmCD5bIPJmbVeDVLd+Xq9//tmwNqejU45Ix0/h9wUKUhQWA9+
2zJj/qzNszgNtvoitBOWVVoZyw8epgVkwrbi4vWNwaMOme2H9CaShOwbiXudYgSJpxV1NwSb7Oka
YeawVKjELL1iS5Tbcaq5nbOIR1Bg7GvpAr/NgXd2fXDPbB6sMZzPAYQ3K0lcm6ifWoIkOg0c200g
kSZcRoSzmGviWK/5Y0e2+6F7CRL73pkGBwDaV8uH3CutEefJGz+/mjB6ntVoOU2XvNEI6b1jcsCK
y7n+2CxsQyTwnDwJO3sc8tPQkVAuvM+P9hEP+Ofl4vVskbH5jTJsMCBEuesS+LP5685NmJ182kiZ
H+JccxUfPeQruocDRIDrjEA5cwEdwDrTfbwbp+gZIosuwgaEeC3Svk/4jZ35G6Un2z7wBW1OpT0N
b0Hh6Dled12Z84UHAcel4G5oLUoyupPr5Eg9bAmWssrC7kVPqH1E68AUMscGjncIUZNsSt26YS8V
KsgaNdP0AMVNyJaxdqVgfJ8UtH7h4MGelLlKRUjHzoYO10nIoYXlIKzdEC30n669gQRvxhnrCFnJ
XL0gxTEDTaBd/gU5ULAa0JHylVptK8DuibgI+v3AoNS/WnW2Qf7mgapdWac6eYdaHivfS3fBkmIc
AnHClgmM117Pw6p9DFJ4OgbU/Fhk5Tc6PadZfaZEg/N1iNb+QG3O1TyfZFBXK6kibM+jvA29uZcA
P6KuDnt3dcph3MVE0G+W6mVJUWWVwmLirzxrQ2MhhGcgxJBMcGYUO2aIxtbdUcM6KpesZUc+i67q
5OZbcPf8/t6WFUPPet/mnKB8ruAS9hY9gPk+nqlYNwoOkaZJxLYH5aKZH6u+on1FU2RQ0wB+Edm4
vBOsQe5pbV7qumxDKHto0Grd1NJgZj6qC5xuaqzEYAZoRp6guXaCBqV+1J3AokNazBcYrq9l+DEi
ki6TW4Kjrm/apuewJ9n10S7ZpXvRa3IThktxqw1ovUyRniVVWOjqeE9sil8JTLiRsg6eDojI96fP
+nJQbi9wlS12WOq0HYWqMRyci5eKTYT59HOBkVPeQ3IdwtTpR0LZ08mtFaD3S1/SbJVHLNQsUoAc
6fj3eBkfsCZvTF7pNcvQ4twAxgfGxtTreKKkX7pDksnUlRJhKi70SUrHImQSfAE9CU50RWgAzT2e
/Z14IUC//HcunFdZrRsNzAs6hrNFxvrnDoyx6JPJrP1UKwKOY4ofeXK51zVUBZ7QpegaAZVnmJ7C
kBYqx4V9D7ZcYacF1GsfIA49wD6TdfdpIFcCqwiVIkegB1yudQbEAwnQnKqJfcrgA0ozZL5nFRbG
XxjVN/phYoyq7b+vWqY1UUhpaSbfJh3305EasBWIxxQ4StKJV75BR9X66kx5pHku/BZnER/jmvW/
bw0hLBL+i1op2ZmMrCZiZ4m8JmbyzVKCkWa359EclhFzxlBKgB8ePx35qkphj/SfMb5llIzX0uYr
zpvEOx2dveFoUrEtBmpvXw8MvFf6mzUTHCx2UF61nEXBFQ0HFX9qN08UQWMNKeNEXBm61uIrkwzP
ZWir/Bf7TOOQ7DdshA2+Susv2iwV/Inrkx0Jb8y9XMuvnihDno96VNk2gFWqkZ9HHNkeRRQZN3zB
wgznHPVgSVWXkEN7grqNv3sgU26K5MjTmIZXU3TuYhdC55vy3tJDNPolvaPQXrHf8N5QvjjsgGtf
lb0Rx5tJMcZzxZAINQ/cSmHkP7P79kVmZ6QNs8z+4UfCv6xOG/9MczMhBbKbgu8pcbCt5V8G11LN
2X8a6Mr7FkfI2Pj+1LhHwoZc9hYG8KdhKu2+i2GkzLGCTgoageLFTXCDYRsI3fzDfCPLlpAAOMZn
svOKHSIyLr4VWXBiWqt9EmQDZaR67zqCXjJgTQqQ4HDXc775xGBqFFMIl2MtkVk3HjzZ+TFTup60
n/26MrM3YeJpJEtJSse8kvB6o6hLl1Kw/G7R+0hhhzMzxRas3Um6UDIKp2DMTqBRIaJ3VsUJCKUn
EQVtqZ9Rn+z5bs4UEGesf0llkN3sPeqA6oggD8CCqt/NzVfm2qryyoh4/oe8ksffmSPWFLwAhVHA
n5F7FUa61XHuXLYAdvs8nubb2GXhtW8pQqpx2S954CNO3OEAgiTVipVZxaO4eVqqBvRNCul52WAj
3aITqnxeHwWdTQSEr59YRPrOEIx+wCqAjRP3XxDVtclzbYQalL00OZBzV51jLcy35qRobQmXNMuF
apr6nnJd37zU2xsGsRXQv6WDq/QIDKdRgzE3YV+ml0/mp7m1d+I9r92ukgyUlaIeb5bnxCNYFGdJ
qwcffCFEIJ2hiv/fMneugBKFPggEe1HzOIH6TCSKw2JpiuPDvYYywl68v3wQi/q3Wxq92eRuda++
w3D13SblM/u71VHo+uIb/pkLPLLCs1E2yEWO8GNQs1TPK+FBWknb15n2xYsABVna8Ij5xtFakFQ0
uBAjQ18i/xkXFUGmlQbCtquVwUl1LYhxxL2rIOB45kd+KedoK1JCtUVowWHLBS/kLJkiFoEmItZ4
UyEyyxtihVGKEeiUV8Uzipc5JGeZUmmbeglM/EAaETPjoTAggQEAwqF0S6syYtcXlMS2GMLPYEr4
wvtJjMOoSKudU7+4/LL5ooxPOtwr/korudixaNpC0R8YoGA2qjYo0eKnvBy0biURAzso4fUZsEQf
dc9l1POv1VjlEJElaHI1VR6B6eaiU99e/zPYeQiDPEUbIM2EblJPQw0MmJI+T9wKelN+E38bQAtj
QJGSirTxCajCFSR2xZ170u1LXx6GsSQWU85UdYWTpAyjZBKsPyUEvulUoPLNmI0NDt1M47ar2Eb6
WDI75DggNUnJ5QI8g9smgiCEfZFmmeuJ5LC+52TW4Ztce3XZCEU+9VvLqcoN3NYrO50AdbxI5ryq
/ZtjpuDc4Eb7x8jnJTdgRGg7qZhhkfEOlz0L6x0IrCCt+SNGZheynFrmyGn69H5HVs+VMyXOd84l
VVUa3wQx3RBGc8ZD65QUsoMrswQXiTAvtnwrJlLexynber14Fby882AGBRjyLMw9WmBn4CA9xGRA
0/dMJbi0jfFqo1dgsIv8+vV7ZgbFtR5+PDvH9AusfKnaO3C6NUvYup8IeUqPj9eFwCF1QMb8Pp9S
nVM9yroEcsj7P7qxzUEo5SD5GuhoXcsmNzgWSrM2jjopEItJCIQxzbhMXsnASqYGPrGb5uP0eZGB
5zaJfPVxYl9aiYrfs8zgCOzAMwTkp7svCN29kPBjshAGKZeM9WUlH8JJK4Jv8Zb9Nvr5IGdZpPg4
9Ow3Jk+4oF/jtJQIQfYes7V1QT7FwkmO10kpag0ROBJ0VJbsaNjX7Q/C0jJZqL73xdDQ3rSIDPgK
PyDRTAo2yTbjkwXY697C+pc0zAogwDBC04N/WlAOqRespnQBr/ASG0R3qrWVrEsIizK0uajYWuuY
vdM8SHTTJGH72m7QuLCLpTLMxNzsHhB9QWr7FOcfVYyuC9C9D9CSU6y1pwWXE6+Nwy2ZBSNTnIEx
5HAuQpp3XckSYDpctBRvgjEJz/JYyfXN3Zp5g1CMOJ0vkd1lfAESzyakESD+bokQX8VIJWNxnVVj
nvFsayThbhZy0TLu5r5rEzZbILXsxGnCXp3NKbzd8yyRWbdVglgyWmM13bmgN+KXuIqogb3QtsXz
I0ZLDGN/vXNUr9WY5NCI+iaNbTbX3rWqHbp9CdWUH+fVVYioFI9mrTmfVHy0OWnqMQI/m5cXkCmc
jCfwNGkscrVjBfgJokEay0FAvnZIV88LTepvGG8Yxly3Yf33Gx9XF31ilOpThXhp4xoR60kJgD2+
nsctnseYWPNiz9zuRPMaioEwb+uJElUasMhbMc8AVO8z9ls/HLba79WFRkm7XUoO1LqvCsrxGL4F
AtN8ZseJw11sgNIJ2Nv5Qe6wUzbjp8HtZe8slXpNlOh+2Bt5h7FXSygB54OT+dBcCvsq/3WmYind
U05vag85Fz18JlWFtnMyczRfYLFSeJ43BUAfNaMbRZ1RpkaZmCahhsc7DpdZtvO7/UqUUbxIRjuO
c1pzG9hEi9fHOEnFY/xMTTWJUQu3l1XkkHZTYXdWHmEZOd5W7ipiResEWUAT8/ArSvtVBhW7DP4P
dcb2Cd00Zi5bOuOMGedfcZYCp7ZXb9ZR0cQPLMY1tCXhkCK8/+8pXeN/0KNHwF0BLJLRkJ00wmb3
pVJuIz2RvWWjRJycoSSsW2QBJKK5UqM0hreuVOt6rZt0KhhqPM03oCfzCx2efRcI4NUAOEyOpnlc
o/9XQBX0TeWDvCL+z5GlsEaiu39PvNtmXBMpTZ7BfLqTNYavnnqi8ZXnBwUQMcuiVHa0NDf+K4kB
9zaP43CBL9u9Dm1Li6jzT49w3y1M5u1/AIX139YXoZWuLDXVOEz61mz9yKhAVvBtl4Xd7jW0LrWo
5cqHbKBlqOmnvHI3wT4e5ttnSQYqwrT5wfCy8K5692ckoKA6cXvwqA53T+XGNdacOavEvXqe8UMS
70zd8zHZVBXxYYqKaMM4dI9nAK5mPyulmzBH2c+t3SzVRWak97uTrvccrW2/ltLKnnWeNJiCQ9l+
mSemOZZ1W8GZDmtbV7vA2QgD08caDa8CyMZohUa6Khvl+zKWL+nH9YlBnp95uD0YvrZFv9s/gIWy
HUidYChqTxlccrI1wgZpuSxqmfpeXE6kdHkPtm8WNk75evAI//bPvjtT97Cuk1rAywNHSAd9+EFM
WN13My8I/SDLgfu5U1xpRLT3mda6gtOqMVPJZNm6BuIzeBM2pQuwrxTYVPgW0dKLQHaEb57a4O5c
aApZVgdfka6fk+PQEVnscj3orikirzEIgw30Zj8FmhgjZfFSZzg8IMOAhV3GJkFrMPnltHMfD1dJ
iyXlR2Qn5SVHiTu40N3nAFDcff/cgjABCxaDLlgYSfHkfKcfmpgEpg3kJzN44FsBFDF+yG8gpMOz
litdcOXDnU9yqCnCR5SOYUMTeT33eARVp6rqRWmqZccnaDdG+QSgWyTrc8nVM3gua2eTWvau80D8
3AEOHkuaUw04k+GB8iZifFfW6NEk3yxhvjDo/qI/HU3HehKlOF6U/qRgaHWkF+7DqXcwkWEpX0c6
Is56DYCLJl75wBTuFgrenxwv2k7almZIO1/73yfSSz+tWJQvhoidXLl+33ZDFddSIi1baRW9K6HR
hWdrJR5d7wyaDMVxAo2vLjSQPGxgeouLat+iUVdOgJ9n9dT8SpJBnLcYXUXQVGs2wikf3M49cmYD
q+AlccCfgJw3Qgc+n9bwTqkYC1425TeyR3cvJEvPb2mwfV/LTRf4VsV0ERYCFGwpUYHPBtnMolva
fKcZY+Zm/Ypzehz3LFUHN4rlSPylwxQ+Uz/XG6grBIwDfohb2DO15vmHtrKUHW8lQJgIcEbYkrM7
QFKyJXDTXTug1ltNchRd40X/rClNNxF5q2a6SBg8XwcurvVYpzVcm0OwE9GAxn59waRkD/Vfib7y
qoIIfD+5RK9A8PNqKaUrA/QSybiO/kqrcXLqXc+Yg/lHUWK4JohywhzpFShNDGvlKMNeu3kFSwZ4
TwgUNR9ap2I49ND+rkSYkwJKrVzQVkAQ1AXFIocJ5uVJz+GSQoh1ero+1W3bo96E3uy0eWRq6Ur3
mmbhjJ8Bc3N64qG2q/41L439BHQjRxy5BDrgGw5hPrHZC1bmvH0pVu2XpwU7dn8no29tDGQz8xW9
nS6sFMPtHz8yGzQlhBkE6iURURiYI8knohQPPhcRvMpiX4xJg3wnZTirfa8SkEvfR3oWzSJ5Qk+A
aIHf2HYHZmGV9wJkGJN1+d7AWvEp65gQcBdD+4LI4QVTm+p44nmGNsAi0f21uQ/1M7/jV2e7UecY
ohkb2m+iSR+0GEwRjNQbG1nZGFLZdVs28WPmi6Q8S0EF+4WnGvCr6Rb/HVTV9Qvpw/9iskeq40Wr
aFHqGTkDLd76xkUyl5eFpsGJ06rOo/NB7nc5el3mAyC8fwYeVsTGvkwe3V8wQEouVu78dmk3/vHo
tc5Gs+u/u9dkDVikSA2a2s/C+msSZByBXwunTve0wgYtSV1rHX64UZxwJ7IfoqPTTK08RoOl3H5v
gKtNlhQ9QFppBQcagW7EKY2IjKAmUdV0D0/PoO13SxqzF81EpGuubjToh/YFsMBG9ecvUzxsvEve
YDcz3H+dbkhB3xo5AF0/Ln5T45QRPUBAkT1QXZk6eKxMDS/PAupYFKySqxXrR7vMBXEcPIoqkjDp
PS0/CdKO7XwzK7t1ke6qzEMJa6rCZOJ8Tw5TSfMqxuQXuRMU1sTMbIPe1iWbZZyiSNpuWO1mQLHQ
Ufmp+C3K2jBBxGHV1xO2R4RMBxq9yStfAMoN3aZhmDVDF0kvVS4snI2VkqNZj8TZExMQsA/EZUpg
URSjiG3nlFO4TV4XJilcFwbw97KegydVaXS/0DpJYxq489hffCR4NOY+rSGHKe5dh7tPRqOe8f/v
i2VELgcCXbBf+vqwmSTwU2HE+DZKcCJL0eZfhl9IvjidoXJ7plrfhNSyAjFRoEh212UsWBbjWv8B
VDaDoRXZAXS3xcwuGs4WmukF7nBIgCOWAPn/Lz7pF7aDrPtySbA53oHgYMDeM0ETYlx5/cuEMTsC
Swo5URCXsTOxw/VrKZkSHG+FU4R5zzdkesNDaZYKo8sz+qSa9wUCavpNbs0I4AdeUj+/un5lQIye
nB5G/eIcd1bYJZkhABFgPJ2joIIKfVfAmQpTYCCgbGliPJ12pZo1QW8OkPOuQ6YcpFgdXY6CL3qr
N90XA/GwSm/EBjtTPJD+vjYMayFNLvySmyyjmsaO/UXcA47b4Xp6ihgCKxsUwjaEh/+u/iVucAjq
rZyCQGlhpQ7WdUm9M4i3K0+aYpWF7Dg7P7xyaaKHg9KMQ6aXS1aWeRnF3NuyxcLnx9l2Qb4tzrPB
OpLIuMRRy4As7Uys2MsuZFVAfTxGIC44jOOToVFZWiLR32uw3hdGsA6tNzCNrqVT3ge8qf9FcZY5
xHngpnHvdicQtd0beseU+fMLrY47d1lRl32/Qwkb0HkVdI2/gIzXramjbffsciZ8vlYzrYNyfknl
ywiMf1MezLVeL+CL+Lcfp/JwR9xrWmJ6z1+xUO56df68NR4od/k4JrmadlTksK3xPKLZFkoUiE8l
cWj83ZLfF3/s9yoNKNSrBYdMYCPI5/1DQp2MtqFyT5GcrHG2rHeNTLfXSwK3LeAK7wIvt+sxl473
E43fxqCrQG+R6nhNebAVakCv7lV0VO3mDvtjgQFXwd0URsRIZa2indr8JpPbuiS+hOv63Hs9j+HF
8GkA6k2+L/FSsJedsKg/Z21X27SRRluwBWwYfhkyb6U6pwVEfc3+2byaJfo4gq6wCZajsmlTQgh7
pmlwdyQueEdM4Vm1vCbE8P/JLdjonG1+tQ+Ao9zUtoxg7DE1Txa2k4656PEY+fJp/N9T5gGtiSWO
zNxGU/eHy2Ldp85ckr+yviJizZoprhAs2I393+JLyI9xRBRjfrOfDvULjMbc3gE7yg3AB+6t4V5K
qZE7IZQvkL71YLF4o+t5EgHEsru+jUfMx/QMKkag1EYLxrczjCbgfXjMdrmZND/3sQFMCwA2n4fx
hHFntxIYrpH1UKoKgqg+bHCN6e0EPekmlaw5OYFxSNp2QE55d8ju3cSqa1eWdkKK5Nz1tRxlARBR
dljpcE7F+sWaISM0UlBGPzrts8D/xQ8ZFVVYcRSZt6pT5fxfdUFTcxfm81Jg9MFPpk3GhtuHldD8
Eg79ziaRY5HXRuIv0bKpboWfeDwwo9+PLjhs2iFc6NFUKDm5WNKqteZvefleOvnZXVwPKyqnMDZq
b+pCA9EE1LIduw0qt9bb8oeYREoj7RnERJ2KGTzIWM7/ArisZx5b1zVua503an8sWB/lEqQpLPwD
+XKWBlXjSlgkQ4yLfDtqbnxTWB86w6UvQTtwu8xqo/QbTw3MbD6yEf/8u2JqlRRP/Yw2GCazV+06
eyjPatR/boEtlS8ucMuww6tQuUoh+04iXVVoEneTTgwtWrsc84Zx61CZxLc823Xb9NjJwidEUNyT
ZXvqyAPsF/zx3KrZFdsy1xx22d+u+7Q85vv5BgBTcw/dqnbkThudHtBHhsJtpCbqNIfq5uNM/YJ5
2gwSz8k9p+lpLoNfDSfMhTlzjF9xIVsMMeKllicLIvyBh2m8S30ZTHgdb74hHIB5MZr3H+eW1zye
V9tgm7Xok4x5J2SHPziwQdYd3vIZ/PY4rmvsBkdzaW4pmcouQRRrfisVMq0rIIwMW21BDbFIZa+h
/SkzEEox/UJwbmOsQ4/6bT5h9L2U898YgHIJ2rnn4zxgTT0179SRnvWDtsGn7HAfj6MDazP6zlVz
utiJ4JVAyoJWI+UKAm5gWYFpOfrCvwOUjMTQ6NrnIoiE96X8CqQiY76RYZF5pSvtlj+L3/P7jihe
jGFo1lI7NQvdA0O/g6/ZT54llMkTa1RAMhkzEn/qtjLgJDrrKFqMs8hzZ0LG+e7G/gbxelSiscAK
WpEtCR4RQn1oUansXvLJEHDwbDWVkIaRK5OM9gv0e7UpE1IsIcqmuTrGN6XCeKUgXrcYhk13CuhI
VZJjbifdHLVVB58LU3sVqQ233hEZZoM3dBS3rMniS/87iCiKrs4tCcqfAzSMCE9zKaDRQ3jHJSPs
g5fTPFN52EGFuJKgiV9ovKKhBrAdwNe2nCfXP7njE6Q+qq+lAM520GgyiG1IbhwPJyhWOmLL3MnN
HWU9kbmqaSrfAIOqTgpuaevB7fBlh3WZp1OJW2JF2Ot80RrOr50fXtRmEsfzbDJGZ1Cem70MwNw6
F3S9qZCmTJbNrRizyPy3hLnWLHoVVMAmsR9KX+4WWbCpNWpPtHpod/OY3dcoOppAN79T2cahczuv
nyWe94cFsTh4QQB+KLhMLIaAE/k17iGimB2sK9uy3am1m76z/6JhRwYEntHffKFyltb/fiZ50fr4
+PjAyOub6TNILJebi4BcFk22PpKmO4njBP2Ot+bqVvKXKplZz7uu/GN3INDWypKNHAk4VvlCtjLe
R6giiNyl6HKjG6iwqW/iDcchWJX20ihr+tWRrCrr9XBApPxLqGO0nu7E6me8Sj8CsFJs5uozLm7q
Vo6V5hw9M7XJX2cdyYx740pSkUFrsgGmbxr6QMmf4tqCXpgzIdusAh37lXLi1vqTwfVP1ClObzU6
48plX74/It4ShuNY7I+ZoyybpRwNCPgzUABR4GxofC/L7vEKwWGSfNyeCnjTHGLRhEA3VV1wzZqp
wACqD8XnHjTGTJ9S+NkGU5GXzsRG2kH7Zo9gOxa0tklKz4idokecxn1PVwFIFJa1YzuF6b7Di12t
4cujidgsSEu+CpwI+SG/NIbKQSDS8eVyotUj/sICt6ls/o4pjm/jmcoXzeVuKPMirrYuoOFvPSPU
5VUNBcVvoNmK45rbdPWAXYDX7fF/05w9E8hRbb5sOWITPaPaZW7e3oeubgYwfAdq+PiTGa98wdk/
LXsgRnlxETIB5IJ8P/sd/Z4lrg5uk00k16UBCfVSbCfp9t4Gfywzv8jdixLL6NtDAyc3b0uCkj4A
149z/TzBLhxTd60b9ccvW/FjlAd2MPH5r7b8tQkEVcL1F9yiqs+Zcgwqaiwx5yhZN22wVpdTF4JC
Ugj3gg++C/AzCfu3BGwmPeVwPdA5JobM9MJmGB+qpRE/VhE47zFRWMUUlX0iAV9TV55nLJN0mjWs
AKFeEb3KWd3xsPh2NrUwVjLV8SZrRyC3yW7ymWYNGNy4w4LtQ1AyD2qYJJ52sqLp8x3GJZWseF5V
F98P/E76e97CngyieOQLQiE8dXwUVPbrJEPrR6vpmXa/0g06bc+4lv3h/zPgUGf7rd/hq7SId7/W
Khbzu3NIi/JARzwQtxrqHVCdIY83e2iCgNnlAUgob2cGgq0LdOafRDgys4TzYoJhDERYnWRz22+g
zY3RwkmWK34ezW9YvcbCaAQYrf0WpK3GOj6xz0OMvOKfc6UHMjxX7Td9FPsF/qi1jYZbWScCd9pF
HKC45qW5VE9cZ+5oYNSkoweFNUwH/vWa44KZYKm+uAVK6jB/6i+bsTa/JlulSzjjmeJKEtybvDSS
VlX3QxXU1sj3xzK+MbZKq40ZvGQJPaCud++RmLqcoQt4hklsjnburQk3TEZiINkwfS/dvGO26Oya
N/yIjdGvbNBzCPB8JiLgV4Fo+ZHxTPrACuOZxRX3DpooQT27/IwcwPOnMITLrE7EYCuL/8FJRvf3
rqrG/VpgCqubBb6DfOBUoEyegujUgsUdqGiP/AY/LOJQBJoQ0+QRMOMiPJSCIywmkEMVFeFY+aOO
p9MkljvKZiPkhynTizMrBHEbtyyP3q1AZPVyXdJTwxX4eh9NbHbO7WFo9BkUubIDxJRL7WOLOrhv
KAGZ8DBrQDCvReEtOuQimFbbvIKArd8osRnFlQ84tOUQ2wCQp/QOUyVFqqk2/dU2jwV27shSwdNC
lcKpVo74kdInpKEfjqUM8WZ5SRUX0d0XBY1YWdIN4OacQFOf915lFk5vSn9+YRWjhXZi5flvk9/+
Nf6eFNcKTJ3TzF+65MkEpspa1Gr0Jit7b5pBSh+L38JeKoIxQUyN8XD71Ndh4Y2zTNwLcgHtv/nU
I7TaeHMO1WFjPLb63l2oju71YxAVd9RTHV5vEQhgQvsvE4CAM6Rwv51RAt2hkUDfKnCw/9d7KBRW
B4gpmQjOq/xAi4lnt6yXETVoduBCTk8PvXvxV8ffipw78oCJVxukTHNQD4lrGvV83QMpsA93S0Ht
CULjmHwzABZ6A+TMrhFcnSmpbuRRwj0PJhznGDMqAeILeBX+uC+vIVAo3Sh+8Vbphyz6ZdbEZxcI
OkGmEeY5EXxLM3qk9muP7oEwvclVklTCAduOu7bOFf66NqlgvDaKk3+DhMIMiDZqSmamT6oPXswj
1T0KakdaIY2nUe4jUm8WqFkQI31LeShLh3a1CsfaHAmjwKLw9LsHEbHfgAqQq4vMbdXneBXgMxnC
56RHfxSNfpIrubktD2wcIVtq0bB3cNCipREtobx8lr3dtCsDUM3k7oqr23DMcoEQTCQrcMaZ1Dxk
kxyLbk/CjeYvQX6lQbKJ7bvvBJhRtJECC3cPrJ4sncncRDalsgEBZRyO8YWW2JefY1LYlti4gq1o
4r8OPvq2aILJ88kp7udwDXViMbC6z1zspVc/zc0m8KJl4A8wyPn9FMk2I7fiXND88oS6ITnmOo3X
aRUyYV/3I1Jaa5SdhzE8xSQuetoPbmxpvEltADZaYXeJ+fbO8KiWL3XRZHNpumKwKXD10+49L/gW
XOwQALmZi8GbUJCyWZTxq8lct8oldx98Hz0dvxheOqtwTerfUyd1QgOHinhd3wiSEioftucBUxp2
RLCWiI9/ZTOcNyeVtKKs+9kQcsDKQBbkeNFTZplbCxVYG8EPyuoh4PfIWM/ImaiJdqn0Zv0K4MOg
3on/KIw8/PWH8w3hvmgGeFCDo8a3d0rW4npy1nRZR4zN6FJadQ8JeGT3PBfy2B9IYPTN8n2ggQmU
nbBXHSYpBrqsZQcH73cmGHq3NaVHaUWmq5SHD2hyGdXGNZkf3uoNC0rHA6eZlP0MK0HscXSt8LLP
wk1UAkZZP4IsBD6lsSNNrFGYnMjtSb9SYxYpY3jswE3tIgVJz1CK3XN9OS8CTMdfp6odZVVKqG5Y
k2rlAPTuQIwM8wq+fSh/+jA3R9kLkJSHbXY49XPXTMQkvlA/g8G94aptY17s9DCIzHx8ZykSntOp
48ZZKsaCjG35mZCg/fFd5hVeMvbgaS1Mu8RbeJle7nJgc2pgsAPLOtzkxa7fDQcGs2NGf2BkaXBo
znIkNy0Gnha/WAD73uomedo/t7eVig6gLuwoLuhw3KjtVbnnvIJIhibyt6Bd3PdyaBQbY5lGYdIY
iLJO3o5lMsYh5Xa8yvYZ3Ht0G1F+IiHMyNXc1kApKpdYh/aSOxsSN1qWKOJWjZXTRtb2kyncddYG
YhLl0SaRLkKhwULt4Swe6H9H+AyWA9kVHuoPkhxiHBP0SwqaTVYGMBzOi/NdJuwh0sgWaDTT+xJu
vuTiLzwe5wLGPTaU4AVpjCwfiDrpDzJaMKs+rGsb5D+Wak0otEEZfS7rEuAjhkmP6lyibaMGOUt3
GYXvMSXzC7Hv3Jpn4iH1rdhoNiLX6bkyvyO0ipfZ09p74BNHzvCh0ETGlY8FAnoj6vA/wKhyFwFc
shnhGDGHXz55wx2wtKl07tkbZtWFtk+lCGDnbX2WtG/lyrB2xRIe+Z5WKmL0PUs/c81GyUf/ThTW
zIxowvW2aLUxn1kB7JtW0KQ63/NUVXnuQUwCHsSItEe6c5fUPoksAhOQBxiN7IGHx8292j2s8Crz
cMwSUvCwYzjlUgbiOcqsikaa5dn1pC0W7Epj+fErqxLD/roEqpaUp7JKp8pA7Kwiw/0HRvjqxErX
HsGROPsnNRk4QRMYUZ6cdwnYo/KYIdpnmP6R29kzwk000w+wBN69xHi8lCzqS0XyCjpIXqLW2boy
Fv1q3ygKWbQP7Vbl26JtOIg24mlLm0PSF7GaL0oaREuJ2dTI5wSIhIGrjr7t24j3CRsxlsnXqSja
b2I5hDHf28ni4UgGeaietFijXe2DsJE9l/Cf4tvx5LU9taQx1HG0YMRawqWoI/Cl1L3crrrSIl0V
ONfkrvAon8UMyHxjJ7tpeLz61YvfFqDc+xFbJ2/pUqQVwJJtDBwcN5dDyaC2WZLZC4K27yMPwHQL
BS8XG+2C5tK7lCHzzkP6wm1ClOdYDUemhHWmOf70ivjcNlFA4aLO3Tk65duGUSBhdccPS7QXeWHL
L0d/BfznAAxF3Y2NAf3wyT3+wL9SI3upEF7QUikemqzTXqHGInJWvxiGePGnvjU2kMCrl3QpNbT4
kjek028ZVD9ONKXCyENV5HL6n/FFkyyxgPnpaEwTQONFPwH37pQZOy/iENuLK6zZ5nk77H56Ev4T
QulenEcvtc9RAGlE8FKkKy+oP4OvCnIm08JOPMQ2xyfr2Y8We0kxaaq71V6QFssNdathTAHhe4aw
tsPsXQ7MUY9HZiI/q+fopksmdQpXMQB+ATXyRQBwbJsLF2RAakErZ6vyZpBSZx6q5BCjq/80BYQR
g7iFf4dn0MU9fiK53Y8icPXJR5vcaOG5+PI9oDj5x32mmHcpw76RhKOAWUhjr3z67kzfXbcwbc6w
6owFeSPiJJssZuwuxWrdJymHE0dgs2OmEz+iaf/DEs8KnSXeLS/acPXl4I4XDxIVym5dy+reHamw
l/nTTEvGEBJl1rFu/jJZCqpki0qJkaKe3gPoQEEwyi0q2iL1JUYoc9A1+O14FD4fa+39wSabdOQ9
tnTtR7Aa8l7eoDz538COegpg8xorCyxkPNe3ujyMbxn4RbvVXU3yVfncPzg1sizsQ/ahjdmDy49z
9w9SW22IqKHi41hSmKnFbFOyAVsemF+TSFYPIpaO9ARFPH+Uh2F9mbz/6kWf7/HjdvhW7+GR5RHh
wiECkHivSr545tX6rFV25tsqVAeVrTXmHmRxli7jkJtWUeaQ3ttZzz8nvII8vIQ0fmqPFYn7Z0k5
fEqg8ulPTsABKuu0RGn8gjIrjplT3E9OphgMHKYUzCSQ0TG8A3qcr8x1RwLbY1E9N/mjexYPvCdc
UV7ZQGe0omMJGo19hT/OA9acWO0HDupnbGZJTV/oVn22A9f3vltywwDHBot0YiwHBi/fukiDKeYd
JWeTYSFz7Iy4sj9Cr5NXjTfRhXkJX5s+b3bfGhqBU4GKN1fCHlq1j1FZjAHbSYqa1qilgdu3OhwM
XYqFfPEsko+YVlXXccpeIAETfONEDyGmn0HiC+2KnlrRul9F5XPXFmOetBD8/0zllVTiJ/7wbPg/
iNeFgpNoffyGC0GNs+VrglmPR9XIMdJmWXBaFv/iaBtsh4KDrIBfxxo4s7ey4gqp0GGT12WkH7BC
VkrsTSDJG8EWhL0PQmlr7AkNaQCN89mzYg95zL7WS48YFwhP5NIXSBoR8vZ7T8WKLgXjLE+dOYKO
GaGckEUE8ruGqw1WasfoD4bUG4G6HzRoLnZ/2XWhTAvrp0Mg0FGYZMheLTn0xN0Lrn2ZaQEVT+LN
JwiDH+JdzNPVFGWabszs84uaFUdw97aKDJFL2elk9KVBbQ96FZ0D05ffqcVVt9XX/yACrMrSq/mH
FJs5gdcNAah9n3gixnYM99RHo5vpcUGqi4hWYqkfR+Pn5x/ScQDzMPYQX71aLtojQBL2Mre0VCxs
4DG6yjs1HFQfNGJEX2j5/OhZRa03kaZOoPLexzPGHqosSZ1m+xmEzm6GuNEvElyJeak3ydjmqHeS
n0df2EBrrz1FzJzTfuYp4kyIfVDuZdwO7fvbk/WINNyMOXUybQMexm1i+78k/rky73iLmJxvN49o
EsWspaJmu6lqPSf24HyQKqj593RUFRTIiRuK46LsqT0ImowQPxWQiWLiSkZCSC9WBaeJzim+Gqqt
Pf9gG2GznsFcHM3Wsipwk1R6E6o8FlRkqvsdmrW2FtFEhVCzflfJEyrgBRkRouH2mRq1axEnvc3D
DUOGZA4DJeV5ffm/5VRzZGArTWXAIorNkqsypYVGl3PZTqFaOXdeoem5fQe9hOUgpLsDYBDC+rmS
n58odDI1Sey6UsP67tEDrLJyADzPKfrgs92uML+i2xdVO7mRvrGcu693YDkVnT78IgpFAavYtnIO
yOzg/M79VU5BHSK5DHTc3ZP58T2EYGG1RBEVZkh9WfG3QjzYI43cizmRFGuRWeNFeoPw2yzP+cEE
JDcT/s5NjEYADhsFDSJE2n+tsbLsHhIUe1e9iIWJGwEtR1cW8lKa5LT+1anQA96a014YSsep0Za+
b5Rq9NPtIxkfS17LgnALSrzYhsHuBmMjW/WjkveXjap+ZDRS3xV9UkZManSBMBwqYld9w+lA3CBv
pogH62/Pds64HBNSc75p/sGSngYdiheNP2Nn6TOrN1OBQczmrP37AenIpMBhCZEeBDLOb0Uex2kL
3e7oCibGkQ/u/1dgODkUbolQhcypkNUtnJq8LjPYTAv3RjGyuUETPr5UFGZ+RZIaTBByjDqfUWdk
Ae/eSA0chZWx8gJXRvgGb0sWiFWYrN+mOqm7LCYTnbFtEq18jNw8UHQRlpyzbYJrGg5DuLFr08VK
Oonz8hf3bxwMxYx2enC0GTmQI7HaGxl4kENw24AZastkK7if4J7az92NCN07LpsnTfHBZbtSRQmk
FLj+D8uFgSV4xeBFXqhKpFclzAyulcUq5KKfjBKwPWKX17M1hnl5qIcCh3iio83SXpu8PrqmDwqL
pmGK2ZAX/aMIO/0//+9Oq1YfVXR72kmQ6V3Vcz4IWyGKB8OoxWn+S/rVrVbHQ37HIGmlx4aQzGo4
KcCbwtnzvMdCs5CAap7XFrhSJGW1RwW5EUjGcKiQYgNcdwYu6U96WQFVajyaw+wab2WqBkbPlBvM
XidR5GB7DaKUK1z018+KPgvkcClz719ApJ9uwrD+ivhdbaZilMqoe+cAlGFaM8e/8DW0H08Ylbfq
F2iRjmw5WkPIwbdxfPMR7zwzv3dVaUu0+NWZKGI8+XlRI8gULnDRiqPizzWmmMfVQIg4dYZtspW6
h4tbX4RtEraxqfwn2Efx0fwtZkmsrDPR3iJMqA6LccFkiM53J2ZJmKBuwacc4y6mt64Ybcwzrpfj
jxZHOLhpwIprPmGGHoUNdcXK0xUadEARdfFfL1b4q/4wIgSNL7Qpvgz0BHZWSt1yQr+BzPOlqjnL
cZqRJdlVeChWtdvyfyKeRxeb6hFLK+L0h4hx6MJhRByQfdaDc9tU9OrnbqKBqpB+0zXwUCSRtJjY
J++B4AlQl15Q1sIsv0Cx0SuWmKBsx1YmCLlk9wfrvFfKTHOQbmtjDJvHTI0uPwfSgI/CT2SH42jv
rfIPgo7iq9TK1/qgcFskCv/PhWpDmib7Jj/oHUecBwzTHV+h8JA6UheW11O6Ntjz0nt8TMMgzIeh
SI9F+NypGODQqwIbazP9O8sIyxRiCchbw4ftBz/8Ppdlwgj7mwvcNYWFkQEf6/7bHu9pkwV3dpsL
dew46cupjwQoyZ95Ns2w9mKRUjWmYwhnh+a26kSafqK5uGumG7e3s4uNAo3h9WaKhmMB02jAoEvB
OxzHUySmqm3BqzeMg30zknfLVVVaEpQCI7hVyf+bkM83LnqGsJ1ZNhmKMNzH+YDyWnug1sxTxKDy
nmp1QsA8fng2Dzve2JhfuhMk4Bix6UM31ea2LC477LTdBdmxnwzikHom9+GEGTATiiGEOXOO1/7b
emsoxmNpiRSKko623JPK9wqheFZq8sFEzXI9Mi+wwgRhv+piUyFZk5ZlD8FfTDB1ocVfqgSOKT75
+0MLc+TwuZpPpx4w5PzyUpgc3pTP4nLpmvArAqMG82pXO0qR/dJKFM+dHYHEb8DkXhUs5a3VBt50
RBfWou5WeURfpc5SGkaD4cryaGwB9PQUIut6WbRze6UVz7duE6O2YYXk7sgdYlevSMxDqnE7KT0T
F0mRBv4VjKEIxgrSYwUUBTjK73w2I/Ti9iBJyMuLcKqDlk+oR69xOIZLi5tUu/hsfp4NRJ5RS3mx
GkqDpoGGHYRtZX1RalaH1e2/CILnNd2ejz1dOwIlXfd6S65mfe395AXol2X9kePLIcDn6X5Vy0Jc
jXhjmE8X+GrvXHvUzvuq7440cWbSUZ2MyyluUWjDHkwyeHteRgTrL3EskgzXJGGcq8WdtMlIR9Bc
0CMuzfha4zgaOe6KB2Lr5Y9wRI9CXWy3sNjAMjLDBYaPMCorMCBApRkdWn9VftsxVXo98m+umVYv
LVirBV1GKB+iuBum5/0hmKQomA50jShuZPeXf77BtwfCNzNsWTLya9RaPR7hhA0HgNX2ENeYD+hx
X8UGhxbUFKskMgs2ueN4loGsDbLJDnfJr75BwF9KlUBDCdeEaROEsPe8ApMGiLBRpEy+bZJOuT0Q
oljBeX3nxHkoQLrMx1UwhCONFR6+y8vvI2VIBWyRLdggCVADBO/oVtCzINH/oAPd+Ab+zVM6F0/E
zLL3GaTNN5JTElqm7pgyAZuZBn5Uy1PO77i7kfemhBzGyk8ohJkNOcGYYKRcuiShCAgLfVAEVLcW
rnR3iryaQdBEIJ4iO/f+lQ1YLcYazlfnYVs1g/psTZs0C3/wzRGsAnAJ2hdsSqe5L6QiMCuEy8FI
Fx7GNKnAi47Y6LiWEQEyPYwaQYJRK456u0iIV3jYct1RlJfN/jqiLUZDvXoctXfTkrzEp3mR+Crx
AKLYxYCplSnrDFgKFcDC6PqmrDIOghD6JyZdWUxnflmtLWluGKBT6hnG3PBjpBYku1U6mW418YFg
RGYVC6jpXyM+BDSDc/aPT0sPdU1pTmqoclZTLImuDL1WE2LsgldDFCWm76W/LQs0ADpP3iJDi5vY
kRoIoo1FgGNs8UpHm8RKkT6um01kSV0lNwp+qcyCZmiEC/VsT8d8QNnSYT9Aip8QWYYx0QcdAWeT
gxrDX9lk4AsBilm/6kzxWx4afo9D4+ii/sEYybkItjopoUxUeyGT7T5/ThIifK0/MGg02qogTJIr
xhdDEFnG+/cPG9nnnHDo4TPy37kgsMBL39v8XPJAz2kjl5QLeypIoIp3q7zvx1UiT9ucoLTF4LrD
MUnoFu+Sl28rZ1CuPrWf+f3G4ibDbUDk0Fz8fhkmtfNl/6ZCF1km6CaP7NBokaWkQCyuYjMHOMIo
XYbTI/c/t7q+bmOZeBrYZv/A8VwI+Ibg5rh8t8VGZuaNeBsYBip0gSE7XgsfBaAGyd6T+WzSlzIO
Ehe+uKtRh916hkU1STPyFdm6I6lPMUFpV6wuV1HliKOCvfwlTwUbXwG9GrYwo2BcRnU2vfCGK6mE
lTNkKeg8lh0mlBFBth3s5FqC4SwZIqXMXeR2X0ADUoB9+h5pBSG5RFXuUgjNS/ulNse65iCAc0en
SOSLZEiR3nAaOvYHoAI6WKRUTHsA5BlZIwE+HsHwU7jA3mkdfyx1K0p5lG8sglw1UbEc0DKznpHg
H7dKuWBx5obsFngAu19xAxBr8tb/yJnouJY8lvoYzUPC3S6/LaSAT9nJD5ko06PjX2HyG0HWwVk6
YbmHR2VDbTEmHu+jWAFGHwaNtg/zVyhruPXkjwWVtXUDE4WJ9zMxksqxC5AodcGV+PQs/EKDHWf1
ykVA0C52Ke+HL4SbVYwZr1ptRcd2OMa+Rx/MZnex3bsLYdcLQExmmT4WyYdhtBafydOimn/Qod/t
XwzXGaTX4j45YUIKhM6Rrw2qIuUVpCON+uQCvzHZV9kR2epe2JqykDNeYyX1fH1E8YPKMRHYZLS7
iMMINzt+OIq/ahRAHMOOR/e06riy+IRDbFM5cLDU1zCng0YMofQmZNnjOzsFLnMj5shFjhilMaU0
oT/VC7m1M2S7d6ZbVZKEXMBm8w87V8UicaLrC3feOXjv6xNG8dfmuDPUQ3bVRWrT3MMSbu5e1t/x
b+HuEM+vIBEoU70jRLvtLEFGnrmlZzWaiFTVh2+igDHQX1mN3GmdtniGLr2XUTVN6go+ukjy7U8y
CEYPGWKb+7ZoHh2kCLkY9a8sRGCAX6TPWH/dALWMvjMZyxEaAUKQ6+9yF1l2jpNi/swWaCrc3zAf
3co4C2qCIhDaym+AQgvcLPj/kfOvAEpgdqbpGDnhTC9KrxjbIdMc2PikqJcMIR0FMnojz5XPT1+6
eA4m1BU/23UtZYRQj35VfZbrgnIDYUS6+mqjRYftNpEilbw/W4xtJurEuT47LbHSM0XVGICmev6B
TUgwyRfjOZb6e6Y0hTKHBe30+tKOclv6YP5nwUNH0piWfwsmnz3QVMg8bit0HLjxJ6xVjhjXcZF0
fEyPNQ1K9IH4fuRzZ5yK4X8Dyz5cOfbGagiD73WPhuwM42NLvLyyOC5tsmZWxvMcNEFS9fdmSPT/
eNTJ4c/9mhUiK5+oH8UXUMP2jCf/1BdQkaxbYWzCK7y5ac8Ack0eM0nxmKm4NXfrQOLxGUotXB/T
ZZrENXYBQbJT9O3PlI4OQVcWzileVE8VJSNaN0tnrmHPbUkEvoQNCPjkDXIbsb02KRXu1fuUpcNi
obDVVQYrEnh38oJK+oDWC2YpbPpnLshBkqo/lX/jpQP3b37tobPGlrOHYg26C8Y+NRwIxJaMYEdW
9TnBpdTe0AzrFsCLgwUUvCf0i1kpQg2Hoh1Mm2qS6V3p40UVc83Au8/7Qeu5LQKtARkv3wXTWRuk
a6BBOLv8PN2lneBaMrYXiRo9Vp2YHm2biBta1oJ71wvZEU9PnVuo19nh1OzKqtORyZpZ19nsdune
5+6RuaRTxyF4nT9H3tmR/PV7sFqKSZCXnFQpfSIdKMqO8R9M7fZi0GZJUWacu4b/fH0qI71I75zx
U3yGd8stWKow42uWQldg14uZ7hVIsde5r3CnQPJA1608J1J8MT1EQ667C/12JlpIozaua9BfBaww
kjRj181pjOZJcTNpTf42dH6ezxilsmgiUNeHOl9ZnHsucL15FyBQL0NBO1MBt5Tc3nLX8hNLLLzy
fCZ25/qKCE35KWzsSnKSl/jsyT7DmPxMNoIJcVIbnC5niulSG7iqB1UcdyFs7j9LSUC+YpPmkyKk
0glkGGYu7cpafBQC41i+panTIQUcupLMhWdbVyTm1Kotu4n9TDlFI8IwvtxldWGHHBxN65aB2CYM
+HPZUeHrF7b/o5XOOiRlO/9SvCnOGlWixvHH9o/nd4wTIlWpdYCIq51kBtkMOTRMSvgYb9L9Q5iG
AYYN1c46TnS2N3BXpeKlxCt7w3vHLkHXyuoSlsBnYcG5NU16WKLq9Ig0/TjSOMEQ50Jmbw9QmA01
BRNXs6QjpFMvsv/Df9WT486ymo7jJBEDvxg+OMcx+woe6VHCtwTRaV824nmc/d9SKvyfwxUBw1/C
9Rk6UqtfgUL99rmYtg/PtIgHmPgGa3YrkKBeCe4vi8dK7/S3sX716ZT8QboEB2xHlAy/NN+oiXoh
cKJDyEzqFtFZiUug3wi9xXJECu8Kjhbe33flR9jf1mWy5f+ziqiFmCQECtH9wRWtPHqKqoJ1v0Jl
LFeYquFTurSBlJMzAVREhkrJBbAy0R/OsRxA1KxDPzkMsTDvceDhegj5AdZKwmGfy9+j6d1k00W6
49URbVZaZqOhp03dP2PAORBOUDZw7Rvgv06cdb8ZL/BHhmINyCVM/puZfGcqMLXixNtR+WzYZR+s
0igEWJNgAS6/mplFtHJ5dzOiFLX/YOOY+o0z8U8tJPJD5+Gy3A4lYtQrHVFRIiJ7/05iTS6SfoSY
xrqvaUWSTY54/V41QPVgFyr82V3S+U/sEIdxOcvNz7U30h110AL7Yx9ygh2axSfPzTLo53SnPr1w
yDH/h5u/6kqUWQBOCIRIyn/1s31j0clx26bn5IKwArVEanTrAD7dbSo5TQaCy05foPUNKYsPms+I
6zoATASIzMA6Ab7uUltnWx27lni4tSSZ865EfYQAeya/BsBNImqCzwopS0ZUWDCbsYGUuysjj+72
If7bo8/v1CexgxCNiWRT5tQEY22L9GK2Iz/EjmasLDQJs2MVEpdFqA+l4zXGXNtqYMjDR3brGz3/
Py44f8IWS/sB9iglASSCvfmXk+ZNwSfN8b2B8tyD/ajmXeFjpVyIknjVE+nMTUdYv1aQ5WS8sL5V
KcxrmvKvXqTqJGzc6zGtXyo/7sVB6+4iwrrYuqzOJpK58pUow6dW3P4am9uxZkCjx0vjYWEnz5nV
I1gU2PwdMKBwRCWlg8vaQmMPFUuGpHq8rodvIe/f37DdNcagVtHOTWStJHDyqjOuJGZLuLv3a8ja
21HnQ15wu95M7oqj7f2uEo2W4wA8nQMt1bz/HRKvG0NWvmmM/bhKUPuVYvEKDViYgJc/712ncFfh
8u8h/5asbXMj+LIo91hfmty2pspaq6kUDYC77f3W8MmGKJ82RvRB31RH4XjquBQi8hrzoulgVUuo
mbtiIJq+SKS1cVuYofnWCg3sRVh7D+nSs4PyuRaunRQl+l55OFWljOjDDURHBiab/qL8BdoQl79o
14mpusC2hpQXK8c7A5iJ9ReaOpRdgRCHzEbytgAhPRrtEfPDoZly6xVIw1A4BU70hxLc8EYz/hC5
V5qIH3rGHTdQHzr9v0SsUjF75kuNAxCsofPAdv/8RatQcctkidH8lQJdpFeuWx4L+9UqbANskN+G
3Uy5RHsY9+ncYWl8PygMNNDfhVIVynI68ImqzauVN8NXIVH8VT95y5dJdsmTufK55K81d+u3PPSS
AMOKnA0YeU9bo3XmXU9XWE9rw1hsfX9+Ybx5Dwae7OLwHrzraumQCvcWz9LomwXDxCtbj4L4wLgK
/kYPdHBvxUc4njfooleaU/cwFb40YfIErYPbMT8pWrPgc1nLWoshVM153rc9ICsBMF7slRAfCgZ5
RDbcsgDHdMh7VMDYP6x+iscYJvNf/85RFRaD2bPiBP9EvM1Axk/UVyDR5Y8TPklKTS1pYBfhwAf9
Y/UAwQ1Utzv48lYGXuBD1LnmPKYAkwzrhMvCJK+uKE791EpTLcpBK8LbiXbgdSyRL8MIqPWFkOPt
tA5ci5r6zge5L+vBo4n287N7mAZYa4j0/IDFAElNVvLKl5n57bDhqmR0KadyM6iSJDZXJ3reaBMq
rSaMtlRhNwySclvFlz6EhpdiMOrGw3q+ceU5h0Ur0S2ogtMMv8ZDP2tBHpJ5djww7JtsGA9tpJEp
ad9C1OJ9GjJwv7FWX0NIrjKVjcdwZKZLO0Hf50CHF/JS7iny/eDu4aLApmqSv4oI1GQKrezOoB6o
HqDU6at7HtROqRsEcA7SkXNi93aKV2HK10cWdQ8++up5y77RxBMGqk/eea+tsMePdBNh5kA0GWfP
nzgL7uVzWtEDANbkOTUEzBZpbGWcxf8eS6b9yMMEYvJ+jDxtxYmS/tVL54rcvOoX9RjaSB95xY0R
RuGBQBKzoxgT2kPZOkBLDZlBvS25zhOLw0aV42IvlpBU+BXTqxhDDC1jwJIazQ3VQ41aluK/28+q
9vav8QasFBb2JiE3B6D+Rlc/zbOdFuIYpARlkl/B5lOCRuyFg6VetB3DdfBffCggd2yaARbb/KKY
UAzpD1PohfQyZDTQR5C0RJt4Ya757j9Yl2op5VwQprVDmcGJrJCYviFp2dOI9i/PFd6syJ4mJ8Xe
AxEv/XPur03HTLX5sZJQwVKM86EnBKwdDIXvIW3gUzHH/S3BP76aYJtACsryvUjC6h5POxQOKwuj
FYBxPxSOat+e8Q0upmqoj1y7ZkgHqHjcaeYJAd7p0YDAdZyzUBnCBzBuEgUVppRy1aQU2i+G3J/7
erba/aHxoJidU3AanPIQC9eajKy3pygfXBeU5fQ8xntzgCsqLczlwzc2v4gD0x2WWRJzkeJolnPs
+FpXvH3EgDnA1CGxxBsI6kMV82WjXbC/z3v3duMj8hM5/aG+fAY46iFUFAC4aPR/V8p/jMSTFKIn
hrY2+kLyUpiO3I3bYeTP2sH3YknRqCvD2jXuxkrg07L1oDk4Ps//0pXkMZujzjZyZ5vZpcZDIP3Z
QawabRrAoSPk3wQX/Xtb+ZPRzgxVF95RnX0kp/OhJL4Zfu+4jQkcM+AKHoqccu5WfoNSNGdV/MU+
CalSP49aOMh5MdEUVM/Tm1Akl5AHmOkvjtTbZRKW2O+7HDpmJ5HON66ZjJrYfZ7oM6Ki6Rxwe8Vh
shWbjdutDKe8ljSd1A4KalGoWqtMOScbVIDMu4793lrmqVTO7cybOTc+/7wyd4tIxI/hdILNX2kK
sFbzJHXLB5xgYnGtGg/6g+6QuQ9LPvvJAichXD76RUAVY2cSOdFMzVD4YOFp/wKC6v04ki57Hirf
rwrMtDeJuha+iAraXVLc+HqzxHoEi5t/5lZK92kQ2TpBfDWCCPg6hnH/IrU0GOPibs6jKovzJb0z
jrTG6dU5K264cu+M6FEEIhJs//69nc+Cnuzr0GFydOrMffL/KHH5U2re/YpIIYzAtabtHHQvxLmL
mDSpEExRu6qWom/FDA9AZJPeBwjqETVJI7Zwn6Dbr4sV7XonYJDtcVWK9F+uXQWsExZBhyLBRI/O
WUz1cssvFt4FHw4HyiBG5vJWqzoqEML8F40eqiAltFEWvbB5ByiJrl2f5jiXgnTxYS/SJFGAYVsl
tdnNl0RTXfkaCTJrpBTs8WmhldmYILiiOzmSU+6MNPaytIdjKKPlgqksYR6sFuXcBccRm9yFobUA
0eh4iDGjC9C03Qeck9hKOmAYeJQVPlAh9qUrRw8PcRu1UJtjG+x1u+QQsfw3nF3xyAnMCDTE2tG5
NWtbgGVC8/FaPcoe9eTY+Wlvchxh0uz6vPlpFZ+UxA7rwNC7gZeZVIRShpPaIJP0VEwfP5JOqqT2
DyxNmIAIJXFw6Vd0+s3cKs+Q6QIXo4pO1RCZS9bMt+y/5Czc8oiD8VtmjNHWLikW0zEC9WHmomZA
SuBuC7aAFu0Gku/bOsbHkgttW3N1T2iE6UIlaHYe3HWl9gfzyuAG4V/cpx6XM0Xxy9TTGcqjhpka
FYgrlKnub+56tiBiOkibNKgYkO4w818gswnUUqtPpJ8gAjrYvT7INMeoCtUht5C5Bh9OAcjeGfit
yI2eC99LuloQV30S/zGD7DqVmuGOPwk6NGqp32AzzRsXhb7318fSL6bkEF902ZDyz+GE0kzlrtzZ
VEMhBdD/3QqanzeGsoeuYwIeClVjDnth++jXaZCM9/VLjaZaFaNinxRU/rJkY5JM801e6X2bizRY
ARmASs9isFMX1Q6ijMbVCGAPMEuWuAy3DT9K/XOXO2FrqY4Pi1sJ5bf9d5rBRd9DAw3jGGsrfXJx
PD6CJ06VSykuibiF2/MGpyKiTPt65ISSyVAW4fBq0mvn/RpYMExIpWLfvTX/C/XQ/mjIzL5Wjw4e
4m8qCGsjLi/5UUo40MRUlN+02BoPas2WIMFhHhhoCk319adwQv1DvGM3UwkyGpHQ1xHxJ40v7MC9
t13laOhAwqHLsO/BpYvRYHqH97IJYYYt75Zp9o1ufVwaICoQmdynfP52+XB5qoP0JMa2QS9g82vG
8xb0Akq+EWwuUt6yFxIrYviiJU4EoIYIf8tB1lrn9OWJtzdMBAdLDSm1bnB0KBlpwgEt500RFLpd
0IkgUjeC9MSddw4+NRa+DRY56MThamLkktHvYjfhhc5/nyqRfZk7nuI+BAUBGMF3Cz3GVvTDqj2P
smjlEIkkYBCQGA0h3RcO4bv9iBr87NkpoQAQPO6XBn9NP0MJhcb5wBPtAwvelgSOSRAbFOu8YN1I
RQf1/fzWyEHyOup6YYof/2DHK1ik1Pa7jwpcUHpsoSIJNbVw3hcMSTJn3U1jg3/OhNtrH/KuSrgh
q6KOFy4RvshjJCCCFZf/iISbSJkoSXQB06cbReNpDDglCvdtXpMJfc5USnsfZT/bP94yewSNgeXc
IOU0pj6BpW8i5ogegN5DzrKh/bTF+esEBILV7RhBwxvUmYjY2jFuvPmBXSGm6E7wrsYFR4UQftv5
e+rVE1MdGUCXF2G/JlVBkl4pcPpVj0v19uZ0TktMN8vSy2v3+O4fEwjzRg4/rv4ovmA4NzaVtmdR
nTX/IAR+idiwb1CkQmy2VKctGPgDWUgI761EopLwThgv3nPxxirFN1sk8PCalrEuvAyAUO3WHa6E
66mo5pqOIEk1+vf7loe0klRYjCcW8KahcAWS7y8EjVxcbuje3BQcC7X9x4iHANImS4nGc7ca/r7z
/Xri6pBQzPBmALBe3tbNcACR02pw5wcYsWPpAzYJ5/WkIk4xqzyUKCEzrquTaubuLRxn5qm+9W+s
/+LmZWhNwy2knqoicilFXtKjdstxkpp9C8b6WuZyL+CRp2/2HPYk3S2BLP1cm6nPcV3Dwtcv88uP
L8KJvNJooRlplYzoOrp6c4A9JJwXq1CwmSxwX1WZ8dy+xBdV8kfEAh3O+yPdR458OdyBJrCUUKQi
iMLancv89ckjlIaAkqv/FENpmdBt7Bsae1c6ii30lNd0KRC81Fve0aw7KKIw/T4XE3RQQKelXa/N
U3oK3Ssaj0K+1f/jKD8AdGqYWwMt5qy3QE6aN06Gm5ApxZkHSrTF96khcxeXg06V1d687j9K+TPB
kKMG2oZx3dDVARJRs/Nz+NxE1onNaYm4dOeAYcFb1CmioHXq4Zq/fgDJXf665b+P9BFaimLKCYx7
WDM8bvAuHEUMUvsJOvYgsj50vCbt519VV1EHDpb6hCuR9M8qLrUGXrTbcAa0i9X4RnPHBgzzv4CS
3LEh1pzSKAnueNkmnQ1bO7wpkmQ3i3Zv3m/qGiPjFnGMmHHFNXyPjSsWhsOSdMHy5/mv2ORF1z2I
UqKBkBuR6xOvreHviGpiDYltX/OnRNTN+mcd2Ce6Ci8fjojJVeP6d5L/Z2KBi0nrtj9+LGsi3JsD
xahx5lsyf/VZK7TZrgz6AsfTHHDDuWc2teQdfRYmmdEB+xo9hfRr5gpdATABQRjkiehFDvW4KECx
bXEapYTF+4rNr+CLnUbY9vfEhp0wLtSC12lVOgH3xSMSsEpeqSe3Lvpus51nqDGWJmaE3i4Uy5vC
quYkLFrfVSSny61Wdu9OK4EoZg/oeP7TJ5BEFosgki8vALnhABJoTdoZU1DF+403jUwvhC/9/NbI
verL6RuHk9ilF1CqPq02RH18S0Dc1Gnho7KiRdUuMhuZUhpjrl7NO1cUAF/4UqMVFvFA44Agwkty
u/TnGBV9HYDsznyNnpohMwNGyPK7ROw+RjqgtVY6V1CrChzz3lrwfUbZMQsCuT2MvwZmlMxo+R/t
vzyth7kurqQY+YKxH1IpIW+SWjvlk87gtjzGQMcH6F/Z1N6MwPiPhNhviVUBqgOV/OTvCX2V3Qzo
y1Nqaj6ckKrkDQM3A/qGCUdKSmgIcsy4MsIzcfheRXPl6iFSD0o7c7GcaPUqvuUnieQS8G3KcanZ
IgkkifbAsv020Gm7OoQRCAriLezPEDGbWeLiu13qCWyIjJi5fqDq6hKTGwiwIkD7upJYJJvGfG7G
c/ehBrmpbics9ekQg1M+KYayMFAqD2iYn4Pt04gToQBa+XRqw4Xkcqrs6Lp24jhuRVPuiIUBM6N+
HAnXRWB2v/PxpgpZ+OrY2ZG2jCXQM8iDNm0/vGFI+DJP0USAnys/uPWEtW/stJuHgmFu9ykmcBl8
y2NUHB77ygn+kQGnKRHxGPWlYTxFVAxXlgHwsy3UX9J20Lv73mYX1eNJmPVnNZ43J/tAhqSJZ9e6
5e1/SYpQDCMZDz3T8D9kUHIjg/2i25smYgULrdQwSCfEYFq6cuYqpdB2z/DuKVwSk71wny21VPCd
jwv3ugrt6yl7GKzybNI8jCtApNtEzgVvqyrv71a43Z11px6029c4iv7GlrPVfzQ39UzK9jWP8YJ5
L/DoDM04rfQTqY7fw1tBOg90LtXHa4Ae2t7+kZTUXwzqVZNfU6PrXdADWD611hPg7FBeCWoLG2Oz
hGeznurVDLFPgl48sl5de/+kP2j4c29cmK8isw9TX3r5cO2FH0DxhjCsPE5CkjDlBWh6K3RAatkZ
U0RO0T1vmuKGKOCwobeD5sPTHbv8CEMhjIIEmnItB5ofvkHvVoCdBNZniVdgJisC5TRJh8zZZJjG
pHfhQJaTHO4fZpS1y+yjCyfdbojLJwELuaMsvAuHQhmkFBYX9qeslisKeiJjCI7jWINXD0vcCUlY
Xd5dIyh1AnJOEVQnZ7RHyMV/e4Q1dYwj2k28XbpJMDFiD3LuK7WZEdT6zlGS7gFybEkdFVAHVQ4X
/l4LjR9VX7hQcs5/Kux9CP7iEu7jeEiamLe1Lb/Wd7IbqoXDr34KLlMmfkPA5Ej4cNkcNLG0SLca
29sHW4oo72ZlGe6r5+n0afSQIHsTUK3fWoBWGiUb460vKgZcDl19+VRTA2l2MXdxOLrEqFhLcVLt
4Pti8/LXng+pzvt0/fq7dSqtNv5xA2CBLKk07B927muj/XYccojdiRdQnQMw+QmHhEYJIyd0gGZY
J78L5DOdPFNOLOqD0naIjRO7Hs3QVVfLLrWhaz5frykAFTosPeb0KS9mimgv/i/Dm700aC/KZUid
6s9ZjBsJF3Rmxn/RWu2RV5rrjgtKoiINuKFLF0A2AS5khtstu99YBj5MgMhdpymga+pEsKtQ4kgM
tY+IdZNwLrh7hltGCzDXhOu2p8Y98eHl3o0yUdDsquISnBgjRk2EQ+6U0GjhsuEQ6ilpIQ1jmGsw
jCvsWBqv7X9FKZuTM4l16uLZ+MlbdYx1rNT9VNqOns7rhydBG5mcm9jq7Zxu6lJBGm/QzovmuWuV
J8isyxmI+gMNqt1UUPxUw3MWZw3hnQY/4TAqpkf62LJtQcJN0308gRkTZSg+wKxGWGd+QoyVdkeT
kuBFTnjUDnkvD2wEnhXUo/1o+PjVmjne9lgjnIsKEMj6YzMw9rZfLJjcDmLqR8FOLuhOsilX7heI
AkD1HnYjQ2Hqy/SCU5GgKcG7UKUplRd5KZ2eUm96PMgtCSnScYMu+EmhK8+OuYZ2XQWoQ8lEOSI5
8lB1MOJtpimt4C6G6nUW4rXz/LX+LnTOleMezOz2plI7A2DruIVY17L1BvHG9UEUjbvpAgZxAcz3
0wCmdta7mUU74w/uq4svop8yj3Wh4aP8hue1H880E+5FuUexrXhBszjNQgUmCM0yYa17CoQlDN5T
ivRuXYAUrHyM7SoGhwuBOQtFu/cw8zbCSd5iAk2NvhdOQfsmeSvcs6ijuXYc+oK+mo0UTYxmIZQe
67Hdx9ZzMaMV33BFXsJolOJe/yefRJTow46dJaXCzFimdevNYixp2aBBGoaZD7TmGVYuzFJGvnRK
N/ALVryPpF8E+DmEAiBQm7Nqyfvb95ZqMp8hZlzho9O3ztJk3H15z6rJtAz022ILa78tvxPBVzk9
/tmNbZF62kbZc7jTIL0IsUCPAf1g+8Hszu9bJSklabwTCkXCmDCTqKe3ItBG/NurigzJ4LYxlgV/
NRNzBFUjkj9R+O93+GcmNn/xo88fJ2UNe6su8kjMjQZd5upSwRxTW4eVqtvNNG8qx1vu4dgslfTG
FVFa+qStr8If9Nep49oEhQAwm7LNZvss2EYwnYEb4S39mYj7ozrwnSFZlGkmXw+AxurkxjMLJCCv
vyN3Wiyq6PBJXAlGfHzHTIkx1awsjJQ4FElmY+NNiMFVF2hRIEsdN9LtHBHb76w58oQHybKtUviO
4yldCWuzoLxwPqZKtLCwH8BqlVRyiLeNz5kkgXE9rbvlIg0PKQiJVcydc92ht/OUMXUu677/p11t
x6+rLfM+N5TToHi4JO3hdgIHIAgisF5LNTXGOlpVJNqqvYx/mZLLWlUtR47FHOMOzbpzDiNP0k9c
fONoMzpwzE8U+cf4BdAJ6XUKwBw7W37rnMLpNYfSFYhrPDQuRkKXVQ0FzxR4iYeHI4U52bsf/6H3
w4aBBvqbi4+E1EH80VXw8Qdb6pbXpKk/RzViogj8ABZT996WH50ag7t2CXd3fZubecJKqkVQLSxO
DDiBQGH7rz0+hoUAycko5jUrv+omGwqo2bCeIu/lZ1R2ARAbp4/A9wg5OsdDS6j3b96ZWookjWiz
tzAyldxzrMavQuHAEsLzTGnHYe2IKzxOMvuX0meOKkynEDOBVvttNEpCgy9Od/MeyciY4DFq1ZLv
WzL119RLxVP74qEjrKVVzELgWOqQ6SnJ0xm++V+2mVpEenlIvgniSffNdv9wH16pBFRWIkh1QfG2
FFcVchFWUtjNh/LOjbTJZBGYexDDA+LgJODk+ty2ynfSwsQV6HUBfHMZRCqWLY7Q6Swxjm/vWgdp
WUUd2NdxOmklpWYSWGx5SeIuTpUnREZq089b83osFqqJCrlJgRWpnxTBCIy+M2Iie8s8qyoniSqb
7nS5FiPVLgphK1ewBSTMpsuZv7WXwgxQeJ8rews9okkwcFbaybpubttA8dfwPa8h/cqfXivKEuYM
iLN8OAPjXK23oTAmUQEaVwJDtf1B8tsW/mBKJNbL8C01L7ggaUGlkIyS5kwzUnnUH7JKI/fzrXdp
nIlNGjpdYMOgmOVLCj2pEe1JBkQHA4n5y9GMvfYPTnPgEL0JXHbWF4zLASkSLPty1/zSmWSKJHoz
S9voKVsYS25SlXZjdj3PDSdw5IVt+sZ3IDPuvL0Z9hDFi5nhTrmzn+vDC0dLoTzOmPYNaAQwN27s
4/TV76JrrWVUj2FnJqo5IEK845Af9poNMUSk5QTL7r2qCglyornQ97CoxjxRhtFEY576DCUDRofq
gQ6ZuLVrln3uiazpvtErcv22IkeY4br/q9dBDgRqPL47WT75uEISvGD0mFUGH2qXT7sRcN+dgZwG
cy6MOaKgV0vgioo17L2ARl6rDRepiE8iz4Y85oltzErd5KtHSbhwg5/KNka+CZh9zJbIrm23UxZa
ZWJs5KS6Gxl1U7w2RxWbEX8a2jcecLHAZmhg8TvX5e8CwQKxHC6HXfx5JJHg1c3zvZ3G5ezAwYTd
U8O9MO6L1HI6wdBN8ZocsFGjyjlM43bLvU5vuxWXHHiJ9I3oMS6Kd5mInw0RwklA4eHJ/z9w3GSq
VNOERGh9pIbrq6S3E0IkLFakvgSuVYJjPRoMCzGjlzguRLcoCp+pGT30/ooGT/j2UVz1Qk/rolua
HmAe9ZzeOyctN0V2sKKRQZhRWJ0nfEzTZWHjFb4R9STw0kpoU8OmojR3khp/6rSnC+NzBTplvcux
cNLxIlHkfM1OUmdRKjpP3qa4okTQN6Mp8iZK+iIz+pxqN2PkdRJ2/Qc3GeDLFiXFfagGItTaOC1K
ZVkCv9iTEORCfqAAS3XuFdu4u6IUsVsJtIRSQVkhXlyL6N2EHIuj2cBvQHCrJIJTuwUxfPKXRBOp
gRtyoN4hdCraHZAMMz3fFjS6SyeNcqNuJRm2yjhZNR9wysEEWFvSdwhqD6IiJoeWkro40FjdOdBt
TPxsCZnIx3vja4WZWBm/c/EIXpFZ3INnEX7kvFiuOz9MZSY0zRqD+k6uwA+OcV6h40pwvtPnk79Q
IY+7bHDfWUdJrXlm0tvH9LSiM4K3TzJg/4YmkNgK8zwIrhM/0fOkSk//wLh3fkyyXiphuy0mwhTY
L6UfJUQb+aV6f2mkvXyEbwbTNyRxC9X+1pF6TrAMNT5WZDu3gDMcIGpPXsu3B6i8pCYB1bHdyDY7
EeCEo6yoLj8Yfp/tcZosFUlR76vYUtIK70q9gSzCvTmAi5eZt63eQ4FN59rTTAFYqVq0Odg3Q3ht
Cfcx/XkIVQFX8Z7WoI3HVn0lm4xpqtadZtsR0wZvk0WeO5iTZEI+A6a4/f4Oo0uTSzCT7zR8Ux2L
kf8Y+juqvVE1AUaVnN30YgLSRxT5kwhpQI/REc39IjlpYxbWRXYd/UBaZ5GSH3gIxCgOonrVMQMi
KlAE6Qh3Iu0AosjYrE0e7J/pF10p5981zCl61OqaHurlYQdXXRpD89nzGpIdnsLfpNvae0MtcKe3
maZbPC6AvXDuaQ6h4SRYpujjUyav39Et1ggxX8YMsE6uTN2o5K/wycZbv7p53U+/AQtXE0H9CBMg
b7c0xAnXV43Fz4ptKuyXPRJl6JahmJEQ7Y0LvZLl1f5m/b7lbEwJ7iyLAZabeUwyIC825J4som52
F8TYbEw44qpT7zDmj88F0aA55SfVv3zipylYxVLwifEf8e+CIql1qoAfCg3lvPnugO0TKX0ErFH3
jtY+Epd0AlM0RQYLSbqN28JT4RJnVjI30ocaWn74z7Cg7emm+hy+r974NI74VjdyAGuXGXpbjfM6
cqrDdr6ihrWfVBCfSwNNl4RaS67vVFG0Ahv/NgbLpm5igERpjndaLRkyqROhbr2hG5AeujT3/RNO
rQ1rXTipa2WE7mBNlnQPKFxWJX4BYQQWkmd90gCRMJbOEW3kimnMabKCkEHDgAJOuBNDzCK59UmF
5UB9vxXywUvY9PfjtVPQYb5VNhWn+Lc3yBhjQgIsHFFtdsVDkIXKkD28Ywe0dxdxTEy9muSURlfC
gGkafrn0LZ3IrG/nHA2InCKaV/o6zu0+6biiC2o4jXZWqkx58VAyCM6JMW48xSI0y+pJRr3htZg1
YaemXOTOjga81WyB4F3E4XQ3uz/XfB75FsKV/D5TXRByRSjXJLhkX1Qqdv1Naf6eLxky7NOmimXt
i9C82/3AXE/zM/qzu4tSILTlcHY6qbly7G2kfdIZvPUtPD/47ooTg/1EFpsTBvq0SCAfH/FGU69/
OaRhmr1IZVWFpLPnKC7XdqrqfP4WdLsJ3LI97ZcTw4ozT+Gfo1yyS5Q7Z5omAq1CCySHXXgy5xD+
rQPyMBSp+H3Ue+wdxcoKqCQpjm9yaOc9OGK6Ohp4rVnzHMRHAwFh96+dWyL5yT0t0ct+KwNT5gVI
un5nAG1/guNyVV13SVlEIUjBuJBT3ZPnuK1tPH0pxjOtOi3hkHPJiEiKEjBr9kw1c4yfh7IDiBGM
Qnhv3YObdxvoUBwIIJjDvfJJdL4MxoZ7IU4hxfTpYU1xVyZ7XnbYnqwEGOHdr+tcL333KhKRhu3F
80b7Fo+DUNZQvTUTYraO2zt/S+aOZPf9fhbR/v7gqR03ja+s5GNaAuMkA6cRFs9mOuFtNdBTI1L5
dahquV+T/OmkFLCSM2G5DIKG0K3vqHhqz4YVF3hmWT1Sopi5R9M+e/mNgv8DXO0QI7TG2k0xWBnN
wlZU6b+Hfo2bZByKl50fDKaTQDrfcbdejWc4Da4AEY+Vdq12oJpBKBImmUpvBcXvz1HlnVk1J4/8
SLvbhknoI6bB6MsxLZilDqtGPSgQJiOqi2BqjdMoS/KN3g7ArZvJx0kr5YcJ5bwRMsf3P5KCm/Mq
ejoZ6H7Ty/Q2kjmzPnbNpNqjgLDiUhAZvcvtvDor7VfxpaFtpSpj798pU9MdpjQFD6e5FV7F/YOr
RG7aeOzX+6XW9kxaS1vA9JqLREDGY+YrU8PtJkne2JPhnEU7RKrYakUJK4USmi21ZRPGXH0tgUd+
s9xuzc23Tx6sql5ZrzmGpmH0xd2nZkW59cuNj5gqRi5bIcyBwntvIY/Rf6+f9H64IJ3zVeRBvk6N
+ddVlSmBAZYOgSlSXvUUhDFLFXg4FFgx4/yZkP0m5pV5SvrRPjIG3N9afeaXe9RESjtyT5vYMEAA
F2Ses/qI++hgVQ0k8HJjNOqzh10VHJXmYfz0OsfA9NYy7zlRDjULeu1D0OllXzPi4ENmCtmkSrRd
HiMUDnz1GN+tjr80/twVZ8StnBon1tRjdZsD27EGF5Mqtkyf9XV6hVRBsiFdZJHstusJkUphzwuM
4qDssk4puHy40MSexes4icXqjuHNyttTTFex+WQnpFpryCZtwkU55CPM6i6x8tZzvDPXzP+8+Pa9
Su/TWn+kWRbNAROw8svS1n4hiHK3zBgmmFHhTckZgZ0TSxdwi9c3BYTqhiudBGbdwH31wZKYWIrR
/tLg4LmBOBpyL7RDLJ/0RjD4CSTIkFbe+nVJ8JOmPra+cJ5tl/JbhaD57lskRjOit6iL7oAarHd3
pRc6hSLg43du+UngXEMoYqilhUE3JKWIZxBI/B/yKu16lzWa0oczM2qiXNPY/DUaDsCnIOI7k5si
ZsKYy4+sVhyKsIsI6Nh6ZxgNTfSmbams5kh2E7C/EUwel4GomOQdRRyfq/wOUCFRSdLzyvYeQvIJ
9IksGF8EuUCee/vh0LctrbDsz+h22J6ZtKAy2+XCQ2MouZd6rDy+PwZsOnk7deVxUETdGqe8V2lt
sq+b9QiOFTGq5nPsY+UPjEnOfEjL8d2dzYVU6RNhCxY6xseo5oOUsxASPlsD+pMAcFqYgeEYVIJh
pYMA5Kku3wE+SAYqr2oIHqqS+D/e+z+ZR98UlGnklPC4L+i4Lhps/Y8BWc3iU1TNDcoph9zlfOGz
Ll7T8PgQ5faOFMyCMbO65dw/dpvqg0XmT0Gy675j5iLKaLGDQOLgXefhEG2XoHQDMDNRRbd61UvU
GVwPcFF38BozbJUOR0lvV05LJbdI8ZLRUzK4+hHerMkdeBcizgXM1NV2hLlQODdYMTJX8idYIxCH
CJpvIN2zXRTI2B4zqAjP0bOXg+IiSuV4sHtl3wGomkZlcGAi+aYvn0vsLVwSAgjm+zkFX4+y+q8+
7gpAkh3RFjH39j7i/3y+TparDOoLJ8P6fcCh48u3gmUEnsw9qIZm5nxyAyFkKOMHJ+dbfeu9Phs3
l7U4lkEkzilpoqPCGgAQ1K4+oXyQrxYhJxqJDQpjXZK/XsRT8B2fIhWb1GMxIbjNI3ibLuMjTkzY
bxZMqDcjVPD/vGE2OCywaeJEX5SFmnJ4HXr2+8H6miLl4CtkPJIrK1ZSxOfYaiQsVqWwCjyjw9ZF
PAydteLjhlihbG+Qf0gARuQ/fuKihqgZvzD7eL/C0XSa3Wwcxt+X1259un8P+gOZidFX2u+J8KiX
kRFTTA+ImaTtfoYi3GxfOpfI7ktSSN0gUWYIaFWs5gxljT6Xc6yZeDVUKqu1eeQWRABpYJVcQYsc
kMdTVCvbgJvMWrCT8kotM+EVw37qpzdDGk3MGeZ0UxTM9pJrRi1a8iGcF/ElgPIIEcxeCTVMOvRj
SeQ593C62lJqtXPKmLmyRXRI8XzTAgh4gFJdDGYmgCSKZ5ar8ak9wCtpaOqKoCYArp9Spb09hFVr
Bg2PsNV8zxrimaeqEEg457P1IJ6TjHdFPOfBUzP3GU/2A3vEBdZbPPa5zWAz8UVFJtUuL0YlbZD7
dsgQ1qnCXsKGwh8ysd+dm+KI/0Qlq80nplYVvZkkHXIthLXThzreXIc23yBKVLdgnAU/ckIwPOT3
+Ye77QhSEGvoDU/c5ArziLLg4a7I7P1TY4VHwU/FJIh0BrXEiSl70yhKOHjYwbtbVw7bqDdoGcpC
hV46Ah4jyb25DgnK31IWBRZRdW4RDbkzbcsWy+GaSUKXaLX/b1tctz6owMNcwqn+++4DVbyvwjuh
8Gv66/xA9K4+4aEHohEQHYl5ISN6iaL8ZQARTI/WAPEMGs8b9JJDdzWG8+molTfH2suVhs0ix0tC
JGMCHh9lYlyWfEEbj1RJ+vYOOPqNPq6nXcuVtM77aQ7D9wsVw1iM7k5rcu5cSAq+H2Hyt0nznYDW
y9tZtmLwRK7HuWrzwMRZ6CCh5002KsqO2qPNinJ6CEVx2R4b68iOa5JTlSprH9j3xi2rJLSqAuop
BMAywZ4yhpP2eqw1pJKtDpcumdXys+9i0akmvVwAkqHxCyIgjNUP8EAbq7tAABjo6qxfLo6kZq1I
8/irpqUbGjbMC6YZzQV4rjdJ50VmYBqIFt6OIz2GYoxlHqjT1O3ZAjXiIzS+V+mJ1g7GlMcWowKJ
2wzAN3fzFvjTob4x8l77crBBHIF3zxRrIWzmeJ4gmdN9tfAN0vdIaj6EIt6itfQ1anCP4U4x4juN
6UMCCCsHFMDiJZAZxkW0yJHfHxTTfiEgtm9VpqhL+q7ByReFv6vfmGU4tFzahwMmk2HvZTkVKlwP
elIf3GzmP/fci3OUruR/2hIN072VkaJNmbnlKdto2F4yYYaVLcSNXRYvTjPnIR86MXMMkYsxtsLH
UjkW64BBAYfuVCZPEb56LRzJ4a/Qls9D31Jr9teULU7l48BJl9PThstAtVjY8pdJlLYm/uZSIP0A
53buk1CcyIHhfMtMoq6usuSpor48MreBD37xvfIBD5MwRw+TSblOr7eMl6fd2b8iKz3ykgfMrvD/
mREifrDuJCvp6jECp8w92SXEorKTcGUk3sxMuICvCn4w/vh2JkRmL5XvK67nL4oC7xdihzoAIbNU
O6qDYTaiajaeSwZlN2vuDluar9Sy+AytR1Ixxv3JBxyIq0VNRg0ivZRhI454yLPYWSxyw9gSVRnv
L5BAPcp+0kOgPww/gD9Smp46H18HxzVAGcw3S23KJyow6iOnzLFy5poNCaj9A1b4nBNsLre+OYWR
JUHZxEV2TdLNutjprEvMH5AkYNQjnrFNZrCsO7812ysnFNd2V4V3VK7VMXpcdzupiLehm4QSesN8
BzX1MX4cTd5eVPvp7b/hmM0U79n+W1jlVg/Wt7XMyhTQFiz38h82tHCvTPvFivDg8y2QtYBWF9e4
y94yWVsqj0MY2+lUQXZkeTjJjd9JKbWJA76UYkHeDclQbq9ZqufbmMzL6Hawfv4oUBF5o6xzyrQj
6MUOO+FtLObVlYsZ90bNlbi4NETRYKguEb2QaWXEQtahL0UEyikW9j9Og4QyGtM/QmWMaBMw0TyQ
Vhei0kPXq5cNbztGuYQ5ewMqLjxXrB/SI5zi7Q3khufc4sxFT0WPUqe+f7k6vK5DWt/JDpL2VHdr
o0MP3ew6DLp+adaLT959uNzmDZbybYmJJrEqUtRiyRO59DOcq0hcLVXc0nr3O8OeUoUCPA4kLfJL
enFcefa2c6lvq7FG73qGHP4nDXjUX/grVvEq/l3SZUG+d5vOxywdWhj1+mnxLyxkAvucMbExKWVx
zTWdgSeT+gz9h55DbnsPphrzdq/kO8wUsdW+HGSj5PZ5bu+X3ayotPBXxCsqufibu7CSzJHdGZZM
/UY7+8Jv92XRys9zNLUqMDY5rH4xcAcd0W82zpmK5Nys3xBO+1lAF5rtiwPYl0+tuUR+luZS7SYV
AE66rjl2DgC5xMsiD+fzS3LmWEgnLRo78yiskApg1PxevDmr6lfjwMnAJlwJ5cYQRPc0d+sCUVX7
afA7T4PU4JdPVFJaK9MPLnv3iV/45TA75Hibeg0FR6B7TFzTDUwKHWiYh5bGEdbxY5eunyn1Jlua
v5/WTBGVeCk6mpfqnPPy2wpBkipSXxM7IBciHfZXx8klYDZ/eT2Mpn0I5g8zHpWxqefQJD97e1xn
hxbJN10ZjxSq4ojlLYCE6NhfMWRc3/9mDcSRSy/Y+WmFZ/S0SMgXtIT4nSaFDUcAigaSEYa+8+wF
tgd6MOhX76GRdKghYrTkW7Kpurt39+c+PDOkeBvRlM5h3n9OuLlRjzPpHLQEuQzZ0/enIAeI9YPy
G0sGWfT+Ry5P7Xgzo08Uh270SudQpZBeyrVLdXOBkGQqKOX8rCHRnlaqD+MKlpbmpQjNzpAnfeVP
gx0xKGnCDq+AiLUZiO/XIlzK7GWUWUXyyYTTNmm4b4PvEyeBE5Xyq0PDdyHvXT+ULctOaTpQ2Rzm
nR3mmTnmYWnAwPK+qxJnegBHayiN6b0vQv0t5huZQT/YENvR9kMyHxj510rNXonhNc2fhgQypXZp
SCVJRhb72Hh4JuUwfOAwX92+4TQsh04SL/2yRN+yaK5WWVVFbxCKdbdbVNnlTPZSlDZQvV9agZnu
ion+Gqy1WFhO4TNcK5E2YttyVo6HApyKShAmofWzfORsL2dUXPz5dsNBM7WlVRRQeXcZA0uoO+wH
sfa2WIAwAy1NuoCrecVWTkRX/E7jTh8SRGcnLq5kNODVoq/MvoXt4hFcleTTLJQA5iRYP7bv9wnV
gfRBjX95GgB3x7Lh37pfNodWtzZNKjq37qEd/mxHGxzWnZKc0UHQna8/hfvmduUcLtKAuqxd129v
wMzNu0EbwrJGry9POL3SwJMi9gnAMgaH2E5WikU3G9zmoOS6wiQJQSGv6Pv0DllFgAJZca7a9y5q
VyQrZdwjOVgcgAW5fOrZZ0FMsIpE+m01BDL9fKt52qN20PkhAsN5miu+B6vle9t2BfwATQ7+VMF4
PpIrjzK7MRSKNRbTFqdAiAVh2K8h6tNRQ6V4244L0XT4jXxj4R59gAqv4gy/t1tDSzyoo+UwSfLe
hT4XeicWM2Q0xcP8QWi1th+Gkj9AEPOlrMseT8FLJayq4J8ARUI2eVfLU69x45T5XGE499sqp/Dz
e6Wmn7hvYGSSvlde3AIyhZU5a6DA+XT9y8MxykKwTjMPXJwQUuk1VoaYouWpJZ4/75fKsEENsaLY
vzlw4iptuXCLKCNkbvy8C704r9bN4GuOrL+1AKpcb753utpu/ihObg/hSt1LL+PBqZrNGsa9Cj2V
49nuwq6QEVWsIFsVaZ/3Q7yF+x86kIS7TFY2ahnpn0JCU3whYE82L508177wR0Tzz4/+/Zsg5Qy7
+lGeU4U+uR9Z60BWat9DoDwleRyZKS7ykKPdyYJ+/sHSEy9fsM6QK/VfYnf2wavlWjxUSO0In8Oo
UytpfF9tK5XytDryCNa83CHFOMHkwKODN62FB26O+c+Jx1zx2XMwY5aT829LSaDOPTE3mxKrIUeG
fmsMg85sHibV0TgQhFL4tNsecbaVC2mSUrUJUW0016+N6OMIj6CU0ShcYJBD9KEsSlVnBGKS7IGv
zxSfvuqEq6JRv4SG036gG3tBI3qoCSFRa/IdM6tnHe6Am910mjxP1xiiP2qoGcVnDMymy6j0ULvi
l01ri2UdJ3Gq+6EZwFyJozRSfIYb7hci87rRS7ky2PrBbhheA2N9rJnh2n0MKe93xG+B7tBuQscX
yBt4gDNHiQF6S7nOSdAdfL2BD3KEx+/lEpgmMac5ubjrdWBeqtRqVOiJtchk7ACK4wljTZ2fpM0/
kNs71CZHhXixethX+t1yv9Wy+qu3QKSsZLsJghZgDr/fgy51pIJyZWmKoKyuVEyc+ykV5fwcDBi3
5EHXSI3mHwLwysz04w1fcZvz3WeOGGW+wIqo4cthfxvzJZ3TILeOfZAvupDHnjDMc8EQ/MNaUgGa
YSlRqVhBCn7yl3w2xIa0wYQDaFv8OeZlUJTm2J7x8bPxhczTLOWnK0u52pirinl6/MlFYuX/O8qc
5pmDoiup7J/QRZYAHlYMdg+T7xbf+mdJ23JY3pPC+CN8cfwO05rlRJlHV7eYB+IlxTA0pVKsMV32
nVVkpALeNf7dTiyJY63IgC3xk1iYljTezdNfNsUSXAMRuDMtDoa+5ZS/0NWeiZVqUNTep5XaynPD
RQPmknTqem+ftzPmo5Y9jVY3MRIwaY9BgWz2UuLhH2XOCWVFLPBXmoYT9lz3meNYu8+jqwHWb7DM
pbqFir6qcRCUEH9hJV3ogZme1iYaCefTHwzHigNKJAylr3vNmwfXyervIdUgHv9OQmni9ba5zkYk
C7OHzaEWqV2OMF9tTdo7blsyr1mIy4iTWsY/nbgP/p2Xvm2InCGZDbyHrmOBTWcNZKFkarZUmZou
LMsByFKnOdb+PQ0/3fMgiUaif7Sl7Fq/s2lyMvP0wwlyk2IKenuLEhogR9ubguni8n5RPk1O+n/p
kF5aO9ZTSjOzeAd5Ft2nlqAlPmXZw69Hj1U3G41DIs1mXaIiIxGQstqeZpmpsQm1aVgWoan1lbsI
X3+Y53aHYxcRUns5++7H6+MW/xROer1HSYxH/SHvGKT+TGsKwTC9Ml+/FlvQ0S/ImJHku+KH20Q+
bRCVpfp7z/vU8ycMRIwGrtV5vZT/QB1FmLe8C1hSMcHJJrCRUM3r4Z5nE7bTwAgLakAoer/Hi5c8
a2Z/pWHEJWNnB8T5wFZTbSUrB28rvCTmxg0chki3K4w4B1+M3ccWoaCuzKJLLPpUFCxnPESp7e23
HqiBpfRIVn/FoZSy1BqgBgHE88WeCA+XD5CYtccIZ9xdCWV5C/9c+fQ5Z2qGhdWrDWfE/lRVyMHv
csu/QlVur2NEK+vty+h4ncEZd8ZhfUwPArG4DlRtGSadB7lW/cS9+x6lfeGnJFCyZBfq/wSU3qfq
1ilH45I33xPsP0VqYukWwwibfulF8rANlX6uE7GnCQinFWVSGeDnE6x0XXev33/J0E5qwqbhOLxY
ZqudF1Xuql5VApaDcpW3ioCx5lCk0WmrdReL3xWrSbezNKhBUjKwvw8nAWFS7WaoN28Zck/q+a/g
laZ2p3c58w86s0d9LYd9neL7928jC92GeqO3jkc8vo/LxA789T4Q1FB2CoUVztqnkOz0nh5Wt86X
iERkKtNIDLm2d4m+pzQzEPc9AQah+AW/8qvXzezrhScgnIi8Nmq5Hd6eWPvZLFYglGl1u/LwVOD+
ZdrTCs2h7pjy+rOvqBZQU9JgPXM1z8LHqKv3I8ykVf4mvev43Lf9fkZfCKEudSTnEgNuc586bplp
cgBl89Wh8NFnv21RDEpVRg5vOqS7Jzps5lNCJh8Rncd753r826WhbZ4L+5hNg2S6R8OKJau4ZO80
n05v0C9+HH35nnlaINP3/LE/OwcK5S3UysJ6T4rK7ApoUonab7PW0eRiniveWwEe7z0VmkfGIVGQ
Zxgl0aSeje0GYYP3jzYI2XtDY8fYFe+WXq8HeHwHI6rkQCJ50b+dE3eGMt60gR3mgHQNzTVzGiAd
vhm0FR7rj3FuivA9DsjRsoVq5ZRH03ftBhh07WaAdEpjE22cCkbQgFBPvOS86QclceNXEAz9TPd3
SVB15Y57F0UTW1Fo6y1A67grRIbqxJ46yFBfvyNHuagpoZ16us+sfo9o/Hy4GRrsYBiHWxxeopMX
uEf96Ol+RT8c88Q4wTTLiPtmPaH+26rLN6ML68BrAGIkDrL02JJh/tT51T1DBhmOOfzd6iyBv5Rx
6cDic2Y3tbYhYqcNTeEz2Mo0IwB0rqEWAIdOH2w0PqBO6T0HvigV5K5mgVGTdJPptoCSvyGUgtLh
1o6PmAH4l+A/65mpRs2xf99mBE9I2MzoMq9DbO3cHR1KL4BuNQR2fh7XTygYbyoAZg06wTvraaC3
cicIQ85UROxt625uT8hM81EQ6E3n1DLlDP5gE6zlA6A1n4uer4tevjztc4D7tUCcQ216D5ZsSvCV
n+6vKA+3WVPD2bNBBimwTfx5B5kEzVSVYOpiGInx8STc0T43vVpBdkGR/5gIrlaxrfzjYjpy3iAF
CLjtqXAEebCBSvLxSnftFgAo9t8Tv7efftSNEnJUMWzq5aaMw5sPwsXo1x4RvXP3TcUIsTeEz8oX
aCFiaMfRSJ8b1EmIW4vJOvY5MLfkfkwhvSfnmdPnEbVOtA8kj3pN3O9tmQ+3D0xyJq1IIRXswkgb
L03AujtawreosfO6ThWTZNYqewOcQWVzD5k8SKyDF6JE4i57jUQHuNFHbtrSLDn/NCN4GCd9oR3b
fVUSYCPC3JsJdlDLcBS09j40a0iu08rtcGho+54QiEamEx7VkPpbPWRrEaKLmS0oqA9HkBFHKRxA
KXVQyNxiorT81UKmJKFQ908Y5JyyGeg0/oA/zhlGQrIeUjthcOvkBysYwBwxqxOLQ6cDa0lLjMjP
Gl3pKGL8dJ7WmvJIvPMbQPybpRpe702wq1wkxfvtpWEo5IDvka4xbCK9GlwpbYpzjcDhjzNKv0Qg
l8rJg954om8p7HDml6eFerSA5+I0Uf8fOwojK+GauaWZ/8fGYqalYY9KpmlDnrHQxrXIVl0tABsC
/guV68/s5e9Ia/j0uG7SvE4x+fZRL3eh14JmTfW9NETS3Lpa6It+fJ3l0/v/krClFtPueCxD1VTv
wS55Zz0K5fKAtV5VBns84xyCX2t2vz5Lh5NBCRU+Ye9r2GapRgYkT88MiWjb44euxg43mJuKLkV5
Jvyeh0Z3PdbCqbT+JyMGqM/owACcDPT48RaWQ7HW1aTB0h2a4nNohXrlf0UZsxgNjF32ngxpkKE7
oN5pz+T4QfzcevLts9GbmYSKlBFHfsW9qjXgbBorcftDDvi793nzcekeaBncH67QaUrPYzawN89K
iwfaOykYsHCQHaLcxBqshoTdQzaRu8FTqiYvANRkKz6JxgXvRo5ApSCNTUCPSq7q0HiCeeXnAwNK
uDOQg7BHWDHBvCRFo0PaYYqXy7KCnd7LJ0dDXh5p0T6hJjmb9DOkqxKyKmtMtiUYRSn+po5pNdMJ
zWCBX+Bbtwb9w+6BcZMjBPxGkdwS2ZTWsIrxSswqUHGcBc/LyYmFeLiH48DQJdKkcqzV93ltW2Eb
WH7TpjVZGtDqCQae49iTS27/zI487NK4WQYFpC8nA+Bac/wiaVvr6w7pExKBYcmmQCuvTreujO3w
GXEFBeBUMkGKB4TX04B8C7Ra3zpWi0MlBnVKUcRujv1j5RQzTTbeIcKm3Ppke44OjMjif8ejaNkS
YBFgPJXOot4gsGrsKLhSk2iTdr64jaNwFr77svLrb8GMfM1wHSbguvApo+a7G/dTl+H+eiTCIoqU
AliyzdJl1WWNuf3MPxTUyBQEVwgAOJXhy64wWZm/2NdRPPMWScU7/g03RlgSU6I1q+J5Af0PDFIz
RiKFiHa2kmso6hU/1dbtWYNStKul+hMG7m6MBLCHeR8+CDnhSgCm9tbgvjT2Fl+VGbksOtI3prDw
cTw0fFWV/Oqr6je/1jhWgX2jAWRJDhgwDuthuQ9m2tFN23f9+3yodgEz/st7HPCqoga2NStUqa8a
Z1Wx+ZQrELgJy89KuLU+q0PEZ2sxK5lvsZzt4Jmk1K8gNcrNY5bMUhUPqSXPeJmQ3dE82M0BoQbZ
yCwS/uc03v109yfANyVWuv5MJnM0NbFs7T2t86cSVFEkNzN6sjoE39KeQHKFSM+uLLUx32bGzlQY
bTEd/0jV3bbPmM1J+9pR6HN4BcvJA1VlIMRqHvt8NGoty4uqra3vDGZugezeOttE4Adjns3hgMXP
cX993TWEHA3Sej2RhkBcPEFRGdwVrlkURY3waN+5JT4Q7r4OK5R450NNz5Qps8VdyVM4m2SOuQd5
f3cEr5mWlUOY+LTgajPM7+S6Hux4g2jS5GhuNxpN6XTURHHA1cLYNLwg65/FnCRiGmVV1QYNPm2S
FO42D4oeKFfaq2kkzIl/O/MkL4MRFsiPCrB7TMh/9qdldD/7kLZBmOLYQopT5tGMw79+nPMvQads
f8koJ19dMpXPW4d3it4jCJou6dte/ywvwhesDMwLY3PgQbentlp8ag62/SBO/GnZGcuo+ojqY1f4
BPAlrL8Jc6yvEbo7ZYQvC9GMfO/SZDSWgmCKsHlxYF5wWG/A+4OIL/qZgYYRCpeT5wnfuibMr5II
rgYaznQMngDyHozEHIzVbGJn6zUB1wsmAnx88r4aKGAoYygujYJaI/OcGlM3wiqc+7d2LGKdMHnv
o939yJyI2Env8aSygWk4OjKqaTuED7lRwgRapCq4VEoxeF4HSVjYBwM1zVljzN8fE9lPL7n75NUo
xivzcucsulVKl2ppHJTptB0pO93xP41kq1yiKEM453ZyU4La71g73IsREMn44Bb38bsZijbjoA+v
IDqT9qQyMThadivC0h0vly6ZUtB0e0ApB8HdsO+83lAtuG3/UINNf0JtS0sNJMYJGn15YAvpzMRH
0C9oMNOe8AmVw+QXtDmFNsCcjwIg/43WjpCiLprUHOMjDjZoas1PFL7Nbgs0wPzgofHDKJap+P5k
ZBpFVo/lEOY48JIzlkwZEgB+RMKg+PjF9+RKWglaw/h4xJN84T+yr2oOocrSeshd2M9k1OwopSKk
qu6nKT0VvYxcWsDRU4m5DqOhpeBQ8EUfSxMGYOi4DptsJvezUK77rYHQ71St5F9hwf9I5qBIfhvc
q24UxuepRpKBcOgIH6lSvcvnqrvYZhs2+t8jO2dwbowKI0LMSb9oZtO9uJXaSTvtOB7qs3DH2jjj
q6XFKcmgC4SRZOlG4q+luTEkoXz4ariJiFf3uv4EXbtcIVsAWLBjawZdoOku2N9Ci5b+9F9PChKr
ykyFA7AJ1/PYlE3DJ3Y8CmaEPIIVLpjEfQ2Q/RxPBNzMfxarZ8ohNq47tvW6rCE9aXoV1e8UxqsG
SL3V6cjbKMbodtGeTqcxb8U10uNFNhL5dw/dGYU06WW5Nb0P0XT0tU6EOnuKmYKuY6SlVxRbVmNK
Z1rVDpGY0ullcFnWqGO9DyE+QEUyjZlQ6C3yNQGlcAHwWbo3xiuRMfWzjcLo+BaoZzS2BHUsx9nO
XpuNSIgUFh2QHWKDbv9jath1YgcU6VVfDxYYEN4TNjPHy1v3zQm1r71JcwhpyoVcO/Ipg0UMtq/E
KKQzTzkXzGaU6Mzx5U2XUoVh4uZ+Wa/dnArYngFoRPCk8/MikOTvMvpIJx7QOxJZY/ibs69MINOa
SBIzBca5Uo88SRTA2uPIzlZqeNs7wROQ1u0pEF2PEdDsLh/7KFpNFv/LS21C/o2AcQit/LsbPkB1
mxkA7PNo55UFOd7ETxqqKE7aKDhdaT8SdEVZdIuEBHl+Ye73LMaIWEIL4Qa82hvg4VpLAUdf2DFD
pUHhtoiI4qwjmbfNng+emmn91y6nv25L2Ksr7CIx7zdOEXFtLfqoCmV3oTDKo/NDqc3BwlsB4RME
tPINB1GMafOj+amtg/WSyF2Xyk3zKUUK7Fvcc+uvpJYku0WDjMJkp+OjPn/HgtfUamB3+qzxGyND
KpBbd1mlgD/LrCiJ2rXdScUztoh1b+nTgUsZUnWFh1C2W6QAhIGm6zTTJaJBgjCAVuINVAxOY2Sv
R68QlAl/Bju1ToycdFHTQRO8QFc/rvDv33WEn25tpI3t+Ji1nQ0hpekaLONSPuSVLPQu4XYzkpf9
AflXEqoLuYDuqXV3WLvBbFvzDMgViKg9rT8jdNP509SquEJumOxMgIn9s6CAB2j+uqXFI1ea1cyN
CiMgBIZdkOVQUxezxroJB1R0+NOnAThTZwVYc2w214DTzFsX/ouolgx/sNSE7guMoBHvIiM3vD6/
9vjbuzetSaYx6AWlaXSQNWv5ld1Kkz2QoT8McUiA9cLBCHZn/iYWyC6M6yCtaw2Uy7fr78ufOL2C
JRJ3ALtU9NxENINOZ9JM2yv9GGZgHJ2BUT7pKfeEo7V2HuqhPb63epkv7rsYDpThH51gkHhNxZuc
913GXnrFfz9fDFSjA+9q/vOIYVxRZgWdV4wZTSm9BwWAMQWa/beIxVToeUpkD0srWc1KnCneHWpu
qzZaT4C9G9/WhImc2mP2IL9mfcHJTcRbQ68xRP0JeK/vzdZWjCZUDj9sO+WOopaRGtnqBSzCaxHb
ut6JUyaDtOrYz94Gb9tVJPIUxkwdwLrEvInOQQgacVtQAy+ER85nDilMiJGhwYQJ/UbD9uaRZw5x
vzMiCy8vskgLjq3TC7c7Gr375C5ShnnGbIQIMJ2q5fylHOkmfU0+L2aaRonXP/zf+Qskyhpupea1
WOCAoswdF5qL5KH0OXfCxUUXOypAPMAdzdPBGi86OsQIPHSBMeIWaggrvsHdJ1JtD6mup9RPQRVt
jEUkAtMO0/MfaVpmPiCGKFAzFnOxYqZUJrdwG3GbsasU0DPAaorqF95NI/0sjwY1fyy6IQsWcygE
s+BgSplsYMG2ONvGaeUcIHLeq4KAhA1HSrsoC/PqvqW3otTAj+XCsBAnvPtDwXPPOIpT86ygKvnw
Os9COBKPQkMceleZiXV/cOjOORf7VHPDA53Fe4vbeCI344rrkf70rqRXKVL99T/oGoQLyN6q4FPH
NbFB9jIxzGr4l8Ub3Q4Ks0h/su2nletrrXs+cczE9GZ9Qo95NPkWHmmo/PLuBqp210TOTXvuxE5U
mqKZVLnoTOeny7Au6x3KaLIeMnPo9iahrTCUIU7OzLQtZPFRxyjiswhLOx/aCBsKOOUhUNDsIXnE
QtSbzf25s0H9Y696UW/kKP0qty80b8QwiTE24bxZeBQThg4VLNsBGG74e9n5hNnxsc2FPa89MrV6
Hdw7lwjyr/LQ3tgovuZG5wGYBzkeGo9tVbINYDxlPmY+xJoqzb3aQZ/tX76B8CuJfvi5ndcflm5J
mf9v/c5N8jSkn7l2kxkSPPy6Gw1RXiAtwokA6l1yel15iLkIcJTr6APYlw34UwXFZ+9CCV6YY5C8
mJlIwwQU9VCYUHubKJJpeEG4QbHxOvVaDg7lP3dAmMgBYvqgXgiVLB0+HHkmDaQM7AacasU6gK6V
/49kHt60hi+fdpI652cJd7TIFskgK78uJMA5SmJwqbNJu87oPbovK0Ae/1pu3v9lU8RiJJ+QctDR
nZIduemA9TC0IZnD+ThhQ8qSvz3EcGw0llifqo3pTWeMQGTFYfcWYyb1oFwzuBxr/YTDF3X/7CcF
4dO+q94CNoIlS0kgInVCZVvVScjuh1yZxAH6TvYfNWBp7SRfClaAF/mzPvQUpCckFzC7mNAUx/03
3c2bP1Ajyz+MpL0p/RrycN2AVCHg2mueCLtKnPa6DBg2oX+8SQAUPvngOoPEC8NzJLpU+DBXrbw/
lu7PS2asp6K6C+7ON5rejHKyCRxRMekzMIOTkeQ0OGyy7ZSWB/QbK8SMTPGArTATZ7ZRU5JPsgUv
+PJaP7Whf9La0PjRLuhUGGqugyjqZwPkKNyOiqjiS35vShc9JzwpQizvlKl8sUc+9ww6Yxis+WZ2
vshbwPYUwDRQYFgP/96/daSpUtKRZgnR9tfXJaKNLaviL7APU3tXWgQS0m57CPJswBLhkmqWGJ/t
j/fSPYXBSbwxcHuhwEBbbdFPZUb5J17LqdAiJw0C87nH1pepDCjawedZ94KqPWXtH9I421a5Qjeg
x3IZaWXueNbPT+03+QVP5tc2Tu0dRsn/RolOPEJh5b4+WXVWCC7AO67zqtUP+Ya0jnG4IH5ZNCCW
GjqhR0fiVXiR5nIeFoZH1Pdrf9b2bzKIPaT5Kn94XXlctrZMzQxdsmvsa/Vmovp07v8CmMTg1Sjo
z+74tVfx8O19TvmaEkyftcdhxdcuPUx1N3O9Fh4WPItyPoYgc2nJZFV2hgCprC/LMNuBNumH9R75
RcbVg2U2dRq6M/Mx/j1WZWqvajcAlmQlBBoAOGDPOJiOvNrCb8LgWg6luuIx0ygK2/vC+OxZ6esw
xjrI/wGzyC+9IX/mk6Oktt2X8/sOafBLgbGKzVBtMVoJuCn0QNAMojwWSCUhSdMStXOahWNUl4IC
qr2pUIMXhUFxqoC99TVZbBxR1n7J3P7zt0SkKjynKOWkRoBwMmzhMM9EPZ7JJLKQ5w+unujGQ86T
GPe4toMKEsmHCTkuD/HtMMFqmFU0WwrUTJtrrwpDUrcP2EI+AC0gJWwTFdrrFVg6pgtN447pykzf
XoQu1xj2plrCbtoyHlkRKjq4cHiEmKmlr0JN43F5/NgAafYKfExA5nyZlWZNlL6AFmJTIoVqGVCM
jjL4iRvC+Ae9VunZOCh1DmVy7pjUWbP+3JGX5bwF1Lf+Pze9UzypYy597bqWHxezTeikH955gmuS
v6LEpRe9wpv1bB7z0k4cviOooZw3OiLkSNzJm6QDVoheGu0Ch7pdZWT12p0+cDGo0nX37v69zgxr
VpwDQIFg43x6Pjrinjz1RKPqeVuJbHzEfor4KctzwrW38Wo95MqH9RXjgEvRvl4kHQIRxp1yN6l9
D6ldrKlQwB7Wt3csZxZz2lL3Rqw8P9Yz9fNFCQSZ4YGNq4kxuKVI1uP6QiC9lEqkseJKA+fqPurF
8uH1ViJQpWGbbLWAwQQN8msI6aGLjdI97tKR3+lAR0cmERyltX9BwB5NOs2Q1QAOi0j9gW0Kfvi/
AevXW2O26pCBTUxrtk8j0uQ7VAWRHYMJ1A6a93tKxOxxuhNCggu4MmSvU1N6iCZnTIE7zKVBaKat
iCSFzL24gb0ZIAMTWrMt+R0K2rsC6w8lDibHpPUexs8pKMMD4UGY6Tpj1sd8xyQYEwN+O+9w2oRU
I6VJiqvmO61Zuq0+ERqq7cN1jDlPBd8+rNn871dNIXK94pexPkairRH8PwEC+HLCgF28JJF4EfXy
98uXAXIbBICIIrRRb8QNPmz81qCyzsYu/xjS5VoJGN8DPYy3nWrEcw9kBFfYYAGm874xXwmnWbvT
6cqno81J71hjzaGTpGuKSvvzd6F9clXVeAuyCUq3d9YZA+MegjNt+6WfiuK3VquxyuPCqvd0LLe2
mQNLgW7XBzIcLjOddeK7uteu4W0siY9xinsUVxDUEUXeyqDZTe64aO/o0rL7LpxkQq3fpnllH91Y
P/WBUeJZcXCQxbEZsS/rmKYrduVbym72x5NvEPq67iUSFHqsFDkYhuYmsVbhDIvfomQM1uKBH+lp
nMMjjDLH2hVZm+Cs2EhtiQ0uIsogjlAThEo+S8x8yyfzvTNVXeYw7/lCvJHcUTwb1TZCUGMLL44d
04IaWmfvC0Utq1pYHtCn7n8FgISyvbBeQj2lonwc9nVE6B2Q+yYhJSz2PVHhwtMTXBL3UBwxdaib
PMHsf2w6hHE+LBXolmgcgHnmfNEEXkiXtAZvyw+1508UmkyYvJNRPGNx2/N/NTWJ4HIeKdac3AeV
8mUWRAoYdxUmEkAsliP4q+5Mw8WEnzWvySIDVkg5/pl0iuAIUCyuUwo1AwdAtzuDlO5t5tKE813t
CL3MnNZnZTSObaRvvaYWptsBCzkjL+g0ONwyE3buRg0qB1JkF3qmMW5e8hPysQOfGKT5ee5+9zl5
jHd3OQ/EaJifkfefJdGPXMrNAmSZ/il9sBSr25oHtXJMDZTmAJZKJfPTjWvT617VDOWiq1XkFpAe
n2aLYjCmpbDOZEHrdsXH4NLG/E3yPvTc7tudIr4LS6BZVisPcoOweUNdbaKlIS6eTEVMJDwLKzvi
m8wyW/NNU3DWWlGxA9Iu1meiW6lNYXRRbsjVtXGaLUbbZfNnOpTGQXdJ6XApk0IJbJ0bPJEkjLYY
4wZ8dL0P7XJAhVOP5KoYSEabCLHHO76iKiBIxLZ4ZQAyhlPu7hzzDNpsjsaz2aHg8l79Koy1xljL
+Vj0A5g0YTstHUa1Ms0I0HMFO4qr1QPMeVIaVXfaSiLSP7zUYSFW+LBjgqJ36ku/audpNEj/GUY7
+C94Z5+bz24HB2tJvPNcyP0OJyAvIkf0j8DIbLOlT5sCDOjOAyCIphITxzXxaotwjo2/gaTERGcZ
cdsUyyLpm2/FoaqYo4Vcxx/bWAZ6jN7aE9dWuOhq7OQT8O+7h8gkwsshJl7U66iU5NG7WR0xBjnR
OMRnqx+jPH/wpxuPQBwER4MQHG00QxoHKlYLYn3RJ38mTXRb9lw61oxi2lDukzTUI9z9+tz/aZn/
yU4H6Olfu0cQ+IhkQIWOs+VtZ+3/kh7oXG1/2GL8bj7R+yUzbb/69hRMIdUEPyaV6lxiQarldq8x
h8JPGmBwOCznESQRtwEPPwUIjQxdJrG+IyZJPfxhgzfgDHvvyR+ntf5TBO52WUqR5gmWcgpS85cy
v1kecT3yEF0ZfiwtH1ZV3tZK//hTOgNxZidOUIjzuEOWR7jp5w1hopvID5XzszAbuS+GWEI2g3xJ
K7XquXKBkvMgB6BY8BXffTjMFIe62GcAJvSgJzHZTV2F5p3vPuf/Hqq4I0sJ/tnBmqdsla3A60rL
26LT7XDH5bZkRETuR+z7WEAKCBsO6g9lvWViJ3WiUKLc8IxnPLRvEIYGMXFn54PQM8Ot0QDegck7
f8ULeGXbtfJmJWyDDQL//sdLpQwpNpqZlCl92oaUnTIXaj1wY5v1ZL9kyIG/DEgFKRCkYe3umaJ2
9irERl/w8LwmvNDlcq8xKq1Xh23/+RbfsUN7cGRfgOVjhQfXzh9elvQ6ITkPXHUVV85FeBKxDo3J
AEn3OXyhRC0bNY7sln9heoQLjIvJcVgcojMeZ2AHdzzyjHZrJf8DOcgqGwiEjOreN8rNhJ70FmYI
BiolCQu1HnW4C023gA/ABxFC8mChWr2GehRXCFsl0v6Yt+gCL/tuZnTHQCXbqv01JkMSGdyCXaYl
H2trsZ4MBpyoeCjVo9xTPoSV8pIwxV/brbJpZ8n9gGrf9ZI7tbNUk+9ZUEIu4MJZIho+M/wF2ngs
r+kFkI3qWOEaf4wh5O2svt2ENSvLb1GS6WdO974Y1v2z+QRV7nB18n7wAG51W7zzv0TJfj9oIMPi
jb1EWMYtRLkm25CMl+VLtmKMQcPWArI5Wo2YJTofI3L838OJRhp8qDMCzZAlgoQeEPH8oXnbz+Nj
JqfQLqIgysPJ1LK6eIYcLrMcXUg6dXF/Szl31q9B2oo4mxZwqaYBj7c5ZYCSclAbtmHHOkOKqxqZ
FaEcX9FLB7vgBf9JDYGDgxYjXnO59nzW/bSJlo9ZOJXiV2CXT73ZslvDrBREEjrK0meERsniv/IR
AfmKw8OHALI+gFd99XHh/BAMdv9GYmo5IGR7zoIZ2AbPiZEukNs+TJ/DMihOlARJ1mpg9TuX6Hou
GJYD1p2+7fej90VjBsUshSvbduDZZUFC9RAVnKv4V7bw0mhsf77sbCsZnT9Unz6IE9gY6daxQ9bx
h4vhC6W0rU25o+SPoI+JzuRREn/+z0uSgBdvj/Ab6ihUpY0SIRrUJUqLWNpUiCaTTyAjIqfTREiY
kT2X5fujZ69Fko4KvXe2X2wuhyYMTs9xVhp1CbVPzrIYcax1kI6jRET6htk5vQPa2Nlpgk0mAvJ+
P8bOROcrYiIMfcNZDq8SWo23oETem1p9rIcrAW5u6J5w0wZ3Udl7nA3LYrn1U0uLouwlNt8Q1qMJ
YZQj2bsVgg8kCmlsfnZUlGLy4rgpvD3w+wX0aWXD0knlgPvnLbXiUxHsQHfJb6fMgciMcAFwzAd8
P7tBaEWKcpnTPh1WY13aPVA0fsXnzxAwLpbaEXvN9V/cYDL1iAK5zfUvx/S/vgBZIR1SEgmzZP7c
lNynYwx7l+fIjNtUK8DhYjez5hitAOB7meLjygdDyPDM+q3o/E/N5PnhWXU2or0edBwJx4KZPuq0
37hHqoPq918L2I9701ORsX/2G92dMtd9mUTWhLT8vHjghp0hHZSuXmYXbFfYg9cjJ9FjQg2R98P0
DmLbPyR42x1lfDWYwEhbU6vbm4mYyfzoImNkwF5tqlFgaSmarXXOrNc3NO9IFqXY7c87sEAllqev
if4eaK3U/pSpyzt9EnidXNHvBYsHKKwCSHBHC3kd/wnuuZ3sujUz+YnoLj3Fkw6O0wPbQ7misxJP
OdbWrVcYN53/ee3n+/O52u+4ij16h8K4Q3QLnSxj705DNODE0RWpzRPp6JtyDWe1tl9Q34YlnYeJ
NjSfB3bWHV8MRB4OCAZwReXCsB4cPFm7vCFHJDAWmrZKN/OdrOoVtAWJXe94zG2T2t/ZwHO9Talb
YzpHr1PkR3QIUi0nboh98o4+HbUqktO5vKZexrKpmhsvUbam0hAeprgXL4PCC2KmD+QN9l0h3GHA
iwgcF9QtaPZ+kWplD8GaVIQ4kRVlz3MnPod330xB/BASd4K/vS69TAIbCp8ORzduQtFFOyrApToe
1DZlh0MA57lomzBdxmP4hquvpLW/kgnS613HrV0WA5DXuQ7bpysomMu4OVIj1WxZu6zCcICzudrn
JafhFguD/zH+kpwQ/ltbxyjZKcsY0TNYyPElB7sAcBeUIv7mjFZdbzBFjHgn/g0Lm6K13+WqGfdq
gKHBLdE86aq6KJ0qFqvTMFMKNxQHz51WYcDOFEj5ORQS7sSGqtv0Bqmpi4NDhXOxc0sevFU1pFnD
NHmofZBJJDtbAeeWqqY6t0FmN16kUJIJlNMoWlC/fND/9WIzU/LLmQPFoWfNm0jOAVJKD8jSLEZg
2TW119l0ZR3S29kf509o8LOBaT3uKjboEr1Q07pz2qQQh16oWbY76f8oOzAc+QxftNad3eRRGLhn
dUYmyNGvdYbquSO/CA+p06dNvKK00q54xeE2jXCyeUj2YQLNrqTwMWR7XR712rE1DI1JG4tMDxPM
Cw19uQzvsoCI8oljNzNWtELAFcjGeXyZJfo5LiKHpKoMNAG6EGOCo0vWcnSSlGToiPX8LKqSOwiM
yi5Cp+vMmOjYSyxKfUI2eeHzG8mN1epTPd9uPDve3fbpj1Lx/G8C2yHQph1Ldx5Q6Z35Xszx4yHd
3csWUwHtUAPaYv+D8Ow0JVWTBm71sUQH+IJrtt5uqJ3XZmGnXl8EOGzpF0jh3Kp2KBvt+L0+9iT9
npzvE5wW+Oad+FdLATEp8PHLxmN8ma2Lnyz/CqX4/Y0Sx7ss5io9wGLswhd1hxu2Xe8LZAF5iKnY
8ja227pBRuT63zlgQL+ZTnE2lqkbE0yDSzsNkIc9w/qEL1XH7/97WaY0hWC4Y7KJc+Tk4ONUyLMa
BaXlA3AOFwwQVKvvyxTXDqz1vP4/zuF2gHlc5EdDPLWXIKJA7lJM6+nCbVk97GrY8gH+ZV7BAc67
QSYr+RCIB47orvgeuCuvQMT+ASdUgD+c4LWvhLijyNEs2Y1sq8cQLgBLGrc7MkxJlill7cK9C2PE
aKccUM5XadCH3AGLX9j1dlcqyoA4oRARMPqNXrKpRpzOPa/M9osIiljiuaY5rGuJ4sVyW7MDVQah
IpjqKntNZn+NxxEtafP+3aMXeO+APdDgF9zoyawy5wZgwM9+jlQWE3V5IWP+B0t3lw3MRMfUQG1O
vmJJnmXOth4DdA05xoybbimTukYFrj4plqSZzQA/rKKgVOzSsvQ5eDB2jBYcxdcwS112nP6zGb/O
Vn+wDTaoiqnomajsffvwfEIcm8Mj+VXAprtP9YFTfryKTjIkikt1qaQ3QxVImyFYwTL4CqAgq5ay
C+tFe+lCppO1rsWjTckGfOPGa4DYpWY/cTxoAP5fqJK4MqefAhAq+l99yHy4LhA5vAumsgphcEE1
jIx/Q2MlUo5XNrT3h0e1DjJkMiRO3fqNFbbqTgRifiZoCpC3tJ7DqR3v1ZCd6GoPBv8nv9gcegCO
ClxpzisbWL9RjJwCqoIu4vAREMQIAZd0UlFs76Mxq7p8xcsJ0tLuR6kRFwP3uL3PFAZHyYy7tNY6
PQqvU9unNpi+ir4OWPRO1yRZeb+IRGZD6EKHSI3RB775QU2kKoXdqRAbbs4ZCSDncjWsV37IyA88
fnJiqzo/XvCSY/sHJfPJ9mECluBnjc0yjUEzkZGRNnLNPGnZ3RPs6DwQwh6XLHr8YmxUQpceJrf6
1oP1taeNZVanNoYi5NC6XEPuohFOOHB06Mlt1M+Y5iBcxSP0OAw6Cv9Qrxf7qq4N8szl82TFkBIh
LdgoHsn2oqV1Xh/FzRCHDCCuIgu2PCt7d4Ra4kQnUY2oJj4o2nQYEZd586kfo4Jn3+ZmAemy7Wp3
AaST+WVASNCYW5iX852zRTg4zGFzmR4u1m2EhwaD4ak+aZAUciaA/mYAV7103xXgua3fVHH09nks
DywAoj781KocTlDl0m4Dx7TrXm4lccHeKCybquQcmtPFWdka5N5KEw4Mvssea4MJGoMkjfa9oVyo
SnLJYxdRqOi3PTDUh7sb/cVRBUzpv65mpqZBnGhcIB/v0yHF72LplBog4hcDYtYdVZAhpOOw09Gi
O1gO7oO+fi9bpT2Ruac9lnFz/Q+WPP11I638OQJnwDhaBF/jBEa27s5tnRCVU+4JKMLam/oxf3LX
4SItVKk34nDXicw/gzhnhC30sTOSdLCCJg1y5iDTj7JUnqE7j1y0LHnG8WVdRusHE3M6SqwOd3ta
R/Iuto3AYIK39pzBb6L8f8LJ9kq0y2ivD5o7IYTUIrulXuKFjvP391YtvNMCNKCJmC8bVSoVb6Jp
Vvu7JzG/AgpdYq/FVp5LpK6H4kmqf+3vmdZFZ9ZUSM/lhy3nF9l4CjVZMf49yY/h5pJ2gkfZNVBv
EeVuKW+seMPPT+1g0lia7g0xHRqCgl/j1N/vBtj6KWQSxwn2yk6+tcpFo0tn7UT6tUOLVsoqra6c
XqpMiksyxrQdpVQS2P//13VyqfJuBoYAHdynf8xB7/pMCy+18J59WWyvGJqIG5y8OQ2hmXZzMifj
LKe4lFx5MKl5nRPCRlxPhoXuz+qsEcDwPoTrmhhuvFUtEB1kTOKbidtp7Ni1wbtl7G6Yniu3aGqv
ddWKNr2dJx3R1gL578/wi8OA4dimhN88dbE/hmdNWxkZbMXRLqRTqG6SbAxGqqNH3a7+oFOlBK7L
Sya6wh8HdzFP6Ai5ipQkN2vXrYEyNSXOcowxLi1MGufArf2fs3GWiRLwnDXZ67JZo9YsiNHd+oCA
4dKDUdnY8nRHD5b7pcaxLC+jrrc2sLnfET2bWDT3lVJ/p2+6BRY/2g8fKKqpMQxmSeni8Y/E7w72
v4Ik5vjsnnZgxV+eK5gkRoMDg6mtc9CtHUiv8va6TKxeFSWbgU+4koVLBbwiNNIt+bdQTyN+Z9/+
2gW/vy2JEbrVFb+6gFFn3RpzWn2nchVLQODTSfo+nZRvIYMgwBXvAFSm07qoA0ckINofCIEt5FVL
TblXk0PXCSz+RHoStapivnKLYxaQtjCvxORafaaWYyWHtGNcY4mWOGT6M4nTTqVgOCwZunXFAmS/
f9B05qjj05knK7mR7m2eev4JDI7uGrd2DgEi5V57YMqq/RIEL9mFbyNBVu5x8xy/ASIvbjQBKYEd
oSlPr2LM5R7PQxUXdsQhDguYZXUlQiyabFThfHMIdJ4UJ7l0pstWYhut982mlECMqjeHdXxgOTkm
dWUvzVVUN6RsupLTRT13tP5O1yLRzU8qYBMV1iZ4fa0UujcbNcUtvVtJmB49yQjM5JWYlkm7NhMB
BTaL+izwDnMUVsXIhKuPING7LQkecILmNYE51nKgCRTuSo8s0iFjnBbmNNXnhvfp/oSUBIiMv/EY
Cp3o8ag+zOJnwjeC2mqn8h1hSoYMfRQx5Vm3dZRHYg9YgATmNs7ZKEzlaM/4AIHoxgfAS4qmBD+I
IrX4GFiY7Zy7x7BQenrj7i7jnWNIQo6omOICjMDASaHXX3k5SDc7OH6Ttl5EvDWN2Mn6QoSn5NbA
H009tPntsueoe72HqZZcq6BxoQOTdAVMhEDOVEbLplvb66C3nsdP0nE0OxSpt/VZvMu2V5VztKSy
dOZish53DV6kMAfrvHAoJ43H0NL4B96ebJWAfNieW7J8T18KnLKDYuKytWE9XqzPKVDUYq7hiPIC
/RlFhexMJqeRFTD2tGKjRwe54WY4oFZtJ0R+58b9+vNcViNXgPmh5aSfx4DW5dbHxbSw27kb0n3+
q8MEIvU/CyJLaKlC6qt0Z5eDHh1HXiCYhzkeyaudzexAMRisqPNliQ3J8oP84xK8JVfIQkHJ8i/m
e29kys7vOAqrWkPD0+VF241cV5Y4tqpJv3FHUNSERKIGJMD5Pqf6EFuL1zUwf6+EgwgqHuJP0X7h
g9U31YO2sD0xpYUCa+9SRqwG9KnuXKVRIOJMx907+LWz5IF1ZxjdaCNpXE+Vzzh5K+/5Xe9vg/GD
ZNkAgPzcXQ22FuaCmEHroF2txciMP0/I4LsYlwM/uSzv9wzdDiIZIcLbOR7iQYmaxYyzYh9heS1D
0S4Fxa0RT1pX11cKbtIPHXqLKI7laAKetYSYxt2g+QDukQ6TT0jsK1A/a08jWAfq41qGJMFCwkRd
5SNx1vNkVunyD26+dKmDK0cMT6uKmU1+rAdGzZJdfI3vRaqWd/u63PZpegs+SGZHQZvWCWJJBZ4M
EkOfa2RFFtps88do3g4HsoFoft6zDV5ZOANviBtsyytlWrlp3aAMg9K+eDL4WTqISgTbVBEq9I0v
hH6PjJ7LsXg38R5NbMQdcKiNIVPh8j97WY2Nek6EB7PCRmMo0l9BUCVWWsxzrJB8ODrIvAlIOZJE
CSbVJqHOY8epNEurePqs7lHX/zEt4w09sVuT3xtrwu9KveXtKH36TDKYgbYiGCvzAJIBWrYjl3lN
f9sF8dxhwcdfkrCMDcEUr1X5PMMer2IYXYS2hnbzX0jSA2Es8COk8a1AUHdZ9zhUJxV91Qmz7fvF
5CpEPISS13L4qcjtEtwVmD7SdjnlnI12H4/GDkhiAWw3pF9NcnAxeNDx1zJCmxb2UijfoDBRMhbG
IO4eaSu4aX1emqix8h8+PXULKPjiPhushV01/K8QgvzO4aqC4tdLJD3LdORTDAKu2kRK6qG1Rjb+
8GQYGp2og1he7GBQQ2ofovSN/Pe+89Ad9c0OXslnan/VnG6cj05jkm38/w3wn6uxulKNmmKp0GA/
IEXE4xHKi4FmijPqsiXSGlkanlJanbcQL9+C7UAAQBhli0+RGGMp+5Dx8guqt6sJ3wVXpC4E6/Ok
70aTOn8msRHHWuhS5hSv954hfuIlU4hTi5sGlxTly2cAtB2VAL8wPqU1+hQcCuSMQRXwv7PPPs2N
2zTwUgOp8/sN3rIH9Q2zZ02SDxPt5Fn9zD/MWn8S5ylC5PMEZ6YvDUZpaAp9RHNaLkikFNCZb3sg
ZYo0ViSgir+Qlwwn0WTwrlDQzk3LWB+ipetrnEqvtWjCfBsaY5Ycq+zy7PSkLcvLqCz08hJIygcA
SJEFl9MUB5xdzcrL2DsFv08uE2ruxkcL6QUG4ddsXgR7IbvtJaORdZsI8cK7gyE4c1hye4Jf7D/7
YK81DIR3cJzhalUS0K1UEgwZYMG3/QRyB8wR5OmkGEwmqEM8eL62BsO5jiYPhQMK/QbjqfcLS5B3
cvl+VbN1g8neWgj0mpIkQYrLVo7jV+dL8VE0gzdxvL4SKbscMNwhzAqPuPkLCDNDF/lYqde59SvR
RlbQsFFEe/qXCOrtMVordJm01jFDvKaGBpDNxNKjl9fIm8XBZT2dJyL7YyELL8KGbFa4sBqDSRI6
7IWkMgVKBba4EiZ1Hl4hoZcdV/SMVlRkfZn/IqyxwjsFBwSMfEbRGBip70IbhBcdpIhaTKKSInB7
pqUofx6Twwo/usnBpoDQtChJ1Iszjtrewd3KmLwS9BMb1+tKsLgubQX2wnaVB8cmzC9UqhVZSuJ7
YvFcaVVCQ8QLaBo0x2qd96CPtiTzKTqAf7lGl0MMc8DQHgNBOxtGwO+TMCCfYi7bVi3YTCiyFhy8
rDrJb09rEMP2gbllPnHcGcmqqRNy+rPCBxQO14JZ4uS4Cl7dxkEuyqeMEzO9O+8UVaM6uiaJ1Fdo
G7l67K9/X3oVtXGAQydaZEekUZgpXd5EAByn9uC+7lI5NhsF2G69BYqfAkpGErTk1um+tlWMczZ7
/5DB4xg2e/wOEck3fgWWSY4dxPhfNKiE8pVGEsQQ+vtZhkQvlGYNRpMAhcG8QcbKOcJv8SOcMmYw
TdX87PBzGpk1MDe9t0xxSwWQTO7+iEUpa+tl9QuMiReZGtOgeBvEOk1Q0kocaywDAhbADt+f+G/D
Y47kQuiGE3lmN4X5t5u5ywGKGxLmwbTVcHyM9RKyWn9+/PnBzmH87cI13JBCwZkmsLqiYorRa6xo
q3lkXi15K1dsSsYhYl1zTvlhXwHfwEahM8v0847ry63j/MN8Pu5wht2hD/18YXV7GArtfMzMfxB6
o60BDVIdffFIHPkDnOqBypqU1G0Ndp4yNO816fMUEgbBClfwr3N5hJsd9d26/r1n/Ip0KJ0hOePK
0s9d9CT5dnSOUPUaLfjfHuYm/uuBKyB5a5KRzAN7egVhHc6ITW+67vITYYXIE98MKrqy/UG5boIs
WKHfg/jSjBen4B1/RxrmU6OmZ6pHt5YpRErZk8m3ywsb8zUXM9ogooPWa5okXQTC8WxzqwZUxBwf
+yKuxYR6XYNhXCGFOJE+lzN/cR2ilh0yUbXtzSBdrgg+exBtlLaqUfxW/p/BGXG+oE0Qh8NE0wn0
SbOT6WU8RQxOoDBxxHeTVZwzrv6nuJvQNF5WHb8VhNEvnRelLU5RXzE5iAJq7B5fOrW4NUuEXDiR
sjsPTupKHfVJNRiVqZE6R3VLZk5tVE59zs7sL8+BCN5KPFPrQvQDL/NThbN2FWMLKAkEeh/G4vCk
vv/h7VnZ009zHnj8OPIiSbDPcofDU+ULqSie86R7pQFFhT4nwU6Zfq2zF55dVKSSOPWvdBAQT6IW
Au5CcgHXG/EWCyJ4NYj+J+DdI0oFsNESqeWUmqmFKKPdgnx02XaLyscQ4Ly/1UPHLS1Snv1dWpj7
lZQwJ/rHwGjTGwJBeBYpLxUspq/U9pnzAhpDoRkSNEPfjoBZbpSv68a41QzGARYD/EN0YHgOGXSS
z7qXA8Zoxv8NoVeQJ9Aoa0zkB2z8OowOUJpwgDjZh9h+9LTvABhitv3kRHXpg5aJDYk+Ve47sOwX
4+vvrY5D3sKfmST01TEA8GwZsXVgro4VDwlWdEMUl8vPy62KsjqPOBecvPozMBi36H3l5z6dz89M
WNq4FxFG9uE+pqQzQ+eNHTq+GtoZXi4ECNkUVr7MlSrcggD8+LalIzbTGGsF0uqU25y2oRimGmIZ
VXSilMQ8IOGViaeqHhhD8c3X6NU3bMF+sTghGBlB/JM5HN8OI6YpbBNTySpk6XI3rblV9Lko7iz3
3jiqvFAOY2n95LhjMc3LpAmbeQwybNn4PTrGKwuHtDRQKZF6YJ1ReU+2KaPluGBi532QMthgt361
uAPquLthZqPfEtnBT7/DXRc6zGQbpIMK28LEpNTCfwrJk6DUaAJ3DWP4eD5kzxbDTLRic94/JX67
7vHIOeq7XHUiynT5rlZOwCGcovPvEcKUeNtqjOHZRb/ICdcVotVFTPWJX4DZpZ8p23DFFEyGgRWd
IYB7Yp0vSNFXgT/41KAGLbFHgp2Lx0dNFifz2cIJQG7QugB/PEH8RpeDfvY8X2RVeSbsh9atyRG/
JGRN1XfVqK8YK8zAcadvpzhXRzrGJpJQ5WtbH0xyndu8dDg13sHp4UlaPfK6xWhgwNbSuWv/O5uV
Lmfy4fwnvbhJJjyfgvIDZ/DhGdGCR9fNkJ3K269dy1qfjJY/XqxQ+g8KOO7zkCWfgAYIBFzhLvH2
90dJ+dZO8ngSvraaSZ5TRipNcW1PinFNsiNx/SvAz5EUBdSra2aeBj+jfmOT0Nzx/VYVQXz6A6GA
Nu/TowfXY26X4sfH3kPpz0Bp26+eyuGQEZlOd7oMbCUh39vwby4+ZYy26gtJgGVSKRmQ89oMh+cB
sQjjuS07G4uzbFnL4c1duwxbinYFBseTp8RjXti2fWrfCi/ucUpYktirR01HozC025IMLN729cw6
g6/oX7gmzWjFO3l40kgG9k219WaoMARfWg1ZU9SXjF1UD4AeiBWZzdnP+6S8o0hn6dirKGgrXSel
kxZHBAcbbXK+M3F6FxxeX3UhwEHVF94/xnXH598Ea1Q944jZ+v/WzdRwWhW6nW8GRtK4WeUXPpHH
3VB2dgOJ6lkII1w+ioqH27K59YXiA7e9AdPWNkSah8bf0RDuR4cLvHHO+VFMf8NfgIkKeSvxcFSH
3+lQqsueuoH5yVqRIbW4dNDLl4epcDsAAWCeRYkzKIzNKz0EOOVx4cdSdM0FFPgUO+o9bul1JSDQ
C5Zgwki8nrCYZBK8S8YcKVdmqchhmAXISxUkRNpMoV47eQM4qVe7TTWs04qXUhOqy3kYW/PQetKe
jU/nTK+fZg1MS8Ys692t97buzbdYa3S1t+ByQrvTCzNo7PPEaZMlVNd9St5bniFCJCA0bTUEQsOR
mpgDbsmJEJsTmjjSKXoYvEGTaebde9z206CTHWGmS9EO3vxnTfzzG9h03/Q26YTIz8BpLnt/Qvie
1tb/zUbzE1rBDAtPAOIo8USXlcvw/I91o1sVB/lwEjv5Rr88oC1+FNfPIJIhz4xwa8Z761l/H8jB
tyTVyymWCe3wZArh5euSZL5JACvtEo6VwoTnQ6uongBYmCsjaY8KR10D+SdR4+p2Tlg0SA3o3ZyJ
o2wybyOHjs99KFEEZX9K9QaeoUwFDoJoGKruAgsMR2a72gbTe5oBlVBzs1JrUa0Xv2kDFQgGo3Gc
p9bSa57bqBiw/IYgi4WMBe5Ce9aMJl3L3mS/H0KH6x0Kp4oYJeCS8YJI+swDl2a6ly04wdeXe9O4
wIZtHRt4P6JhyDVCQtHNn2uQ5bwG9rhD2h0h1N9nwvLw7D0Yj1tGyXKFdbICpAQcdjm6yVETZsm2
F89sHHuKIVT63gGKdUJe+F3yNcxlSiAyIA88Ioy7uflQPfQLF6Rb9PM0RH8mqoLpS2xHOSitaFOT
UGQMsW42UydI3vOvnrOg9YBngH1frLjUZLvijO2PPsUiR1m8VDFLcJ94XjP6oYGTTvjYw2FKBGd1
ZkndyeCna9X9uGgrLJjGgwroaOSaWMc8CswdT5bPbND64L7OPFzGedb24zE78FHtC5fmgku+N/de
ElX7HXCafdWNm5tzDTp4iVwwAV1o5bK4TRXdNPvHdlGqS/FmKKh9xBV9sGgEy9JJcDVgn2IR/PSo
rbjoCPv2miu8Yx+7UouGBmlg1jgdfQyjSamcBumY9nF5EeJ5FFcLHVPl6AFzardEwiTR+65Illli
QcG6PIZ31IrSTlRJaTwdt9b+mTX1/4GEqwHm+c3pqE88aHyLh/717fQeQ/w2yTCKaM/xyF289o8j
v/pHOiMsa45PSzbpVepXKBamz04O+qhr5uSlwMxgAC2DEM/jCR1e+x3c3Kfbgulitq3BkA0Bcp3Q
3Oy48YpiVBF5WNm/HUEmPxzdCnuva5WwLrkrtq1XlQBvSiiZqgMloDz1wUzZ7bSTdpNTtj/9I7Ly
qbVHIuZ0QYCJ3DYG1kw4gzv1sbRTstyWVr06OlIca2ooSbZmj0sJsZ1icsikEpdTc09HXzCk1GwH
DFfdOJ1tFm4r6SNkjlma3ItEpe7C2kuJWxVA3ZmuLG2sGC52+qOhjEkikwL36Mcx04/jPzK/sRYb
fgwY5KUOBO+F694oQxj13pjwGNbv4S4hknKQI4Uvc0dr6X9IMYKQaKW0ANjQJ45NcqfnR9NQl+oK
eEHUzL+xdXB5YTNAshxR4l0aVT8t2F72QZqeRRnq0bFMl4VbIVS7KUvJsjltq+jmQB0t7abU0xmc
sTYrVzvVFaClnsqY1qjAZZpLD7RXBhQb5YSR58mmdvo/4p5CxRqkMPevIpUqhVTm4W64OaIlg5lK
Pg/DbVaxYZ2z8BjIl5toMF/FTTrN0sfKL9X1Iae2eV56mjSK95diRuBMBJQn6HHZ112m1uVbknu9
XssBC4kosUXDATfiEvcXE4RLXr5TIolCMd5azQnUV/DNMgLjeZ7tlHTdxEIDtKvhEpTY+r5UE8/S
RfJ4pL3yXgt/N/IwgLLarJiA1eyQnhCv1hYysXFlQGB0ymB6mc2q+slTavgD4DAK4LzQqljo5aRa
KEvl4EljgddGKz+jYfIL+aa504DjKUMhB8OTkbGmT5/jF+ApKz/kOVFY5Gzm5C+4Cu46X+ZquGC+
Q4wYR+d8WK7e4sA30g8Ws+X4fZLwHH2+WIwnABVrEIiWhaDqbmsaIVPFWRy8oXNWC9osyFXmxaZe
rSOmj4q1eZRF9aBhdCj9pLqNcrxNHJ5maChRzq12NFJtnpcYFrxbA0IBCILSFlZ0tZ/3tgq3Nbxy
pVVzHvjV7FgGvRzFzHiF3pwFwHCdAuhkhwx7UnYvgUV0nNes7HjaPYaERdjgcujK3En1cmrby9sv
CGc22qWrWfCnKfjgpGLufhvMb4fBl7FXfIfWzsPCVeOaMTqJLFr959We5I1G3JvSaDuxTJ/kntxf
wWac+rkPzS/ZAmNaZtXP0jNcBRwDrHmzY6pXHF9QBrWR/J18BdoVfFEIpQWVR9J5DrS/SIij1173
rlBY5tuo/4prP1D+YqevkEV7j1/MrPlo7lj3G3u7N4nCIsHbxfy8fBmMMLHDuRu93UJlPKB2j2M/
r6oI7aZWoBlg/6S324MtJzoy5AkkvZ/U3zZBR2nCfeqLFWeQNb8zapRSo2rQKXTikPIgD1yENK+z
KDNNeDwmOv+Dr8K7VWZpntWO7tYFxzyNXkXFM6pM5khLPQATdTh4o9Bs9TvR8R/LNV4ldkNO01dG
ez+nGVP8v0KkSx/JbBz66dZX7TBovn6AfGZuFJ2tGd0ofmbI9g9D6Ugbt8SY2qTofTT4JQYK2YVb
J4rC2gEfdHSyII6XwL9L+DAb5LLlJFNEVHdm1B2qlU+Qe64qVFZHgjxV7LwyFx0zM7R9DNyWPGCp
dIJgpSs9NURofNBgCjvHdn56rV37w59lRl3ho82w5HIGZJneEr8R/wVHkujI+GyGkv58pMVQ1hg0
bxGXcXhDXJ/H1Rx0NB+oOny8qVEmH2hlQMWI7Aud1NCI4eirSgJyHTpClOfK9Z4UPK5jCfcb1uXd
64TqALtl6Wx8HVm74Poj5eixBh8mDTagOWwdZv3bBl+MGhSmj8UJ0zkdD9JFPT1iN0rvcR+Lkr9G
EuBn9Awc0C1ej8PlyucZU4XPvziVfbuq6SEJHDQpwTRbD+GGHdubd8NbNn7wlOu/w/HfBWd7HAOX
2oQBerEnc9VlXsKth0TVLtyVC86rH/OJ7c/5c4FmZOeUUm6tfHkW+8OPhmVcJbptnYUwVZ7Msg/4
ExcQt9YqJ+xWlHVNt+azdZUXJDe01DiKXyCiMKvGuQap2rReOQHyCsG9QDojrQZQNFXFYnGaKoAn
lb/pBYL4yPOO0WoSD3Ha1UL1lXUEXhY5AwXAhvt/37gDCANfUkR+MWPAAY5ZMcW5VHXNwbfywljg
5dyMZL3XAXjD9OlcZkPcvME0LZuT2Wz6dLfHGRZCR+BdgLGsagbfVbYTeZAxX+ddLQLFekl9anzE
AtvQ7QY0dkGqsGE6c4iAwp3SlY1CwmIy3rUvN6q5SofUDxyNF+JSWp8ve50mEpRgedlQ3dKVGjOS
7MBNR2Ki45k7IHOSAaE/9V9dwOiswbxT8VvQ+qUF1q/HbmO7XHjVS30DXX0QEwcFHZnLuttQAViY
8RnIgG+aiqdpcnamwGMGkKs/LuVEC9mXf7mKT0srM311U7AzxmBxdZJRf7F5NAaqCEI1ELhHYpn0
Grc9CGc9R50X6dFdVfY6hTIRVBv/6zteomGNfY26B2FNqz4yWq8VOpDAxG5u6GC/6djN6GhD6OVB
ZCKlG0K379r4ubZUGdZ5zxwXDT/3LcKrrzvBfRg/xuDrEH7ee++rt8M+fU+Fzm7PZEaHEttF3lfl
YzADLwY2Yp1oiJxE7p9xGr298FnvYogpEkRpgXGNmcvNSoGFKaTuT8XtUW1o4TURccZm1ymD1k0C
tXRR+y7XmC14OTVZFnJxpNBAzopa25Mj1Gg0WpkRSgjMs0ybD7nsNONjj/FpGCwkPdiFDqFKCKxA
4KAhOJRAql/8McXpiv1RLtBjIqBDPkkgfPFDkazlU6DUFK8rdJW59n+g9NWyajtPQGdeBRv/5I47
uhcRGbRqHI3RU70WeFdXpXLz4rKICJ8I7DJ1tQxeqrGTvbJrMGwVti4rKIbuxreHHG+FQ4GHLf30
2hHWTXjjdXuw5aNiHtbcK3VoCOxrl4wpAPLTmb7tmDUIF7EyoA/3lBLrH9ir5V0k3VRoyf2UVMP/
P8PNSx41r3Gu0LTKrBaqQx7eKDt2TL6ShDIWSKUP70IG4D8FUCfSCg8cx34efg30ROC2KNdb4iSQ
NNbhpbAoK7UaeiMylDEZ4zBOTNPK9eTIyklsB3PBOuVKPFVPIeKgiEE3BEWpOiCjZKvRr440KTH/
gn2u+PhFT5pE6AZbyvO9t7GI/SaiQbeTfnKAA22PKOXLSsVeegPtV+qC989ojiy0RR+dDYuVWrvK
6dArd/OrHknNICGsRgXPMdL0NSH9gcHQFf8F1cfbkGT9Vj+5GC2fiPFPG9POVUSTlZH4DHbiq+P2
sTKUHiLUij8w9nc9PYZDoE6Gs4OaC7lMVEXAebkqrtU0kXKRif/yRf4zbhTnlgnOdQ/ZDTjWLuCQ
4agbpSyVWxLn/dIm/qEIs+EBrte40nAWmH7fZgNi+pOsWhhRDZzLEq307f3KbWWTeD37FyKvK2VD
xC4koh2Eyw6DPVqtOgywpYrxnsdIb4XYgsSOjCi6r4RWC8HDRuaBfBsIIP/dhnX7vzsqdd2tqGFY
Yj1C6c2aO374xWc0LiKVM0x/4qWsw9eg0OPDWDW49zhYRBBuMu1JSzQtahD84dQstAYYbenl+7Eq
lvg0hPnyJh6gVwJcvu7ElGwYOwQWR7NEqbI2JP0yAZ6FIp7sylZ8XVJO7VPF8ZsuVz1C2EvbOK9j
w2ZyT+TIpnv27mFEYmOEEM30v1rYuBwq0Rgr/d3UKkV/2FNnovIkQ3Icj6ymptbItYdBdWRvohug
ySbNyX56SnFYwxM/2NPP81KrprTOyhNXxPQirpL1pUumxGNe1Xxs3kaUFDsrAxv4RRwQ+IwWIXIu
rT2veaFQoARaTIOoVhQF/Sa7Pj1nc9K6QNGd32EQ5aW8kza9xkcvdxIGnnH0Vjzxz8agP/31i45P
lM1vAlPty7ZbMwjYKTaQVA64XOlwQnF92OTBR0K6cfxac4ItnQd6FpxE06uULUDzbiCDgmkrld9N
h1yBmgy184FtKCqZGX9VczeuLi9xPmAPXIu3GAJ/eDzJyYY1Vc1iaUjxBhGqElPwbWA/1z8XDHZn
1MEwt7wc0nIFgcR8gSKZbLSKK6+m5Jrd+qlpeESWE/zmW57LAxzBEOcAT3eqi4suyCmDi7kiLuNx
iGhMdLqIcbjAN4fVazh9iBsxf2ltCgG24PwWX7+FcsZCtmpDnHXqN3SntiLvRuSBsSgOSRdL92dP
9Vt1V6Dpwk6qB8gkqK0kBYNLzoYgsXPciVGpk+n9nbnvwiV13Hf5ccKYGEN8lr/XsV3o7e6pFY1n
zfq+gUJ9Bb4L8AtmkhtXtOaQguVPIqRfvCANsacgghDZD8pba6CjtOt/mY4CmNOvnYxtqcrwCdnP
GK7Y1CHipuhMQkbiZ7LiK+OZPo/5Yr8WpP9Vh2cneP2fO8ly47DtlgP8zhpgL/csKmW4lFSzfHl7
VpRbnsYtD9TK1DLIMIHBb96ZEzJDGgC4odpkxeTQ2K7fXZryQKY7ApGDT2dOLhOfiLnqwrRfu/EB
HKWJzNQGlNXX1q/VcpVWj4tvhxt1LIwMQ+pcqcqOXOtLwZXEozVTSmXtKc1Co7dJhu5x1BOC3zeI
Xeo4RTCFUsaRT0FogrPrLcNVMpACRK28zMnsdtUbCIyTtV5kLVtRZm4sSZY6sqKGX7Z6u+2WdyZh
PEkhZuQf41TUypDE/xZBdWJFX1XZuA8kRFKbo3Tzs5/2bUIu2vOfQVR9HgqJAUV8g8rsX2Ach6kZ
f+EGRK+TvNYQ8GYz+p5+gagfO4riyy7qjL3zMqhELxtc0WShYa6L3W0h4/ZvwOXh/czG6IWuJLmr
WN7bl6UgwzzVBa+/aEXWar1wLwUV3JU1y31u3kPClknCkHaX4rzkBbuAlkU6WDU+2SFyZNFTkJth
VM9vvlMkuiyMvYYB8VXwvU+XBDfnK57mZrtqaTNP3cLOCUfRNvkprIsSwPR5fPfhDYH5vS1pXy4E
JZLDFU5lM3itdb88LMGYmcDIDWEbUQFzjQYHQFQzoaEIykUgbiGphW4yySKawvOVBpT4OEXy7jP9
opHwjg7HHR04kEPlViHjpaBlt5Cf9ZRrgMWx5qqIVojAmlaIQAmfemHGrW/gS3tFcPMaexiwUWnp
mgazV15jNQ93gEnBCvA09B5vAM1gSx1crQBKcvqXFdN6jj/dNckzOHB/MeG5zaJpNBtOu9H1nTnN
HbVfdYvHyw7ktHSP8KR1sXXnkRob3l9RU0FrE50hy+0g97MsE9d6R6d4d2euSRtfkdPFUf/DGGJd
tmPJoXWG2Pr+BfHuRgrGUra7vqprzgJp3jQA+hYcO86MVER/2VsDU4/MkVPYYuMitGyUvUtRhv7C
wKtAjzVwMzipOdnDtNmZKIH2To6FpZ7W7QHoT8AKVuRR/2rWuBFaZ1ymIaAY+24KAyyeZUrF2qCS
EL1glWAsFOzW7d25CCgzuFNPk6/SsBBRrHR5pqatxwtZbei5krjbzS9qSrIY39l6dBhM620Usbgy
T8U9aAtk+tkTCPDFkJYeorCsL+3nL766PxpJM+Mp1aEBkSNatVGqht0Jq/y0k5XG19O2y2+pqZia
vvkiMht9ZK7kn6zKsWpNHq6oeNMXyf7BOapYBky8rbMgm2itic2mJMIEgcz2ft/wEMp5n7JrxIA7
Oslv2XhbFRH9lmJ1/k2A2rGNt9D9+NSlHyVrXwfj80e49r2U2J1l6TrWyjfMX37l4okHGCfiOLYR
uUpiSCx9RQpKCKw7PL/T0PlthhP711axbz2lijxXz7D8EzwEbw2eT5I9EobyikEfyUFpg/Mg8epd
mG4C3QT250W81smHZjoEKRlFklhz3Or05tmuLSbbxr2cmyPxsz2iP50qfR74bXpDF2NCPi7/zfLt
xEn0N2jiug9Bvn7TGNj85xMXaD58Eji9/aYNBH5LuUIUHo4DZ5RuZKMRTN8rJ1OFEGVxykcN4Iym
/URBpAHM4ZY7zhlsFtFzIVp/0HN2avaWrZDTPkg3Z8CbeutN7BFQWR5TuOuBfRrzVZCYIs4Fiq2m
54zXc9gnOdmIGpxXJxas5vKiz393MnAgDmJ8qR9BleeRyB/7VzZY/Sb/AytPd/rSOKMo+MfpRzto
AvO6WEIQKLffRUmFNTQVoui5Db9dOZMltIQMkaCnZG+y6P5UTZWZH7+1pBw73QIyK6DYgJbp0y+2
dOXc0ZEcYLU73NrohS9zlbOLyeL2cxo2yPn9JlFGFL+BF8cDBsOV+qyI4UNyfpLaSCKL9rBqZrEy
SwSQRtDBMXpmvQud0WFnUyF3weOctO5ExpGV1UXhcADEFwxBPKkeXk4XENajd5blqQnFAeA+o7yv
9WWVIsRXxf0u6CyuQ1PIUcdsFHcxF4gN36uM00tkZox6eq+viVCEVq5To1XXjgUFtRkWsvFpc8od
dRzxvIlZgEdS9soCH/Qu8pWKzViqQhU/unIIDSP+waKJP24qo3+4fU10atM8VrMLElFcPHjbpkL9
DqyXPlVkKvHQ3dP4wLZNwhqQ2eV5Ze2PKdALtFdss7Uu/EAM9y7is4rvRTDOKB8Hwzs+xCIiqmdG
5qxXbyWz2dA+wYlf+E1M+Uk6nC3pJB2rPAqFhzu5oc5DPCNwv5E8jsA90269d9q7xbpoQtl9NoKD
EJUCrTYWLv4AUtkzlk4IMHdSxq7sD26YJMVQRC7Bq+rWsMo0sWwQ443YWRSq1YrkAVtyUAESjrfH
Y77viWieulbHj6fkwmPafSlSmVkHXpvEsH1UURdsTdf7B55KhqMeBrAI6I7jWTKQx7dWhyPRPN6J
On+wUcYQnlsZYI7iXEp2rE4NRzkL1XuwaGkfBQhGZV+8NeWe36QdZXr+YoQFhb4k+MY2pCSCH93i
BN5a2uUHgcO6qlHLIBoPcNVAs97EBZISQX6GZcEMqgEEUI35GzNlEtde4K7ohwVFjPhEQ6kkRajM
6UKlFzd/Eme1DkcBRNQTVdAmZRXZlSXN3OXAQ6Bmzie+wmPGnnmgMz0vlVf77qU7SCVcBCLDE1MV
1xrC3MpLlKqmYoMmyqAXI2TevC3KGt/T/9PNGaas/uNHIEILMDcoehy2YsOQN/TlrYNgHXVkYRcs
PBdIl5Zwmaz1K2UTvsTKAzwkz9z0Dk1vOeVFpviI/sxsPTcJs/avhdz3OsaV2K6oHKg8DaQcn8Dx
RpcQFCRrE8/0xeQqU4erIb8xkLFQz+UmjkQ1wCcxfDnhhRG6COCI6kiH344ak6EPOjGQRt6//tr9
77FTlr+rPmWR875mRJS/fBJpeBPeMM4OIAiD83ESunCXrD+ebZTLN8zwz6T8ibVwdmthav+TgOMF
iiFHEdrsZI5NGRq43E84oG0abzuSb2iHBjDz2pmLPIOB7ftGL+/rsyaDtHTvdWlLfAJJ5jpI8E/y
Oj5WVWVoPlmR+AzVfSvIkkSWX64S6YQJvn0b0vdRUpWg5NAdQIbR96g2P9MTX2VnVmJGweXvXpnE
IDRON+SyKqgpPm22+BxuhJAuRj7/yBBiLb3y3NKAQu4hKpaEYC13S9wi4VqF9iVvwkiszC33G0X5
mZzN/C6yZrKxditPoQSCg4O4kGTkN1RV/aZAwLxpzUMvsQacJaZH2flVhVtIR7ZTRkxsgIPAOKtA
Mirw/lb6uJXLAGGF+3HHy8ck5+xbwysr92KPCKtubJ81ilq9BRlAm8mAvsHX82eX3M9nBrnINK0v
lm4mAl6SaCZEPRc19iNedcWfgDTjZ8DuVI4Q+PcaHKmcT6soedv/c1DEr7MPRk2Q6NDtK2p3Dwvt
GgmGYKg9vKNtgESCCjUIVcMCPoIXxO3BLMt+DCNJtqvEA7W/FIGHqShWJVTlSl0RfNUURaebT0Sb
/lB1FAMHmsmSIjO3yWXnLtIugBvp9on+H+m12zRP0Sr7lS0UWaxlRrkz53hJLt4V56sX3D2ggSrF
k7y1Xp7jygjA8eCQFp9jvaV3clGvaXGk2eoshMUMf2vCRledaoKwNqXAXGddRsKYpMglvSOAP2Es
Q9ejTzdNwJ6VGi4MjLD8lYibpTHjKwI/iRDdAguYeg1vGdTlBDZc2f+t9ETdtOz2wBp+XuWYir7K
0GDDvnKQQ4jckFH+OAbdZbs+MwLTlI5f/rmf0ERJCQrsJDB0QiN4gRORTG3n3jalXTJRDYLSYpHE
3CLz3CymDVRN5EDX+wn65WYMnAgrbUsC9MtLiBTao180Z4l6E8ATsXXEmrnI6RD6RfWe2Gs0+dx6
1BIIqm6xvAN3nDHRkXHMH4BgLSBtgR0CZZc/wX3LRjSNQGWGd3KwopuM6oUOyp+RtOT53YNWQt1j
RT71YUKj1K46i2RdsHHXqzuMFOoeaDDecZ+yyHHe2ajj3dT9n9uVdXKxeWmZUOSLUn5uK12RDBy/
5oaeYn88/UHVHLngWWQ1KdRh86mZd1KY5vFY6rP2ZOmtad4Y80BPEcyD+4tdZFngk+Yx4zrfMA++
cEdYSHxqG4kQX85fUsraNLF2WiOV78He+X536+8tu0mZM6QLyh4QoPGjaAwA+TAgRq/ynCEGNMyn
gek54W8+iP/hC9Tl54Qi/0NjXRXrohvBuO7vkysv4HmN+gmJc81SJjuMex1VbOT7/4f03ShI3iFB
LDa+Mt3pg1OaegA/J4AsmWmvEf8FraEbhRwaqR5WJ8+KZO6Jqwr0GPEwFWo6c9J1vE9TcvFE2YIe
OFbEZf6HhbhWFEp/3qqf+DNufcEMIsR3okrsXYA1b3D8ZVC9uR6lPjPrjhOV3G/So3g1GCilv2Pt
cSBgaWSE+QHw7dNNlRe/2EsxfO0N7AjsXmYYp6a5NC7pEzNMsssSToC+8rHBXZF+i5GS2JAv55Df
1b9bMrEMYJ+C7yFaOr0CnCthC5EQ6wlrX8xo1g6vFkfmmfN2LCTCLPMOe/nnlLOdm6duHnqnaO6J
pfRG2noD4pRF9cgD8b4jzXrc005wo6BUBE1GCO9Cwzpei4SylpouHxzPRl5XYztA65WHXeBliONu
tCNeCAkIBzJ0k5OAuoLdPtmOXN2KIMxAK91G93YdKfqhucU6Ae8hR0kPccf5Y5MO2XOmkhgoE9zD
LGPEYzdEEwG+f51s62vFmeI7QmH19CjxH6ViVMpFMgJ+LZ/XD0drM7CLeNdJV67X7JMjwE+byD5V
5KYQaackRhcHEVfHT39CRxkR1gnD/9w593I5W0uqLNl/GlueLPl90IM5aHHKLxu/vB0EtCiwTqpY
+sQmXvWTLPrshDBNR2V7FMfXb9a4clcPsoimwAxht1VL0I6QokLcTzBTo5hQxFZZBuMLmUXtDLB0
u/sHAltR+/Yv8nsR9f16m224LeJ1liczb7l4x8G5KShWj7oHBwIUPCW5pxczTPvCZ5UaEj09ElBG
V2ekBr48nmFC5WCd/eEaJOrxpZWDKHSmr+8jUDm5ocow+GiKncSGh5Io4R3Ca+ca5MeegjqSVksV
YX2Aph4njSTb2ClWPxJburKz1DfBdRVLvd6FPqXizwGSnhN+n6QmQ66dziTab8zK4t9XhnZiTzix
q8qRqoQh/4BbroXVeuz1JbjKdTgGAY8BjnpDCqOeb6q/AAW2CBHLtycDPtA7mB9zWVMdPjAoHuFO
OwDftVZQH+IVst9j9a3opg8f9nHXO34BMyEETnX87Gc8RdgbgNMa583xWDs5xN20liw5GvPi1fza
POoyaW7+tWf/3QDUQvBSItYUOzvroidGPb8ef/ElxuNu3y8pRyrdvdKzWrDkBU/Biah6otdElwis
EawC9+nslytJX6TJa4I0hUVpw2MhB0PxXVi9Nejw1vfa0xe0oM6MbHnD9kd60XRvghrW2JZrPCSi
ODbDTPSArZ4B3v2xZCQeYhXd8MlO6XZAqa9Tcp9nku8jbn+tk1Bq6MndsBVteOSrmsknRMb67vYy
UIfKePJxz4Abh+hG2Q8vyGdgpoiLDnhXgvYyE5KNj+FN2SfSzMLhKIk5rP8Za3ImpxvwVF2yVHmO
ayccxmIltHnorOU5EAZLFK+oOPb4Fap3hvieVHDzud8L4PzJZ/53srh+cT3risjXCnQSnuVgfKCu
tvKEpPN0/Or42/hYvDApSy7YqHRH3uN247LatVXVJh93/exBHE/Qj+foJKGR4rgX1yxDfFsNBBRU
qZ7AMJR3nOx297bRuevwDijwfMrLuZgcjPb0330kLR4AmgkF9Jgs+ACCbD0euYrRLrXsrkLWf5Eb
KCELM0KKqRw8Ei6ogumD1YOlO7U/j+9j/9d+ZHxIyd87WGBWUXTjuCJN0xzah8ci4tryXPI2njDn
Grs3Qp+Y/8d1ReBdDLv8pCfKD/LtZoWPhLe69PURZ/Gbbe4/tf23O4d7V5uXj4/tyCLq5EN5grpE
V1nihxjW1pAl+s2WoOBddRBKfh24SV4YLjIXzUdfIr8ImbD9XiOJjGXgvt6/B6bDlMs/JcctgSb/
sfVjP0ossbk2pDBy5U60ve2bv6uiNDGJPniKN/kTaA8MKwfiRmzySZYGgpYxq9j0bW2HQLLE1Lau
Z5qTvYrSFYxiH74X5xaF+Y4JNgNVVE3Xlvm3FCTiSyKDJlSTD6wrCZj01+MU8ghoYFv55ueMOOPx
D/sNQQfqYSDsSFp81oEN3kZ7lwDcvt7PyhqGlow4/49gXmkhAJsZJdI9F58mMr4yrqo3StyOFHYy
AKA0FCAhm8cZuR41wh6uudLjBjbOsbF4WwNDvy27V59QIlZKcfsKCL/pGuG0C/jmQ9SDCAtL/xN+
Yj+k5xXUXLoXvRd8eEpeC9RDogUpO0kaHLxqnCkLagVUHVWSEccTUj9LUdabmT/KVJxEILh8r48I
e+KS6TxFbWMk5X08lxjF+r9Qn1G86pPqdaffl04wgAl7pTBEtIrH7qJA9cHc5TkPrcBdK9Zid0jj
g/AtTFxIYQhWV/T4Ea48QTINauwwa4p06UnacQkAgObm8zCkWFvsfG7NtHLlr8EtnzxiY+lG/ITZ
QEAcHNDH/34KhG0X8h+tYKRjsJnYrd6X+/dy8ktIF4NKwkwCrq7kPTbZfQZwBcJyiVNZdtYbh9j9
7ZmzjbGTGZvxJSj7XM1JyLEtHg0jTi5HwTYMBOt7ZOlsM9Ujirh7kIcYaJ/uVNS3Fjw0e5+mCPGm
YLE9+MFHpyXe2cu0etmjtn+EBh4hOlECNiOSbAlV49i0ipI3SA3FZqz1hanviU691eAizA/2h71T
iTC7dxNqFTNO+LIMvvzGgENOmk9F0/8JRH+1zvhSKhU0hxC2F0rLqAhlUklPJm1m97FRZ31eFyWY
dwraf7MQ+SVPF291mQPq+KbECgk8txOLSuvy+3Hz3l5s/+muTlsCjwezoZH37xd1rQZ+C6wK2kc5
Huz6o1lld6EmGnWmGZqT3ebTmzkTVgdfTh+KpTPkq84tJZCpDKresR0ArpcHJ/RErIejAzBkzh2k
s693d22R2u72o0pwO5wiOc6HcPWhUzYdRmyiCosHVwuqr4YMrPCCfmZPj7pMdRJM/3d54R8AJh+T
TYIgxikjTj3pDkikZmuab7dox5gOsEnZ2521s5Jt2dwVrkYB+EppzJlasmKSAyw3oppI39O/ITxy
N56cFs7dqzM7JB4yueNf90ReFpcN94r2ipY9jb0JTp7BpywEVCG4cQXyu1MjEmKcDV4UNeEOrgP3
qh6/tBGdH6vQsGi1szEOv0uoCGPHYHqZvjZUkZYSDvx83Clm8Ih4mz63yx31UgRpv9zuUO/Vr0Ax
sZw9PisC71CcbKdmCnsHxafPZZneqc28dU2v/kt+ltfut/NAQUvS+eHnquQF1AxJyCqo++Mcls13
t3XZI1IL56itdEVzdITgAjSGbt3HCTyLtMgt8HC+FQ4pw0CQS36ZIgHO87DasCPh37Dy+OyhCdqG
7hkwG/d4TJcs5nJW6VYzyQfiOWqSKPRWVVXRx3UgBFT0l8wzrYdiqULCMmyTVEUYgJ3xyWmhOdNs
d44THQI8q53aBmVkhgT3DkuHKia9HZgmmxXLSnkOr0qCyCxEY9axW7Z7B//FKLgBXH227OZmm1j7
JmpxC2YAGA7rLasp6yF4rTmmKjzrZYqgMLxYhGnMt9ohMWekJnnGt9bB0SuNWAP5niqwYtwW/EzL
JTu/gGoinqnLYqP57HFFMv58/Hg+ktUaG7iha6tuv0eXb1qId6pjZNtGeLtEW3fmr5prUCFdi7uz
27NrqNyFQMAtayw0jGvFpXiZvP1q0L5x6Sugs5KiTZQFspOOQQzSxjM6UMc79CSVgbcBOnSw/DvY
Mii1GccGM2fN1M9L53ypQjadHMDjZHDJ1XARKYk6kd0vKNvg6ry2SZZsCTTwAMBKsHGxPsaWGU/N
dgWDzrB9OthBu5VW159ryqiElv0PfyhPLSNRQG/ljX7E0pxcAZaO7WRlwIPKbwY+DLiifWrz0Xfk
0JKXaJeb/Ms0S81sI/DE+SftZFHTsQ8Y9ujGfj2/qxv8z42PqAFYiYmZvpbI69+RT5t4s94t8RWB
7WhSZDJGPjaOuFi/Z6sk4MFKlV2o5/nVuCCAULxEMrrhf9JjLUfm0FXOmX329Yvl2fsBJamUE6os
BpOIA6Cqvv/zszIWbpTS4QTPF6vTW0SMEbPXXBwmyuU3JN/3nmG0+E4CoA/kqTFdztMeSBfcHDSZ
8hCrknEqZy/RKsKQ5gZzPq+C2AZZHggG1zeSVflS8onUWLZlAj3fH15gDXmkF1UO49yMyK1rvU6E
zMzEzdmwShLCc46YytJbDzHv+Lvonxni5m9dVd2FwEk/4OVS0BwtToi62AiSS6t2zdT+dRKovHjO
Lb/P/rcaZzKSeRF3nukTxE27m243ThdZNl87zrm7avfDhExF0l8eWX8+DrzWgoDHsZCBbNGKSZbw
9/+IpIbnUoCq/SgXqKBUWO/XjIEO2pNW0WaH+jANndar9bQIkIDhuf76B+0PQjrLl6vdJUWXuufG
w1+tvn4d9U4V6NAi89JeZhu6XKORMEZHK1DX1is1qomOLukwKRRDaYZjUfo6pu0LIdCIxEvmkP/P
++7BxXOq0QmrmCe2yh4/j24EMxsQULTYtGH0TyrXj9rSYlhee/LapVelHS6ZWq1ZdK5kspmzr7iJ
KU9qfkMrE25ranEnInx9AAse+p3ZSUjP8P9v+f2Ae1g9F5Jb7H1Kr9ayo0RmUe2kS2x1eqoYKaLI
ebbjgPd4Ps2h0X83Bp7CQcuTEDIREcdHOSraBqyRsIHj7wPrBfOxyvm4WbV6Wf+hmYp6yqp+fg60
I91XY7lYdONjg+6X3Mtbb9tp9h8GdphQ/ntd3sNDFQdyZ9Q0AfdRVEJtZktin/1rT2d0BFrWkmah
M8fG4Hqs/swOycCoP3M6LB+W0u11jV/mHvDurgD2zfGvtc8QhCTTeC+epR6wFInEi9DuwJehupQN
yBuYRqSZB8d71Jhv9ELrxV/KmeTc8bFtEnDNBYKLjYg6dJ+hOAezAKZqVclLetG/WeZTys7IaTST
djjSy9aylfC1yLWkqNClQiVQBT0q9J/TrkqBz8Uggb1lFPoecrzlIs+yY449yTr0hPKb+kHqkM7R
TGx9dlNJzKuT7Ylx0ARcek46qiUW8x7TZnf4ei7m5WFlFGoa4YbkA0JuqdLRFsgaxMZuOnOPrfDT
NusuRG0zF6I9twlVrLgA4R65LQRgRUPkCMxKRRiEoTrs0sAiYW7HMnHFdSNdqZJEYzTBHSSI+ptr
N0ropplfOw4h+PtYhr25ZlIC3kbsgDtv2YydLekwM8/uCJwAiJp7duF+ek5o5YYbqVtl7rmB7f8b
oRC7rCLnh9tqjgRidt8YSol2/5e2n4OXxmoBCOcFvX3lo2Ideju6qlCDdGHvpEe9AjRgLPAGdJbp
0ui1hfT4xRArrGo+MhxF6O3HH8dNT20V0zSfzBHz9C+sQ1uzTV4gCio+fJipGbEBVh9bkSE4uQqd
0t8tuITk5G5Jq/ujFcOV9S/MerKvfMKgnePvkQZaxjCuPuKEw7iRNy9tSXcvPe8crK0PXsfpHUaS
sLyKZYDVtW/NUaLuDhoh9YGr7nrYOyx4LtxVcg+foZBlXr7cJtFSTh9SMcIgyFger+MMhGNgivOV
cah0Tr/IZ61TuPzUdzG0UunjojTgfpmWMB74Olw97A77ACw1JVxF1HxGQDWUpk/8lyC3js40AT5E
1OAsjsfCkKoz6pc68y2K2WoBAOJ/3aWNwHedA6DSf3jWoEXSXUkjkup+GQaV3nJYJMTFZ5sjCMSV
2sFKgX3S+Tkl9YYivxbGil30fgKkmaHbFGNKDJs5UVdR3NygItuo2PwwcTBYKidERq5qqmWATMaq
8F7lyANOGdsDx4VjDfVRAMjsv02wvtEUjgSqtCrE6KJBAnEvEmEM7ulBICuOZvvNp7AmohxRylWZ
x4Tm+LhfWRo887+siFCvvPBGHVJZ862rG9pDk2StkoHXGOCLHVMoYk7U2ZFAoeGvAlxwGAfdRogo
0FvVwYIwSk2yqBuhs2NxSz41KBtkxP0XX6/frWKz1llCCI4omODcmh42CQTYsKh1v80JZwCsIQWa
HSdIfXcZaN7DQZGtWr5u8kjvWIibKbgdFbB1AzhWw09SPWbJMs4lcefdB8pAqqk3nUdBk6jmzm4+
OP2XmK3TxQzr+wk1qAOOhxIkYFHv0DyQdFoUdNJQUHG/Af+QEgiX1+qL20/dj6K1KwDI+e4/8Cp8
Dnev+5YqAr+2mgoD9ODLurz02yI/zC8qgNwJxGyDPc2F2w/7UcVFEyL8QmxnHQ8ofIiEkQL9e5wd
hCkvoVFq6qFoAhX6iTthhlJIMDpCSqUzDoPKycMbUOKtYoYxMRVeCaxlB4hbWd9JoevPX9SFq/2r
R5dEOPMmEiLYzmYVteubWK6bgJaDm0XYRtlqh7Ig+O4kuG0pzRk8O3ey1D3zPyyXYyVaMe+sD6Ji
UgSQvfCkRCIVzy021DdLo96qnosx0tn/wMcjjjjCAM7U+9N72dySs7F3mvSfMcP/depjTR0xmYxS
BizGIz0C9swEWkqhqZA50ACPOy1KIN4RATLFOSln70n6dboA9fFKavAMpnwYrdLr1+4SB5Whoo3p
yMUVNOR3kV1nL5aoEH0ImYDQlXETzbJIYStIBQGcAKRq//HLyhbiqTfhilNjXJvWeRkqpuO+1eYK
sOuL4QaxSR2j0D6jcUe2sSm+kwJPFT/EAV/Ix2wA19f9EbRfWafvheBM4O91sBO5F5xSYwomxcOr
2M1VxJDCyOHBBRJvMjOTMKWKg97z9bBXg//B0yzPCzqSqQny4fKYBTRKe8d5mgaXrSd7h/r6JtgY
lCEtqgFgpAn2ryCZZHmTphuXCeSvV/G5/ltBho6rjjZAIYm2cpaeZtWQ2P6NcCSpRq1e+qyPIdqW
GL4FjdxoavFhdFxJPOGSzKkYu8cEKxeCkPVe+SdVbMXtxGLWE4syVQATzZFJHfXapkoR7cAtJno+
D5qlx7tJHiaaOic8XNcGMBPz8Ud8WKQySKHrmwdy2KyM9zuCuO6A3IIAAvPARz5clxs/A3OKUqPU
/H9tk9N3tLStRBxghVdDcaEVoaVeBBIcjjT6Z0s8yxSQUdgb+rb/yIKNRQCQzoI9H9/Fz41UlNLg
DEpo0KhakwmNYIkyRu7s1XIwIBfSqH4g6XxtxeZyEw5L6luv7Uj4Hm5SfRrcy2y7eeF5Yg3+0kFM
JhVbiUR3tdQDBqhRlgFe59Z9QgbxkiotH/O7msDCn6K+iAcflpXveIvpTp6n8etMP7Lxj6QfOQER
7Ukxew5bH+CehR6nUCyMFi+0Dq3FsnYQmHj4xUZJdJaaZ3nOAf/5wY6Yw3+EnLkLARtv+YMedUqL
71fRWgc+GK7AEeXihb1zTKcz3YPotkcOLA3bhdHGGWkcft3U0S7u++g9wNYqr9CHJHpxSCE0r5Ca
cyD1OtiCuAt/4BSyN3pxVXtzNGy14tmQhMsLXWE4VLmXryUCTKOluOdjUys18tkdhRxnPT2F2OI0
TPEsRzdbur5oCJKdR9Zb6W69GnlQql6laSyeGUFD6gX3k+zsahto/JJzfqROkAoeByNslT1QcD8q
TZ+3chN2M8Xu5fmdXpObHtB7+k4FLg9OSvoHmvUszbQ13Gu0CKf95E3hJxb2KyQpndFiRHXevQzZ
h0BR/M2/pQJscvkFku7GlBR36CQL6JBuzrzS5ON4WZPOpbRyFDlVsvWWbgTSG+X2kvatlEjeOzeO
RgMrK8JN7/+PkchmxScuPf5R40g+fZpJv+IoMbH8mEdpmu+KSHwlX2DK9TcKusC8b7KmskFzmcRR
oUaxyzVsQ9r2C5oc+03R8PqkohXflaNyZrT2PsvmQSrhWk3GsFTeGu/CI+xj1lcjVvBvU89bbSZF
jkA+bUc5pxD44laRmxAcpXQjkfs6MgeDblvuBwzSM+s8St2AKpl80Z32eEokoeLuvro08wIwVwPy
UfHispDji/42Z0vpWShvtUN24dzYkL1Jhjqwp4rFsJUDSPFo4wJN7EtTgIFFFt8/VoW61nFQ5Skn
fGABCSuZy7aVGOgwVTwPUoMrU94tNTyXSMcYBNJWnm/WEB185CRKOTbzCVwCzpKBDSWEGUVcdqKI
SfBNcq3T9d8gqGPryx4LtpRilofzE+QZcb6NvhwCL79OH0r+Ppul3K3G63JFUWNmkEroM6dN0gXP
J0fSSygodYxeLZ8cN9sGjlnyUxa/P3jQzY2FJCikk9zCd2Uy3YsJMZRncEyeN3rL6cEdiMb/Jp4i
mBMP2c5fZzu1N9XUFqUksqoBrgFTfxvw+fVGAl9lr40C7ymtOyQQP7A6UM/lIIpQyjakO56fBKaO
a/cVwMObNSf/WmEFC012+z3meaJIoPFnbnM7p70C196gqhc4h46RiE3el168i+Oi9f8PEmEqz8JM
Z7yyjm03k45e32j5mF1Wxp6Yj/2fnwRcDaDnLpb+6kILRiSgx3Sbg2avs8sESuw+JMlxg6L8kpoc
OSOr/vjXWJBdzuERJzySO3+nUM5K/HYVEYAAtr9HKFqSj8kxiGyCax3yVksdQbq+2A6DtRNE8Ksd
y/fiHO/edy6SsAG8EgLuz7CF6FLpGDR9XqFpKLfYw2q1Jgbi4LqerCG2Uh8W+hr3u5St1aizNYfV
/HDpYmFSN79JaX+oiUL/WugzfrK4SQ9oftU806MU/M3hpepUfrzjFqP1kU9lUMSv5IkwqB3z8XCV
tnqGjnePxlTHrdCvhY6wyxqowTYc6q9F6eoLLDw/I71ZESW8YmvvWsA0D9Yyfha5uLRhRWCUd45w
TAr7YIf+Svprw7/5G7a2BCaUttRXohyDN7bKJAStekK/YMCKjII8pUEJ3JvHVawkKB+rTbZMGmxn
F+bmPwI/wSKo/+x9CLKwEjX0pC8oqHB5iRKQrjBEewwDF8UaiDxBgbYUESwtlHCTs4aYi1nI9A5v
KbRtAkshKl3ujPc01PqPmESgRDGKkJDqcQCllePrzb14B2laRTMiuIWnn/YGS9x5Ae4EbCBtWKlf
UCwm9FQJ1OCtVkItqY1eajrXFSmLpMjR7H33WgR5Ai6GAXgRgFalMRpz0qQ6c643FjJmXco281wd
kMR9xJx+dvaKqNRBG/HHosEDfY+EX3xSKRTx0umGOJEfgqob1yBCrZJbNsKYDrMkuLu0UTgK7ZGY
mCnG7/DFNRW1Q/5VgcniqyF9M7h1kF7xaJ1qfCGbE4zRbfHYtGjoujmB2zmPTM+RTXNjlYHju5Cn
GPm2T1MX48grZq2MdI0XuWRdX/qbcJjF7RiTWHrocEp5dDUuv4iZr62f7y4d9VukHfAsypLTTE8l
DKMqzMp9V6PYf0Mn6NTQaDlEdqhXjkVVBRhwlsWVshJweYd6sLODHdzcYmbxIabbGOwjsBPm35rl
kNvhKq6XPBf5KjT8VwxwXTSi4S7/Kem5cL0S+7xXvH5rjf0k4dzq4juxYqRnKS4mYTZVSF2+zKWC
e3xDVCfJce6GluCSqJL7rvwbTs9T/2f+UXITxZ32emOyEiEbZlcnoPeOQcqh35dSVcqHNRjSeeoR
KItB/2XBq8ZkjeuSuAZ8zaS4eZ9nGue4j9Zn2Z7XQ1GLT+6F6XKXAytJZo9L8FZL+YbRnL7wwVcR
PNFMuNH40JvW2Z1kuFGxVTse94c3xe3b8hUeIEHMdwRLMowl5ktexM+0hHEQlvot0BOAAQFTb2+s
pyFPiR+ZAYcRz7vK8pYqjXhaQpJ60qpB1ckMhlpesQpi+O5nfwciq0OUzfOaJoqI27xONePwYnwO
fg/AnMmmoGZwSVjEn5cBeen6CwlmYV0Ggoj3LEiJHZMGqq2ptGlodcljFyJbjpfOn/jtdFpFJDYU
ClzE5t0KeNtL8H84CfZUSm5Bnhi5czMbfXbQ35QXXl4x2ePuO2prg/owEJZoVLbZ5t4CFj/dCAuS
hvUiCw9tLI0+MU/fx0R0zhBOz/gI3Qi3Tb9xXkc5pG89iYoGCH3gDO8ZF7Dh/o1M8GBWDo7KNNba
GIaRTNz4YB3gAqXXcQvq0TGr5zfBjlPGQ/puDf1d1ZRUnCbqOOAeMzjLui4lCeJ52+sLy/b8fRdZ
2sR6LARo8ghleh1f9wr44RZPhhgopJ0QRnWDSa/4qwd9Ax86v+vOYBSxglXlErbObtSKXuqsbs6p
9XyTrsqup1dzDBHP4z+AOznmn7UjaWrvhd+JeYG1STI8pmRai3Fv3Frze60oMbPyJX6U17lwQ2JI
TO+A0EiRojW38lkdHDXVUm6RoRI03HR1sJ7sDdUuLcVXaZcxLSBgEZwjpn7S+DIw1JYfrtFkusnQ
o+ZVzP1bLgvnUwhNMO5uZuK/m+d7J1LFh8x8z0+r6XU6a6neU1GsHkXnjhQCfYUmOIvHtgXfrkQr
YFLYLM/U+w6AbIdtRlKsyPulG/fF+n4HbTBl1XvaaOyY7S6OaWOwM3baMdWZkDprWzE+Bn9UZdRX
jHkMltpzl4NfwjjePlLVqr974nLYYa9oXzEh6iDzrggAjv7uss7NkefUsxuwmwosZzHT4dt8XXeo
Cg2loc7fOIs/bYSsSo10bkbw0n+XPCjE4Fbx4jSkB5WtzhARAwj/wyeCVzRftIW7491P/gjMNpIM
8TFliNPplWSvwxkzJDyn1qjN4E84zSJtwSNCn7JgW4+YZZ50jl3CuaBOksSn4O2HbH39zU9bl1mC
vl9TbwvpgIALXzN6eTswhKvRiGURo4n15ix9h3bG8WdsWnGnqdZXy731uxH/BeC5lT/xWeG9Cepm
8GvTE29dppqQTtUSvq5SoO9HY34WF94fMKobhRTsK5J91QYYidBA3bDgp3bV2qX+0RCBEfS4v4uk
a0ZoGSJod6teaF4edcZqh36XSnpLzmOJPZXc7YNQxz6rj1P/K643T7+fW8B8IC48ODT+jhTp+8HN
WRd/5s76XuzkqsfhvfMim3KXnU5+L0r1mgbuIbyTRCQ7A1mZNkWRR1bMrS3heLqsSjGeG08DQVRQ
p0ZiojuhUIlE54vNTv/jRpHDXhZmH8XU9HDvLm7UVDADtT2xijY08Mr+ht8JtadbzVt9juie4sMq
oRaHcWkndx8BVvn557eX9EvsdylxSGH8/YiTQsJTErmcqlQjNm23V2zy+E7USrSPzs7r3p/xQsZj
iHWb/VMp6y2fGy8VauLvx44WZwkscxH0B5IhNTFNvFuZPkCBUWki12+WdzIjLVeK2UNODFmywnIi
sqcoBCk3kdqENtmpnIzQgvFO41AnCOolQa5QnFZitcWNwuKdto8FtiKwHbVYgSa5//fVEcvIRKzm
vcM4RTaqMst612O/x3MGqYpD842Aj1K6NVJLJ9wROd80oW3MBbuBW6LtcIy0IhbkfZzGg1Tc8oBx
AApaH9tEIj6SizsxN0u8O0EsgYKLVR9TX8rPx9Cl+3oQ2wUM0Wh0XBWrK8IaX+3WrHPq9fj80MaS
AjCvqyFIxb4Qv/KK2XFGfbD55h8yeua+tZP5eI5oYEqHOpJsjKnFgjuFLyobtSnqn9YU7cR0oY+p
t+evwnliypG8uXDvplJOUFFZq7Vp+guTqG60Ds4LAMtznoW/UWAFP18/+Wpn+HGR8bt9LQHTUT6R
jn0qlndSxdskwgK9SEDzy6m4BtbztHn2qFdZRzn+ugX/Ae95i48cWoM6lJU/DNuTwpLrmY3bjfLA
C0WXrlI0NcrEF3D8XAzBH3CiORwepQkQzXsXdTOWR37pePpxvaip73BYK16AX27ujF9dAXEklHtN
TmsgsJw8a5E3lnGY/dgR2daWEO2ktq1gkcW6ZTDSRl7fcvttVsuMTKS5mGkDNFYUYwAPQFOXYhZ6
bruG/vh/5J4fOXjCKMsXQbvvvDFN8HyZ2zo/trsh9VVmB29iPWbqxXnqGIx716tWkIATLVd9z2hP
7+QeYshX+idGL9CnTS1+tBmRqzRZFxplzN4Wbs7pcXn8U9VT/jRFwv5eNXY6QGo+IMk/0AWSLTSh
2XhBvuHq1xDTCR/Zh+Wjbjq6dTPXURucsWTsNaM7aVOT+ib5nnL1R2Jw+l9h8DJ23fYVRMS3LvLH
Ax45z8mDZb0K9DPg2OANCHCGHv1bxADYzEDP9dUB7/dN3pWy0ZkAxdLn145ISqtEOQr459xAN/vy
pq7w+QbFhqWeMByyNkXJ9atNlLCDjaXaawnAeB7UY+kDqc+jgHrNFMIF/PWBZce16cSun2YQk7Ah
fxMQz0XFK5R7X3eB3ILDE6YZQ6rhHOmlpcushBhaFzjmLm9YLzw+zu7cR2Hdu/OLTTUrZMi25+rx
5lCWfmLCs7NVoO3D7kVDedvG4TxGO0xBz+2MI0M9BGS1NWaAOoRxTR3PfEhtpogOx/irGoWIDvEH
v2fe1MmY+DSHifKyWdGVTwILkc62e17s9kUcq+h25W9bPAfIN4PeIDOwXGXtvHYvo2iHKRHylP4i
XByAJdX15PBZwuk71hmXfLQu1pzngv5OJ+O1vimT3Rw2zFhE/DK0ZtAlLVfenELhEQ75YA0vAGmP
zKcXegTwfkL9/BvbYe+pnfED+x18ZNotbb1qm1Qf8jBQySpVwxo2qkN55ci0xjf88KF5N4yhWIUc
iNp+Lx3AXoTNFhHzO8gBo85Py0M8e/AoGjnRaouviT0Hj9AxXpgXTUfdV3piIWKNW89p8AVMFaok
y+ZVYeB61P1/untXBV0h78oy2BTryM2z0KH08mJQc4y84/82Sf1t/FpLxM+uQMI6Yh66aNK59jqx
j09PrWipVO5bt0FC974yjuXUiElvKFU6frDe9mxgGiSrFHU+nfmKLq5RG03oopunfPmlA5On8qi9
ncpFO0xluDPJ+L3olbNMGtwlKv/JJE/crUwISJCBfOHwZbeAbmnXp3UYOXV8KgrYJJu7L3gamRNc
ixsRb5FB19JjFoGkj+flivZXB+KzNftZqakGn3FAU0Sx2qTAcJKsW/x93ZUo1185q05fEu8i+TAy
yrWAbwQ6zf+J9uvwfpBFO3Lbtfi6EjLa7Wic5bw0p1yh4Gtu7g5Qzc5qyx064Kmqjpo55Kcbbrj6
2UYwCGpgT+9eeVUAKPLbwQrb9fSKJNQ7XfEvxgUMVHBoZIK3OQurLiRR8ANYElgjFeJEh51Z9BJc
KD9zF/GkzR0G8VAhSjY/qR/bTTqGb/0FmAoCrxHkjgxYyv4FI1c6vTfUCOl5VvioBnkqGdF7THEH
m9sR1KkiixL+ZlTBkV5V7zlQBfWFRuTMHQEa8WMBVugpi9scoleV7gy25gKsvjHKMW5PI9FCLc/N
/CmiPYk6IZCeteyOu0UnWqHAUZYyLYOnqosCWYOZX+UPl1yWnXEBvat2aj0IlfQWaWfpMF+PD9Cs
L5XOoPD1qlKK7932GkXafPVtqaNtM8cXyBGlSreIYmXG9kRCVJFhBpupT1QxEDoCIOIIxVDmLADK
sahvg+dhggn3sHuhne8KWMGrkKc8UgcvUYGaEpNJihzW3JpYZ1GK/F4ERe3jpm9bdFcyaCImBRF4
0NNQFYJvegfPGFnygtJ9M1TRFh2sSh5s5/ss1jeMZZyLOifLtGtlVC0P/YZXgW22tfuOpE/reBav
X9s518gokjVYB8Wyb7EdYpUDL2Cukk7A05QgnQVfXQGupN/DtnNkfD6tm08653noExI1OV/NoySV
q4QYZHMls2amu67D47crOCA//9SojIy9o8EG9smQy8T4z+iz3GrQI38Z0oOUG6aDdEOAbBSqevbJ
CrkE9NROxjdUISGV+sQgDgmRb4PgLvZSpOUKxUdaCZ7OWn3LtpDeIOprEvtMTsUwHTEO0jHqz/V7
euVR0rxfMV+npQXPFFVTdDcEgpO2Ojsr0O8NZ1JazEgvN2qYFFYODscM2ZvlOR6ZZAT5T97av9UM
iWWzzOdZ84SJHaKQZcur38w2M0AKT4tV3wRR4HbGWtxdJVKLPycnAyArHGp+R4TbWzGhm6K8j/5Y
YHUbS6DR16WOqsstHb0kY66aAUAU57ulGAy2THu9LpWtB6r1mjXlxt7wt46W4l7RdstyOMlyK6At
rxrBO4I9USiPlg0igQi0VOz4TVxazzEmIEa5f2tMA8pH802iq00OtQLYPnW6SvQx9Z2c5a1oGTRC
JodPz6p4Qq5k+7Eo3w2F3+8E2KOCgKFsJjGX6+N1dBkSpGBT4CWDoNe3ZX+S+J0ofescH4xI/W1B
IBBs3TEr1QdWRtbwhYPcM+V03hqNIlUL+KXFWPv26N0Uhsbo98G/3huOcFg1cnuUub92J5VNxmiH
77DWA+SZA7Z6RSg6xkMVSKAtr7j8veWKVxZNt4hizug7KrixM+Dnw8+WFaY5NFKts8y2kA4gxIW0
dlru3PGKtYuwv6wQ1KEP9TvoYm31W5j9XD8KbWHfnr3WlNxEQOV6dcWqci8r+7LyIVLHddJb6ZHp
SG9RwlWmgSi73xTxzcnrz423PWKGEAJ/VPahubMoUB51Z+qal4W46Im+m7N5DH5mhc0NACgPDzPv
+nZwott1FWhGJw5Qic2nIs19CGLlBTOGtJoo5Hx/4/qDE4iGNMbgabFiPNo2IFaPUXbhH3pfN9nV
z2+tiglrn2rZS2xAhYTkQYqwe4lqQFRZsfgwV8Xvd9q5Dlh5qpbi7KXp7/2HQDqRud6JE4x7u4vb
CQ/pRjJd8VGrAk8v+mZkzlSAJRA2l0buyerpRzYy3Of0WZvjsj+2NtAqyYtadtgkKLpFmCrd7E2r
68PDs9KvXCnflvJrQvMfjfVeH7evNowq1mKp0mtL/9mbNOjS8iSW495Ny0EF0H2HsFFXoPJ28s9b
iceaZxGa6pmI7aDSrdcNXc1H41njxjpvCI+sgmk1xdGssYWG8Kdln56hGLiBgaiLsxQZ7O8YQ+tY
51aHKw3xI052cgNsNvrn/svSbNXLngaj3N5UAQyaChUNkLeLDcheKwRizbGqFKi9p9e79YzFcD1W
kT/59byEY7urPLGTw67ZbnJFQdMfPPxLFvBMYIIPByAG62S3d66AQWogkk40/eKV84qXv9YTRkcX
BhH/SgKtckxMI24mWF2a8nIjutBe0mjeEeKpbqiJ9UYSE21vN241wG71Yp75QqZWi8wcTZnsWLbe
hmHbqA3ajF6rLv6/E7w6KwVpMVqgtbs/fVnJkVNKqFFNYfS1+qLcsgo6CDNCbduZDt4pKXzyq2WZ
+42nVlPGgV1y4MrzACMOm9v+h8CAkvWva+zI5ENePvL/dEiotvscjGf/KyB4Nnwi8IvsCTQ+GHOp
EhWON3R3UGr15/KrzYpSY27CcqxOI35FV8pyRw9G2imo2H844IwPhw08MQ2/myrggzEHpXI2Vhjt
osipSxrVbcindBQ48CEwd1mtbE31iHrkHgH53kH+hXsFRPvUXF26GEUVPJ/0l2yHjusfGhCSK7oh
Gp7gvEB8yrBQAGFBPMx/Yyfi97cBZz0qmGm+1Yt36/yNjcD7E6zbylLmG1dVnIw5wqA1vMW5VOjl
BjkEyBERPR+5YCRFH35nPrwaVYu1OAQjGxFaDihxDo2/Q5xU1Z5f1v+rOJi2B01DJ139QOWvbxI/
WLdFppLs71aRiHDo2SQv6hxBzNIcizNQPJPmmzzmr9CEbHAvuqV21s5qDcgOzFu24M/a3T6O5X13
g7lHIcx9jVj+JIWXjyM4cASkazfodagANUHwOjVvRSecdv/pxCrkJM2RIAKfXUlq7ZDdLUrQtffo
8soolDydFyCOLqVq0kojiZBR6Aqtvr+dokIxLJEajtv2brr9UfqpaAGVzXDK8lCYyQr/VvqL5+zL
khMmezf0L+djHYz5HWk7DDIkveV2MjzYzNeGsUlErsYGOkDr4eo7bs+/Qla3soa+HHiBrCFdPQf6
nnO9NsSD29a1WBJp3N3GXxaHpf5ShBAAHctFGEjBFZK883ZZ+KoZi26fcux2Mxz8kft42LLKT7Co
9d9X7/hUHdh03yAP7sbZ1O6rKB6bgPKqBtH/tSziEhy5DnMbhSzTi0m5GxFMJq43/vPy0y+Bitpw
HFKOB0pTM01p+UUSTkwAZiETaNEOaBXuyeuin1Z6B2B9yPzD3IHZuaUubxjapXXfvC1Fvfyzrzdx
9SQxhADTWgoj+tOE9kenbPXcMXJA7yA4dwSH1CjGrXuAtM1RCh6dkU+pfMx6JTcE7/OBgMVdjq8G
tB27kOS0SE3XCrAk6gj7CAHMCn6XI6qMTGLZiOHs+T3+wXtSYkUNXeK6tVnseGbc1DAkOrwfqoE+
Ri8CZnoeZpXbaPbNhXtnwuJaCuYyPMy5twxDVde3HrRZStNWK96wvf8xmxg2YaMjTjAWQ217yVjr
i/HxSuidAJuB2RKdlmOOw5Mkwl7bgEmYz16Ewd5Gsluhc53gEo/48vpbh9sg38GM3ixWk20VX39b
Wx1WyHU7cP/9FXuO+eL5u9SQSf5/+IHm9cneegCIMLtkqwMJ7xX1zQxlS7vOWuWbZrrMdQu13fhJ
tAphC+cGU+W81wWH5zeqUNvMzBUxn36chMf27FFjomOcb5gIZGFmliqj9apK4jv30q64wOQLAUoP
+QeOcCJoDd1K/vT8oC5b5TqSv1DZ9wKTa0jC+cJ0JVw2E1cxtQMAKY+3SQYRP91u7vmpEYml6U2X
GGj5zw7QJqWmcFRs/LgrPerw0NecVuHwltda7bGvME2EagO5BC+pH0fvtuZpo9nIxtnqldoajydb
Bcc/pgVjNJTJKSrKeQpaTYmGOg6likSlKssaLhaObQ/RwVajmD/hcghKp0wHAnL2aezaHSfSTbe0
mYw79YX+D8SDn71xzIrNSHeEy2VX39FjwltqXnH/L8JA3eUkosaPXRP+B3+mAWdpbBNC5R1Tep2Q
RXhQVpkfrmHmtzxSLOMUMsSZC4vqLvGHCgfeyhaUqzlt4az3EBlEQpUElXQNaO7KB7g960cAsWLA
kVUhChTVNVL5MU2HewA1HH7KGup329FVdcOqdCl6XK9aJ/VNVYalf04xlWGL0Muqbc3pcbSA3eji
LOm3IMhWc+7905aWZ2MNql0rFYzeg72hyTlm2byaAvX2MxEA6kYznbP5cVXm2CDLnxFML0L3up2d
nd9Hae4v5zScbOGffRBNow3Dvp5NBp5E+bRcG0R25NwihHDQQFPzjBgcsoR3j0Td82+bOmHV1iCI
s3dFSdhwok6lsEK8/RuwYiqF/csEUvxvNTKcy77TEq3x4pF+Krc1Zg5BcHY7CNixv/u+NzQ00tLC
cuuMAI9R/t9U+ab0DEz32wkB/ky7raip2jvnQYyVVRXJn/fnjt6su1oxcrAAvCnULZxiBz0gmF1p
RTYIEeHrLhS52N57dgVODgG+ktHy+rnR2KZxIF9pomAW34vCA82IYkko9r1UzyqsjAd8ngOdp1h3
+A5Fbbj7wjcmmnKLTCuz6R+HfaQujeBhiwxkbMGBKPEAiKpwXgWK2fUTTB+eksFFSRqfBxXEsooU
V7w96+VK32DUVZphhSAOTLv718KBBS+8VBBy0gEJyz2wqTdSE7wdPr55gUV6DrA60gSnbRL6ch5b
AsqIQg+jsf2Q6vIeBNJuNQ4WPz8yDgQMatwp8vAmT6lMZzdvAMxDPb0A16MOIeI7F2LLFkfKzVCm
+NYTLRshtMMOV9FIKAxj/dFRWsY7kfszhjxURn83mBsuhRB0J8IFLU5H3vrjYxCzEzjbUu9UBG5F
4E/3DAEKygXTouWu6D3MWbKkUCHhng2hboM2siXnU5GTIoM4QOBvqvbTCz8ZtO5UWFU/alYVA1si
N0sPGGixgdsr0QR+khJRf9zmYau4hErPaR/ufwz/w1Ts0ATHA1P3/QgxXU81Q5kOL8tgawxu5roH
+0pjBzwJZaqgyFcd9etM9yrYAKCpdXNk8BNaYxGD96k8obOznq8SrxrJDH2YClX1Q0Q6hT/jX1o4
LyyZmd9rCAd5v2iraeUusUMqSYhT0K+nWBhoK56rBdXSxwLwYulNoZsDuus5LdNLzVRKqxyPVxrX
3sMrtnSHyA4Lw5rxW6756DqncU/AZrkBe3RtlOPTui9aXiYaEIus8tVbM6LYaMzCEmMRevAnZIYt
y6ynmD6SAw52kJzi0yyguSrchLwCgqU4HN8k6pvmM4CUF5rB0pC3lP1BZ0MZ+cuQcd68Vze73hXd
jQ8Huzlq6oEkSZfnW7zSiklAG/wSbMqOv/ZdKMqQFOufgerdSnnKIw0msrK1JycCm1j8TfsQZfCZ
qGN9jL85tx8iT/oYggJz5u6UxkpLZ3TRQ5uQw9SbAIlVm2n4VK+g1ALHhMojnFgy/9Jp7ofeuZ2d
Oi08i5mJn8rOSHo6PSVPOYYbZUpljC1CBDGeWBB/GMCn1jAfmB6pRoT/cPdJYfZS8LR1uUKycVCr
pCToAZwrkp/NrC9bjVC5TsQFru8cWpkI9/0Duk+CRh59KKpcRDHBL3x+EXxrNOQZZJ0FPEswtdXZ
ivs7el0BNNQOZ1U3m21g724UXppKR6cVByR8B21L/gADBvFnZgj1sVWFR6H8c3+lPFn9kg9o2eYo
6fojY3NZIl88a0sMnB3OFlBnyhweY/BIcbuidzasEzNk9WYjY8avGRyMRVP9cnDgAeTx2JwSdqjw
UmWs3Y+Jya+mhyG/9D9CLWnTWXAks7uacahetBNKAUa5c6FCsxmG8v+W346RVm9RF5ZEdatEY025
b1IRRMoaLi6kYwVndKB36upMjVrr0J7Ni/p8WivmGM6qjRiJQpP0/kfqgTCFlV6iLX3M1o6hwBwZ
ezd6pXEau217p+RIEN0lyv9HQbzSkVkcL1YWB0ohbJq1IYOLIT9EHeRqDx+eAw92dI5BVJI2gAE1
9e7gd8cIo86COrB3E+LI0MlA0r0XG6YC6liFjl9VwJfNykpaHluu7C6sztdIrLK/GwWWd3Qqs142
Iw2Kx5uppSt4Uz3iPjmtUj7RuDX+Kxky/JvV60XXge2tAjmP0XZL/BpzBEBlSTDVxhtYUrgCswIt
8l1Tm4yhfIXTAuVVIbjtKTmbHrhchcRq9ie8/wMV6BcjRqBV5JhzbinQGX+0bDcsJatn2m3JxCZb
/g9K6QaeEaXStMXVvAT+QOZv3wEllL6wxx3jgQiF4HtjAOEygcV/cxDgeE7O2g3sQVpGLpxxXnpv
muXnVVyxVJ5dbkbB7jrGLAAYI7O+Jbj2GejOid3KHE+JfaBjcVUwe+JiU9kyRZIlamVSjlwvmqKt
+drz+qf2NaHiwhqcLM+e8rNGCpwVXMwqYeRR1a84TxcYfZwKWR30mJUVHW8fPvUBacF7Lfo7iOXV
Ah4myxsE0Z0UgwYXnXmCxNe5fY5Q3rdiR9Bt4ldlbu3xq/YIkSDF0xwrWM9esXwP6Hovf3yAEasQ
dBSqwvPt6t7yOOJE4/aBzRNPMFdoAVV0msbFTXSPbSzZzYHBPXyRNDKDySlFBa8I8UllVO0QkGC5
hUYtTkyGAZoSamT+8qkNXWrzrf1KBaXpb88KPYgbVcSqe9/lW9ORl500yOdHeu2ttOPQOOhV/TGz
4fnNVxX895qXKuGBN/86OG/ekGeUMuUn5f4jMlUJnYfBQi2b7Cean5am2LtXIEfdbkiJCRZUPWGy
498TJMUrA4qbwFG7UUKfOSSC0TByONU468CNtaak53Wq8Nm3LvuUqW1QXim4zCBwff5EshOOgKDJ
pvuS7YoUDF3+VBy67AB63IADTfwuG9/n9zWPgGgvAxj/lmsy3NA0pQll9V+buV/VQtOrrlbGJDeR
GRZqvXr5oy8sQIJxK0UF1QKyEf8TfRcRzuKvZ1MWv8omHHpeQ/szq4dGniyB4Uy78vgTnOtj/tZz
+KiIhNRRWi159HjdkHfo7cucM2gy5fkHx7ayKAkpTyBelLD1C0YdMgHqM49/cLyI6mwbUqW4YwCT
jVLHFtbDI0XopKECdWO+SKFFkYguAiHtWyK99/BNi+CikKFrsjTaaqQDJiLanncQm81a/5Z+wEyv
uC2w7THVsWpohhq83nQl5eglCOTWl3fqvYMpgb6UE4itP+EYszF+FBpuTNWl9G5uVOa+pGzIQtwK
1v2s5fWfxnoLXVfQ3nLrKcSGHUrBgO6e+QgYO6tRAhsKUrUcGutAU7vhmIu/uJuYS5dRFGazDDQU
mpcFaFVxgZh22r3xAUHUg1RPCNBMR04m9T3bDWStx70+WQenU1/OYEaRYSvM77E7MpZHWqgHnPfa
Fqb7mdeIatH8t9FbwrUKYIE+9r7tb7XTpgzQpLaFPZv47gsvJWvbwJbzOTeRDrjPL8DmGZJIMEYl
5rTvhL42pUw1vf3/23miRC04TSzMV8cCoIhw7cTcMkX4XsNQ7NGnUA9MgIP7j5NBrFdo0L6mTSTQ
gg0cNIu2MJ2O5N4wDyJI0g44NyF3SxSlgZ5v/IZzPn/KH+2gYsclOo0pFIgBiyrgFk5pFHcq9Vuq
DyZAdSixv5VJtJ0QuE2sUlnq18UFeIIjTKagMiY7EoBBi4g4HfhEdnlgjRaK6keaAi4kRYr+dLcx
fgre0M/lmMmZQQsF+82WQidghnaSGsKis1WhaPifpLsxoar9KNyR5AzNn8/+/WgXeJ3K4zV3OUeJ
sLS2Wi45iIzj/Hgg2Te/8VcCd4hc2Vyh+h5l1IeYYv0JLeMliKTHfbdx4+vLiNLsO769Ciobbz7w
XK+/q57OmCd+f4vOW0aFcbZRA39tpXsckKM6Vtir4lC8sC/vv8FsiJKbrR0izsQJH8CdvkFsgcDp
+oN0lyjaahFJwILJsoC0cscmfH287eqmiI0nw1qG8t1hnP25OprXFOn92KgN2OBVx38YfLF6ZTNX
8IzuYo7YyZ1bRKcmKChmPDyMkvLqvhCRvShuWXvwdXLjab80AEAXGy+s+XCbLdBz18lSe1rVGYG9
QJc9GFsKgKKl0IikWbTyczhDOGTJetbEKC2htEwWm3c2Naqp+xNHn4JUj8uFSp7TRz+RGDMJBs6+
+OgQIWjaQvnoaFTakYktvQzMD6xe9S+whtec3mhdIHpgkv+8nbF3A0iWa/3KLnrNo7tC9K3AyYMb
4AmI7iyFF+bX5y5GlX/mqj/0YMoZF0IhnvZU4LayILJ8KVmbiJBmCh3lfDE7h7FJIJaO9G0C++h3
GwigaDVy7ZZ6LV8lDcZeUD5GJaxf1ceFWipNa63IHh2VCMk2EKyZwtQUOkCiqt1IYwgxEC16O1tF
8BGMFCyhoFl56mv/vC6hou/PQAhktXBAa7xRvPPRL1QhKx4/Wb8tMNP85Kk9mK6bGv+GOQmiPBpW
vW1DrZkZlted9tGU7tohj/AMBn3m6hQYv0GqUkM8rgw5tRHem7sNpkzUBtgRMairxy3+0LUinmFI
frHac0KVKKr8OFC1pI6Fjj9Sx67AVjdJ7wVLI4gZ5eTntfWtmjSm3HanR2SoagIRdE9BNQzm3G8G
kEUD7+6Q2auZqeltAghZoNKyUJjV94AK6Gh5tIlmJmResk5IbgwWl2FcEKf8iS4JPEw5L7uqzUSP
WxZ/eq8RNJeBFtTeA/oUSbORFSvUO9wILUKADBqZTF6+mVdRmPyAlzJxZ/uL+BKXlXK7O6b8TY+w
oYEO2XcTZ0G6JyzuzBgpdKRZVQcpSpjjQOSDXhNC2PejKu876GLS6Uq7SXPL/OOZpXb+BcH4OsGK
8B6IcxAVJfKl2D29VTO/QVi+fWCDvBTxglVWH4W0Qc5TdiwnnfqVcoijrLhR6wJXdKtWDqq9YWeL
HQWBfbrOXh/We7uUz28dPs4p/CXCBY6sWLorb1gaQ0peUGALQFuBEmI4zq7b0DP0DPrZT8kMvWy9
5Ykr8xpyTZsi4a3shlBojVI38k6AC7Av0NDHkftZBQL1yM3zJ5bvxU5U3c55iz9HAmzgZSoWAvq3
/b4b5IZXuP16du+tUW5WGs1pgtPpYoUDGqhytAgzCGWaENOKkMyYoH7Tplvz9+JuHodTs0iaqBSz
YjUA4mblobZfzuCxHRNreDfwrIByTGPx9y4mCRi5lLmabs1BuGW7pxHVfPxobKXybHd0wB+ajq5G
1IbfOcpIy70L6HUfe2AU5psX9a/VAyMRhicgqT+XvxyPuzcjWxk4Z2f6AFCjDoduvLCHWqQoo99M
W0k/fpEwjP2hXlnuJgEnz9PzIYUCuMl7sMA/F34Pt8rXbfnX2qh0Uy9XQB9Lr0+VKuGs52pIP3Oi
ARobu7HuWYJ7q7mfYeUq22TnybuE/NuuaCMcKdzyF8D1URehmXuw4x5N0+fjz427c/ATxyfRqSco
vUs0N7A/ytHDMd06Cnc2Yy7B/K4jEABo4DOamGF8g1XrWUV0TvEjYohGt4K2863HFz6ZHJmJ4DMQ
d1C+x+ogeMGQta6LSVpLToYdbQiGUi/U5PYnpa8JKnRsUdchHkOWi8jBHBdJiOFHxIpUOD6CaeRl
zowdF6OSFauVV3JMfdtmnRD1/8PPanJXKa7KdMRxJLHRPoeaDk68Qgqv+CL9fVC0r78V1O14QKvv
+FuTknobsLOyUoYdL/RJxnaB2SrC0BJTJIvuNuJqMivMrAl8wIzloJ5BEaTtRaoDEEALcB1HSGFq
IKpnOjNCZdSdPleV/r5Ipcv5Y173PMcXCahQW4UJWkWZncEkvqbCypcOb/BrPsdTaP6Poybhw9n/
Zx2aPXTIKvmTT7LhK/IZReSX8rfJbuDye0vebrDjlHMGCZM6ZvVfYkFW5G7c0iEd3aNMqQ2JXZNo
0xvx4rgnMqlFJ4F9vv9TIyWGPJRXeuc9PPGgEhju7F/6Hozp0WcWQugCz/2z9gfEdDI9tMRJ+YaH
nF8ZR6lDmaEBZzjWzXgJIuw6B/J1L2B+mMHUAfsMbVTwk6464IxwqAfuvF2mSzs8sLVk5TlQ4MJw
/p87PvK3tY54KLXzrIXVDXgU03Ebwk7tPGHpVUSCEGPODVj8QlyfzgIRgxBJAoJIE9FJv8zChEkD
D3caEEfkhlhEM5k+skmvjP4uK+9G/1M2M7C7hJRm3Msd/GUZ6BAvq4RAodTVLZtbp4TlN4CDttRV
rpDb4aYYCmK5bzhCbcnNy23mLoVUo0sYIM3BKgvC8wV2hkNRaM6PTxdSV+N7LI+BSFW1bRlEbWE3
e1GIIIJbiJbKw4mxtXEVguGDyVoQGp7kKLOqAQmXA+mexTKY4nXUhePCsfFH+CaIQVVt8IBkv9WR
ot6jQO5UCaN71SYBnUKIu34HB/GeJCkNOFV82eUU0BJwlFSyMpaAlpoEN5zKeO0r6BKuQntH+Wu3
yCNkzEXGBrV0oEGsw8+GK9gJ2ydpPxeFxRP1W/sdofJy4sXk36Um9Dgb2USL0N+e2gvaEvQZmc33
MwYk6SFAqU2jBaqgMqIzQP+IubqafDz3FfsdA+xRXvGm9WgvehB86oZrLpx85T4DCHc9b54sKb43
zNOHAE+IQUZK5RhvqzKnfZf8QtuVVIVAnrKDFWPZD0HwNE+yzNMCpjZ1TjaKrPHcP4h04t+iGu2Y
LlPu6PTj9c9EmGhZ4IaNgyHluKMeo8VdLQXoFuiL7bDR1fAseMF1XFfUQs5+yQ+ruUGgLlv29/Jn
dqVY74SPoxQBVyVQb5SBsx8oGxIUkbbhmMDeaku5c5s7OasOdUzoGP9bclSMCHrZVoySSy4k1Cxa
JwkZ8iSPdu5DpRrBDZspZeV/BLGQ4Cw1N0EgTAZxRrSCcFsON3tgXe/D2GJnp8mYMKpawY4T72SD
3bKiyKgFkKYo6TRSSIkriFw6NMYz6U+KdQwdQnNswLCIqr99zCz4YgEiuTAyyEah0K8jqnnsbY3S
iUGVA4UfIih3eT30Gyu6taeLkEFBmARwaBrE+AhRNieRVFgP7VMSPOLpj/kz+rEcdvo3biGbBpFx
1Qpk4s3JqtqYzoL1VUyz8FF4L6B8omK4pplcbcIZY1IrH2GhQo7P6F0hbtap0KK3AkmpfRTUqGnX
TF+mDcaM+SQbeb+PG5xY1ggsjrHKZ4tbTyNh0mqOk5tZCstWmy8sGL1AR7gjQ33bMpRXBu2fuBwT
wvVcTvApA8GDQsiZHDVjN7sfYcChRDKklOXZMiYtB1ohnrmByP6Td6FFW01b76ylHU2D/8VaI+Q8
OBxJf5osRWZSH3V8ajKNYD208d5R3RQaTNOVH3WqxB3RV6Ha0szdFF5gdcOea1W4paUtZpOL4MJ8
xTp9Foel2sJ9ssotZl5zQr280iquoNiqxBINX4VV5jbECYzs4T4v5hoW2tXyQae6QTqnzJhXeOrb
7SVTnB4tKP2k8z4BotLh45Q3xy9echy1XoXB2RgEDg3qF09/wS5HqpjazvUv0+EySfi09gy6wLRf
zU/QD0uvjS2M0bidXYdLLOpsPHouLmo9sA7GnGR7r0MPTu3AZ/zmwkgZvCNXGlOoBEWzIgD2NuGr
Fro5xnixYZr8O1h6IPE0tG8QD+mOxdYJAXNtXXplgbZIj4LxFBE/AYxPNhFlSl+qyr3XPddZXZ/v
zy/mw+TZryAV4lA39priA8arRFy30jrGFM3lu9uVJ983svVsThf36OsjVglEYmFeM0PtZhSF0ih+
h3OWiFxW8r6eDTd9ahmPNdg7ouxKLdOqYj0wltvjODgLyCnyomdiKxR8UEc7H7LI11zFF1UdHGNZ
JKsXsTo/jPJWuVR9VXbrUMQupOXrOuCvY9E5oCPQ+/9HGDY86FqVHpLCcH5Lg6/RkBDDJMfmjkDY
7Q1lZDdWtG5Q/IOKBMe5bwxgBqZE2ePIvtXYkj47Y2cWaRuD0h6ZQA4hyzD9QRKH3G8UjygxD4Za
0uEL4M8IjfhTrOwW1fWNj1d0xOUEoOtH5JHaiMP63ytZuM73ZBhfLt1N+aDFqSmVyy2Je9sAFPfD
ICtlaoAUEaDxN9cq7MXYy431m8baYAElM9k+3+eugY1Wu6P9Bw1gt/Aeeq3cRQPiyxAQEsca4ggs
6bdj9kEIHpbwbd/C4d1xrsSznz9cRucbcoUN/b4WgzG70HmkdnAbm/1FfVHto3zBWsxVhDojLl7b
7T6gXBwUodkuPU1rbS4I7ZsgZZAb8lj+tHC5jlkMf1guC+kMzCti8Du8cNb6ms4I3caDPln3OG3P
X91Dcm0KERnbdxndscCd3gPPmwRiFnNa+otnAiq6xX97TmpXaaZTmQxffWCaX76Hfh9ViUGU6CSK
tzUw03ZKXG36uOAVgSoj1bmEgUayc4UWl2PL5P9y+aDrlV93GFpAwn2QgD8kblOzZavAJcfSUTFW
nbSdmy36Wrwg3ZRSepEgbZioXpsXSTHCbHbs45VuISCqBmRvp53psqZuB5oRvzmluCFxSUJmpmin
Ey02TrHQMAqQrxrzjDQohTaLuuJfm4v8kCE1TsdXmXxzl4reajk5vFTawQR9iDxjpKpyJVt7hpw5
maBxwOgWTeuXEwWRQG2JbwiOFvatz3EGSk+bi7DJEkFalpDG2l0DOanbyqkvaSVf+Lnk8uKOspaq
ADWbbbpMYMjoGauWRpI5eBI05W5eJ8qSD2aAhARB+/TOLWQzbEdOaAoC2YBhd9N6ZZ4yuXIotm8B
BaFU3hoUul5/6rhnfxgajV5SHeNvwlOFGcj31Ooqrt6YJT+Rhm5dR6UUEcp2WxrvMdjN5fzAJgmd
ESKecbSHrVmpohSKB8CS/X/WrYpdzpBSL9foBxS5LIh4Ixmf4AO5ZPwgq16TOJEQGvciumeEertf
L3p7iapktwSzH2JmYcxGhxHJh8kF9qa2SCIQ79liDzRWHkknBn7sNBrtFIj7uUvAXcb0KcFNbsQU
aZ7D5v+TEPsbIGCaBx9beDLMBesM33HsE/Nt2KNLOfYY9Pmd/sHlJiAhkHtneEN0zlR0+gC3kgwD
fnIAPqFuzKon4HKpNKkydEtS+Ohx0J/qjKoBkvMyMlrf6t+1EHGu2yybYiAELmnxp5CGFJXkwPeZ
p3ydre0sZzcVyWAmD2ImqpL7hHz436F7r40k2ZdMuoq85WtfFLO8tTWL1yIN9jNAUa4AuS/os3VI
SpvTXRBFbkWF2QtQiueXuOBwz2VZY4QMY8ydTW6YtDW/oXlAtbSXd5WYWLL514stUU3IUZ3WyDCr
oDQIQISEtHg2Pw1TylvZccViw0jb23OfCBxxxjzfidO7A8Q8vPf3iLOkIJp/CepFdRhl7jN6qAHk
/fc48obC1oi1IgiAeV45l+JSBrtY/l9/HpY1Vkr3m9jn/Uy2Yubgn+RqgeDMaGjJqhpedMvaXqN6
q+x5kRnoKaUt8WlnlY0CVG/zJ9g9oUrsflKXEiB3n+xuDJWmr5fbRRWg3JGKAYd4sA+qf4DUCFd0
JhN/41CEOWRg017LoQlwWYaJjAtw6WZrLJgibI+OedJehe9Lu64Etbi+IUfqC5iN829hnZ1QEXIP
UzQoEdLpUIMSByfIIkbXby3gRK4PU2X6p17Zf3xiLtVPAKBfKyEKXJUNg/XfIR5ytHPLr7Ir7oAp
no63IKwNM49sxQ59VJZYcpbMdo7K+LKvMH70c4Wg1Thj4JAIh7jiifgqIBFh/wJaUdgghEumny+I
3ZAbl6f/niw8IME/txIP9j8zUPIbjSaJTHk00Q5rPH0WmfetIbg3KcYhtfnYTRon5tJyl7I2+ix6
ltDFyYX9aubfP8VuIervtm90ko1qRDCi3xmtFvFxaSAYf7QfOKt1tLftT/cBV/DIC/b4TtFTdlhw
DwvIQ60o7xmSFq0awyXXR6lK/qVB8h3vIwMbJMxaWZ9SmAUOaSm873j66fvCgk/cLJVAgekMb2GR
k0b5g4SkNdDKJn6cjEvCqd9XARGR6L/wfOcfaNY7ltrueC+BegebhRjbPITHQzavY2/JtCZqv5+S
Ogzfnfswey0B+GPMKjxaHsq85CWAHRBCwQfyIMgswII3EK7AmAuGz09ShVX4IvLl0bbXcKi1/n/M
Hwivr88h41R4EnIk2iwMRAogt5vfIX6HqHerS2AtbPeV7r+TepYr++pyW7MfpE3Ii1ki4HygHtBG
jg8b6NaRRPqUVn4QDMB7o6iI7qVRSawX3awsLMEIQMe5EoLF42DQ1XOjkTPxyOEulKY4i+bNt//t
xigDGDUffwgR4YQM/xU4msQifBnckRJCoYi2OCLV7ErRT14YhGZjK9T0GIrlIwYpvqOn8dm9WqLM
KF0vP/nSGWb87Xw9PFdkiJNRjez1Hw+tpfBtM5RewjuFdOlXVpIkewppMe8ct6xlwgaOebfMdm5H
tLmU1lfMDeJogeT8O4/WeV4o3dfZ7LhpYpCuHJ1WgPotutqYckjs6gtYKRCiNt8SES5kvtrlnk/6
8IkHKw5eIPUPDphgSZB//moYSE/t7QfcaKCdslihq8u0rQKrDUkVfvfxVChbxmmCHQDfwcwf7oZQ
WffgWPZP7I4Tn1gNiaLBkuWLTryJamQpkiaRenUNGlxfF0i/90T19I3T05eels80L7zzT6ewDNRu
wGUzf1ncdyfuPD4EE1fNpNlB5U+sj7i9LFjXAbQ+DFijltp/ZeRMmMAEzYORY8qA5nqeJMHrNRvz
+GTsmRclxpvwnEuuHWeH4PCQgA5tr0HPtvIZLxn1d4k+v3b9itT1Ohx1A49IaAWSgNy6I4qRqX9m
vC6XpZLa9f1GyuXYGgp9aSrKqQouAM8QiPTB3E5788YtE3djQv/K9MkvY9uUrxgsY+zKWd7NsQ7F
F3bStc3J612AGfR5xBx9yREz2nHmiCKBam1oZX2ZyQ2yNi8ooig8dGUjrvYHKML6AsfATV459mm+
Gz8A+RZIgYbAF7mut8EIc5CYbUDObLlyQJl0ZjZu9RWiKw9NlKCMWh4I59RDf4vAk+DREUfsvrHl
OLtx5v5Q8f7zzhQDfXWTBa4mhDTWOY3d6IhhNCzJn7jV0IlMe18xibuRxwuzeOGC2oAjm19hOFCa
uqyZFe8CWkREO3bpi8WLvdLJY/5vDvS2cVczAZl5QVIV78AnXPB1MwWjJDkhM28LlZofUcUDPnKJ
HZmRqXSOTjB0CpAEnn5ySyr1IGrGKAIvVcfG62YcvA1gNxTyk3wPGDGmooKRarsieU4xEub+JqLv
pLHKrJo6KeebjFduIgyLW3KE+qmNR6yGXUuuSTLjv2gS8no9YGIvGHTeWsW294h+0431XK+D5Pag
d51zWy383VwswS4YnlKxEnfaEC18RmH27/yQrXy6HIEdA3MIlY3/+BMMMKiKC/9IN7thK6+iwiyi
JSSndWCKtRGuNKG3DJJPDqPf5cMBPgfIRAIxYz9NhdfMeD+bnOBHnYDMavDi+ENeall7MH+RbhGg
2uq37paRToOX9Ykyklti96WmSPrPxqAjjl7CcSzkq0Q7GO6kAuHFXF/tL84yJOwQwNd6rnYoQhJu
MGKEZY1eHsWAq3Qb/YnenNIYR/1I6RuKWwYwm806DvJDLjX078rDouS92d3kM8P3kN/oRrxdZbca
ii+7OnHdxrAQGgi8KjC5tX8UKmM5wM+QyEk5M513XFFmVS3HcZfmtO16vU4uuKyd93YA+wmvr9BF
hf8ClPEGtmg5E6EskX0SYLHYzsdApiMYiaNT2dfZ6Ab7o+28uYvbODKY5qKF7zTvvYK3VOzgKTqW
0uYxUIg0xAya4CJUcsOMmtLq/14AzXim0XfsWCcRM17K6ZZx636xJFUUBPjWLDs0FUltneWGG3bs
D4+BGwqgCMRQVubdYvmdl4mj9FSeQX0jPreZldGOP9dL0L0Peqf0aE9Vc0iYXVcO1LjrPKIDMicE
8AJVTd0EQcHPtQf2LFeBoM//+IuiZDiBt1kGzIMar3XCIwMJGV9oxfY7qb8pzfZ4UTr7VJm0q6Up
8bXaYH4/5iII+QHMMIQoXwyP7vt7/z86rk89bRjSU+XEHNFHZ/qtP/xkHw9VoL9K/2NL2ZYGlB8r
DWBixUmzPUfBcPg22WQj9UTy1+Jhd9Y0vB6/M0Ddc2Rz7l13U5S//L+8yAddA2Gm0lmz8mMIclJO
W848APLHaQJ5qj2up42WYKQ1h8nOgab6dnr1b2lnVfDnuhVGi0Fccc1tXkW7Szzi9EMs5C3toM2t
ed6nGbBO5dDpDG5GSsyUg+c4IJSn/Ji/3PAwoUbe8HfL3Pl95f+w7iIO6lpSZqGHVEmTyPqtklE1
etLgVGsOfBWzQzEkILMnugGWNeCH4VYAyFhXJHOdw/LVZs7tugK5mFFLGf5Y8kaKcZ13I3GGUvmt
seJBA34yCN+alZhqHjZRcdjiOYzLoSW1lQwREdrw9HsLQkGFl6tKOvyuS4uLaLpGvarvUHoEclTc
1fwWJHNDIQNTnCJowRFGezT33O1xf9fJIrqNmfyQ8ucO1LnaXsR3lj7UFXV5buUY21duTRFU8xQI
nSz/nrgYne+eV/IGNE21TYH1qi9m3D94iDkq9tMNCsMxvQxHDoyvZSj+wk9vdShbRwXkS23UTWko
SHY47ITtnPPJVPOYPktSruT+qSEqL8HucIXweRsu/F7BPnqBm7TlR+fbs0VnZ5Kq+0VhtAlpmANc
WnVOLTjrBvQthb7AIEkJMMO4jes1JQ3LKFOO62fGJD0Z9TsOUKSg7Ah4Rte9VjcNqt/BkkkLYapl
rTAFDj0zdi46hF09d0x/dAeud0zyVYaVGud8Umys+OhR8bQc7rM7X1Prrq3+zMGtxxnaTDe2ixmv
5Tphe6QmVfXTum3k+/diY3QStnPKreXJ8oyiEYfLjY3m6WNnh25mnZXxAAN2MEVOjgRicUbb39lx
T8x9G63fH2K7/AXAI2incJa/cgRu4pfwYNlgb44k+PMtfhNHf3Gi0PrJ7JlTFp5SU32mynIxgEF/
8KEi6m+JkZOSXwLJ5cti0b8HcNQN+s/ZH45BmcDs134FfLDkRdOuC/4Jzm5VRj9BdNcShYemCT2K
ccPDOKDUqFefVtgRHqAxTway9D9KFEZL00cAWanx2pJOIDTXJkt/WLis2b/9ILbcsCndBM4Zpf83
Fekeg0MqjSUmnc7XX/lZ9r+MVe859XBrTdBfg95R5NFQLj8w1f5OaHZ4STvijpsRcKU9Vr8/EJrO
7yfaJIjJrBroV5AtMzNRnF7ekx++9ZNBi1n3lVpIEc+oeSShRRkbLKBPx9arpYpjB+GvOq//D6BY
Ty3VWCxGdHYUAFRthENnSMfLstSayDBe0BQoubXJXLZhwcXuJtpYBdMNO5i0wEHmHeF+WXxz7m5m
FYA9iECmToD6uOjpAukKSYHMBkrbX4y66Il9ncrpgxa9P83WJmSXJgPUlSt9+TG+bYQ5pIMVhN/u
LxaMS0DVnRQ7FuruqNEvZ2pyJHOdVTvueBYEWyMtNvW2Tm3ANfJfFUrJpKE/ZXEvhe1UFHUWJ1Q8
L6/pzoblIxM75wEBiB9Ar1xDrhEMpJkTKtkV/0NxTfQwSg0/8yANVZcpZ6veSp6pzqHIKuEEUIhJ
he6/iBAEIimX7oveps49Fb1s6Dw9Opq3VLUTpoLOwH2gqZiwrXbO+v/C8LyBFK8bgoMIAg7zq/xb
eRd03q/hwOzl3D+eGxKZdRDx/vNcliZaJ4REIDDisMcZMcda62ytDhebaOyvUderzrLh488plbtn
vTJ8FfoWaKQ97mS7ff16m6PVd9jOw2NpD0TP+g6ANvu1hYL3pEkL1hIktvi7a2dhApbIUC4ckcNv
Oc+fiY2rw1//OVrEH9/ROVRQMtKiuCYSSJ5gFJCZCNi4bGqT7fAVJEQj5i/rT0nUjRbFpZOitctY
fntdPT3T596ARGBec5CfWZcA1t+R6zXqIIBiVH09r/NresNXpLXin6guEZM53mLkEwQ5+P/PMZXi
NJ8ilel91KHT6JEiP74NVwQJNqw2JgmY5FCx1BwaYdcJsS9+6iVcvnULfXEUzYA2+G+Ia/AmWfgM
owQVEbXqVcffQg4kBW0xJGgDt4rhn+/fkH59XQKPzNMJ7fkzwP+nfjy+5Ma1mdyI/yf7UEiRAmUa
QlDbonCqUNZzK/4mE6CX4CgjTzqdGcGlIYanPMI4wSGtJgNmCMBohw4jVmxIFHuYD1jK0EACLVAH
YsEF4yPy8qmdw5zJRUBdsxVZt0GTnwxwgBTlJYhClBqdw9pE/XwEXN1MHAwxlUwfYxA2HTmLOtxg
Kt8ULjS1L0MpiEtwumBxYcK1v4kDkQaeXRdsfRjL6Yex6b7JqflQgs18nZ1qzuCBj7D3mbLXP2af
Y0d24Gak9N322TJDcLhjLj4VIUAPVlZnQqyJbDq/rbZ9LFuw3vQ2ujkB4eSW6WnXQh/nLtEJJdAR
UB7nTbcIhMacG7sWdZIxQJrZL+YOPahOTJQqn6ebGJuqTQZdp7bqrcq6GiziHKioA+ETq/BJpijk
VKdrd/E6PukZgVXHyXlyVHpYPpYgp1pq8pKynZfZvpPbnY+/H4M5Gl5y23vJEDqkUkTKOAyIgYNp
zz1pTNE4+h3SKmewbgl/U8seqEFkQY7YaVbOelpk/2TD0HKSYJjay6/F5PYNNjDEVNIahLHvgDnZ
STLQG0XQIJJmw1wCcdria5oMuvJCkZbw5g2RmmxjZ8HHy3D4hgBaw7MTudytb0Ismsi0OReCo4Jf
TyZNRpzLxs1M/lAAqWD/POXO2ZOjTvNgFnxvvkV6Bm8/wSCtaW9ukFe8XqtbGROlhhy8AqpDS1cj
0eeYg+nQKokePzmbiPibTHOF95jF0WB4BPsQUKh5eryxzit176TWIKt1gu9JB4ljianYlmHERMRN
hOktBSA1d8ip5lisgPyKhGtyFG4MEdp9noBJTKqMHh56ddKJeHJngJz+YhSBWFbNhkNjFy6R5pZN
k4Uf4jJSN6wXqvYfdVIdToLSMBTMmvLRfkU/Namv2DXft3dTxbq1QLIW4E8a9pgWBPPmjwXlqRRq
KmQOYWYhoPHlnytqqhNePDkE955M99EmJUFjjVI5nGrmIj4gE1VXiyXv1kkLwL5Mq1qB8m5pPJ7o
YjMDiRLav7P+V2YTTMhKKS2hmhic3hub84q+5Scluh9CRwA4+yaVbYPUgF63itxBydTy5oFAYNay
XXGU8PdAn9SIGcLQQh928DSbJFF2E+ZsotX6zZ2xkQ0T0wYOX4KCQwqckiMtUCsXJxnEiUN/sLT6
/JJM5uCCvwV3N72PMlKngRTUwfd/Bn3LXY2UjV78z+lXHPU5Y2FBRZefE0xdhD+5l0OQQD7ULEzf
kLur9G1CANNYAeFLx3BGH/fcsgzfdGECPoDyQSxMAVe5HUK9sE/yCdNsn4EEaKy5xwpFyZhSuntN
KdeiHWxF43nWFY8fjYtrOiDNKlZN4Y3d7Rz7RkLnrgbewt70yIt+FbVtw2jwQmeUULyljALOjHGU
FhOG+/U3Xc1WbXeLlwBuc+PYDdbAXll1KoQx0pOWOl7cgwajMUubqFo34i/qhggJL0CT2WPUpEZg
75IuCnF01MGz4ISuLMkdUdJM5kIiyMdjpT8JWnvSy6RLFhI3dIay8tQK3QwpBQ+eHUftQv7MtuqT
5hkJKJhSi+yURm2WbHz0W4u9DltWn6dkaSkua/iYKegJAuywx0J0tHSi4+PJrIJi16pzCwpp9xPn
Yt0KBteN5XEEuDETclzBnzY5LZ/n2pN1nIGBhKRRFBpj7UxjFavfNh0JoOQ61/KmpTNsfHa/8xKM
EPYR9O0IsOwGE96pp5vOrhJRJiiEqEl9/r9PFCHhRShqIss+iBYxxIkdB07kZVsVQIwUor5JdimN
9if1lnbYiwnr2E8Xv/Q3uXlMEd0q6Cin7GB2ifL6gzUZ53Lyey8LQEbTiM9FCYW0mZnXpHALPKo6
bGVOMSssWtE4Qt+PGkoL+bq5PRwiXmO6sDBbgK1nUHY2TM4yUslU76kbAXchGX47kPJGI3+o78aK
yk0nxgIOt0izna6FZ6dlhMaAaycLM6OaAAECRH9mt5tPFPdUxBIFlCX7XBNEumYHNSPa6zV5b5Hn
kneM5IJq4TqlAjt+CESk3930gQiCooQzhUNahdJxcdVDbksJZ7+9FEuFnzU/vtAwLkoEKo0pSNKY
qOoXGBGUFnbhFbgu2WtfqYpHMZQ3oMNfIjYt/7AkC+Vba5fbvv4i4FGfh/Nys5q6XvwFw+uiOSUO
zhfAGIjGgAJEwaPQ2lEXLSOSBkzGL4Za0PGhZrYCLB17WhtqfyxVziQLLU92dXCbiAhp7Wv3yv3Y
TYcg/woeWc4unz8UANux2+Jey6qFtJpsA1coR0L39aKTUsBYytF7WbaJ03EhY/imYGQXJ0SjrV4v
lgfsBDLPcP6b/enetvmS4ZsxJV4iOlLxalznMU5hChs6NdPBRei00s6+OlctXXs/0qK+oY4eK4bU
xINYu+p91B8OD3aqBDQrEei8tcYOMafY5iqq97InwEbJ6t0gqwepDyiNMHDDUC2ndR8u/AKkIZew
C5SfpcXrRLUnTMrPVeCwGzi8T9ksKvnEzff7uTqNHC7z2TrwJCe9hxP+yCVv4HrOUU+3MqQTxtkf
9+Ry+GvqLk/ShlVJz0ZU1t7MaeBpT14Qk3muMJ3zbM2Sx6Y0ifBJ9gkA36MHTcI/AtGl24cT19Dx
v4IPdKL1rIRCLZf04I6zTBQOQ4MswNrL055TF2TABrR5LeVUOX+2kncYhXyvzM6b/ARP/Xg5jcmp
gSMHkcPWuWLOG0ZQ8Lf0tlCR9ef9714bnztCpGJ7P25KXVeOugeEy5YqFjs7ioTn6UcQMvGEdRe2
3Y0fAnRmdwwskUCpm+6m5KDhB/quDVzzMicK40OZEp6a8cd+fwCtkKrfBJD8ueCA0iCFp1SZ9iVz
aPTjOj16lZQAGt4Vg5LN7TzeG32m1zAH+h+v/haDJ6wktp5mT7KNJlL7yB4pd9v27ll6d5KP7QRf
oufWLst8IAlv8P2WNiuXG9+bEwf9tyOpYYtTqDx+1ECOTRZFB1yO2xOZjHQZtFTIj8UGWHKFdAoU
Qn+lBKncE0TwXd03l8NNzgN3jUuMywcFsrJWSWj95ME4voInnKX0Djf/yaEGQP996AIKmwPiLtU+
MgbQtyi4esXzbBuuSU4iUDYHbIlRn4e0dofiwXb9EIaUlcdaeOm9IqQZVz01ckX96w21KaPfTKoB
mPjW8f1eue65yKLcEQ+KZ5l+d6jZIPwnUFlGbaapSeVs4O48OY44TRJcHT29bjmCUUeBAZx/HsSU
v/8D0Qwotz585bscqr6NTBD/U1EHtXqYmqi0UDQHMUlgWONW0Snxvnoy7bvuynKeag22GHnRNadg
9kOomq1Ybx0mTGdDxSNW1WWmWCEl1GrSxqVhgD8Y99cr6sjkW7etSuBM8l2tizhmVcYLWFNUyrtO
cd0usWydW/64oeL/20JzKv7MEX+LOIF90Wyuq/bjbZN8e72yPXpSu/wVMnaRYX1UQMNWS8Nfr7Fh
iU5kSysyTqDCg60mdmonUgtx80ElDfiEK7LtvHwvTWzaiWYmlH2sIhalotm5sZYynMCNhkCWgLpI
vNa7mL7vkqOnHpXSReo+i3b9wU+atyhYZYldS6YdQzcT8SFUzjgYj3VkWDHgIZcSx12vrBKycetX
hkJ8sBiCCAb/ftQegoLgY+elqGpBtucNYRtu6Hh59dNPvzVRjZk8E8LcdyHjkKq3CcQMvBvGTgwx
37uKM1X1+GB7HpjUC3Q3PiHZoqk0aYPxJWD7t1holNcUnRtwhMXhj19VWoYNTSrz29QZw0mD5Vxl
GZvx17ClR9N0r3wOHoI5RSJ7loXMr3l3juydsu5YZu7nn2khw45hAkPpVgh54E8Me2kTftgqW+B+
2eeY/58nhHZvVUMEz2E9Oqa3a+eWP3QqSPJ+tInpocnwBs8JjcaUpJsqZ92/Cm9hrCReOYNtWm1d
DfcPzKaPoybFOwZYMWPxL18yFSeFqMjImHmCrIpERJw+nYWS2NPElH3e0lZEUECSPDVvwaZaS9mJ
HWFUHXEcZkeR4BztVafdw7LpqJT7u5WaelhDvxXLZE6zA4rxRsRQbmsshQ9OsMixkgUsu/AoqYrE
8JXxLtgIHbrr7XNCGuB0/MPFEX8HIV7jKjnvNZtJU9QwN6g9WQqzDUSvQ37U5tOOLGVIk1dtXPbJ
JkzPMQPqD7irHelrRSI/JD0/YOW/0JP6JkY//ewJJK3h9sMbVuTJQ1cDelIS9NOFPzyB8TygPnKp
s3RJJp/waaJXMZ25Ioz80nne7LnuQGyE6yCrtmhkjzW4IDxjNzTUdqhAmgO0iBYGyDmHtPXcGieA
LAafgKxUuFAv/S1HGxA/Ph4Jg218Dp+45NboGRKtehqdNCo2tJKwpKm2z63s1zyPusV1tkfAsGBq
gVQhxmNTyBQbrCb3w3MTdvrcQko4TfqlIrQRYE2VFV7Ay6B4OnDJ23Ppn3D//1L+zE0IYZa6tx4R
GszU3iHcK6ztV9769cPrkIbV74lT9bMMof80JsX98KWEtftYYzpJgs9ZQ5vd7pRdErJFcUQJLaJB
c/YxkFpuR+7hlQPcUAf920DbvOUiIajwUcQIVgxJY9PpLxBLYnbyRAcO0irdLZNpmC693uBnoGCm
GEt6O+D33qCxtKVZ2k9jsnPBrpMKJXpvB8mGjNijePCeYG1ti6S7sKoi27WjjiTtytejW2Bx45JK
AkXiKZWZVMvVaBDSHUIVw1L7Uc80XNUI7FLdfzjLb0hsojJsLHEF1UHSm2ay0N1Cl4BtC93pTr9I
HdoGMRTYbfyVCyrAC22MIO7ke6dcmLjH4luHlLkMipBqRM5WZ9pM6oqj0j34qH3HZQ8XUyFCRH/5
DVGr9B1uSg6mGH7WtqgQQ0mx01jjXsIpzsZKgKGSCBSNk2TyPSuAyy69p5RkoA6XTtobwbWdHOUI
LTKUTE4Cy6Azauvr2BMP/oED6h3uqBCbORXhxPQ4Mv7Y9LXggLLbCL2uxhT6hf5QFMnUo+nGs8Xx
TG8qg4teThRgLloaqBkf/17bdOTLdhR/9kQA9mfNerF0i30lpvegNVyCmWIWnl5Z465oGxhsemZo
vSS3UO9dImZ6D9heLncTnEyLF2OWZvIbytAUoMpQHaBeQVLtV7Fw2H6R+ebmF4Wj++XLvUs+uec+
cMoGc1uNRGKilT99chgX0ADDDcvMr9hqt0tx6JwrTz7Y5ixjpAqi5UeYUHNTArzBfrKpRYnMkYHG
cL+Yw05k6yRQAz3PhK46oNJ2b7GZKUT7vr/m5jb6uBzdO356dEGpOWQbKDq4c8Ip1jSsHxcZAAVh
wOHY0KWADi5gSmEECPhbfrYw6GMoG3dXJu7IBwW5dfUoU1o4SCeFwLlsaitTp8m7T46OysOut5XT
mWS3ydK/IQkeErab/96nCiR2JmBxK4WIj5Z6pC8lW8ezN/dbheEo8GugTlyupe0BBlA6h//qI72P
JMt3x+GarnDgaBHPv7W/AV+A9WMn2+MH9D2wBmiDoTieMJ1XRrfBdqg7JW9vqC6YTcJD6+S/q8tx
5EKWvzmZLzuQBMEn9vxZZq9UCp2eU9gwisG/shR7XeVIfwGyeTQ9nX+Azk5HADwAWXWiOBrOd3W4
sQEFFU8oNjWxOXS2GEsB/GBWk6CDHjq7udMToHUbCKTRlpn7/o7VZtZluEbG1On8UaSIb6Ubt5g2
0s1wmybVw+lR3OnbYoMSfTyFVJOIf0n8eYV5Vj9oUzE4Ha8JcJXU6U6R31Yy28RkTtXA2E3hEzej
PDEH47x1kLwG6gH1/Phee/a8rWtW3YBUsLYfqD1tdX1zXt/u2AbA1AajF+zW0HVNINo+c/9hWdM4
D8Q518n0HJu310FafwM+8gHCcs1IydkV/8+dsuVYKIibH/Wa9OxCeaebTxOgEp514uX2tZ10hEtl
ucmT7YZo7IX3QNZ+ljYgFnmI2kRWEpn7T404upclEJg12QkKGoxc5TRNDzDZK+boW5ry46uWoFG7
rS5fhC0H3DiEXhU9kWJ3Sd3wFD4NmzT41flaUCOg00WhUuEdJYsn80yMDx2h3seXJ9eGmexkz6FD
G4T5ppCo7A8GQVtQajr5rsHL7wm2GSPsmztQjwGa+5qFI9RZAS7gQU3hUVB9nwNz9uJsVrBHFzTG
aWCbLz0Or1R6QX+OPaZJ5k66c3aLjtowOyvkNz/D3rB5AYSc2wYvQUuei8dCIkI40WDBAFSTc4/l
neKKrU9OjnQA66+GwCWJmvi9Y6+NNy7WS6hrtb7vwwHL7XCrywPxdR0ijZj/55I7bZGn7VLAHM2W
s5G/k/k1h8998PrqZaNcmrf5xYyH94BdQSAq9wcd62ewuteqL/fCkQMrmTAXO8xDVR2Ec8r1zVcE
VuAlspv4wCupbYkQH9tqWYcKmc0uw+s+4Qa1upiBuwEVn9P16NLc+0KxwD6SKpcxL7nU0I00MeCq
lRJbb3A8/4e6W9woQVIjbAE79i5zGhmNxNRiDM0knHJ7FGV+V6KBgGFHFOIV6dho0D3SF7m1HR/j
zXy8yHyYjPTxJc5s+JqwFGgNx5Cy5nPdu+5bV0PAFUuH1WeUJMSPQCRY3mppc4eY/Ig/6r7NzVRw
cdqq5hUk1+m5LKQ+mqs0zzkYCo0jsHL+ViYx4i3CW6kSzZWNUQUBubkTm32SdBll3G+0TKL6xyCq
tVhxogR2kcOAwOWTj/OjxgJUEJtH/UaN0PMOhTAAwSS6b9h+YedZ5qF+mPCGVOH3xP76UWlyytiS
B/z9pD68HrBV1S3rVKdcoNcfNI/wZtX7jgmWrasY7Er6C9NbJ1SXmpM4dVtEyNWBZKRMwKud0zut
KsD9enzBYkn2uo8Zs/bV28tUZAnvRdDB4olI6hcge3E22GjwhnayNgURgif2CGJPbS38i1i8D/99
S9bBdCorqBrdVwFB2S7p6CEVT6+yR1ngztYznaz0Bki7vGCsuxiq53rzSwhGVas7uPOi5nV1pz3K
1eacCrwj8ivi0IbxDVLWWU+/tA8gj/9N5VAOqHJBjkP1ofBg+HTuf6cSgnfaXbhNzk3CLIWil61H
6PbsCpYgicj41N82A+3UIyGfKgiyjdnbaY/c2J4OlawXxt5gu2AIopINkgrplfLKlX9fPlOYWggC
Q30vPCfU0Pv2rwSOuL+rD1NzZlubLTprInOeN3qmd9myNBvtk4o+RlGuOqOVcrMI6xmb+K6deZtz
/Q+sE6vtG7i12ly1NmVBidg9jkd2gN/YBJOZ7wM62xDHg598zMNyMQeBHpr49r2CAvZFxQNF5RaQ
xiZOxmwqe6s0+RrTZe8fRH1xNd/y3a+y48WPiOC6Kn3N3PW6bWtUFJi3KKhlFKqCVNA8qQQ9lZF0
6Dr+kD7fFJ1snlHQjsv/lPdkU5t+9IdTe9RkCptQJV8hU3WH8T7PsQyF1U6m5BSh5IUg2CL36wCI
/YVwMHwx138MlSJUxnnPvHjCmXtHm8XDzlIodakEslhG8B+2ybwNbBc/UWpUbpGUHcZIs3TTQT2E
IQ+QFiQ9+UsMUcKmYliGcxDvAZhJp0+NnGx4+7i2/iS0Urvk2BMr4gLSt62B8LKjK8eemrnsDYmJ
V1jHA0xlXun2cVUQI97eYcs7fFd1PZPMDTkUCv56po3hKZrt2h4pBGf//V3L/42lj/Kip+LKyOXu
eCrUC209V3HD66U5rmtkUvF3KXO3SBYZSxezPDIosd3AGMo3AdLgCRyFK7ZUTyayizbNzPlT+G0l
lYb8LFcitgpDp1BWfqKwElWa0Iy4gJ7q1PTmeHNASpFd8cw0I10jQELdeMEjg6Def24SaiDgBayW
R+LpvPtfSqJoycuj9DkJuMdEMSDHk/K6tXffAntgjk7xuXO2rvGuFP+6rCvXyafU3a42KXhGMoYL
1Tr3qHEEHxcNcOX8Mawh5XH7yhfuYbjWnXbcir6OKfVgkH+bqCsqX8ck7DEHhwAvij7u6UrhU2Q4
k5q6rmk4VzYJG0em0PFiSRxIHFwz7IcJlcMshrys6ZObvay03tMKn9OGbzSnO/lCjr0nRoL9r4q6
RTpNpXkUi+KMcQy5AjrVHXl+eWNhyZ4wnLzwUc3oJiMsAmGZaKN0wQWwItrDrHtTC4lx8F4mzZFp
BQhit7sIUWwnVyg5l8xZ2al6aawf0fSWhPlgI3Wajct0WhIUuGOyU+7QC0yES/HW9g0GeDkIXwcR
fX1VNKFv1+Bdp/eoEgaLy77eBfp3p5gbhk/AgYe+4gSrYbMMFQYXCHs6IYkBBCuHYJZSxx4CmV9K
1J0q5v9RrFYK7CtAfd4SpbB1opXqXPaByZ9jHY1wXVbMhj/USEItTX1+Z4HvuB6hwmwJYRfIv5+g
0EbVwEeBYDYEaak14z3tzG+zpGvXuW3b5VbX9PA8KcmfUsUqVtgWkJxUGqzIeJhSPk2IS+eLzVQt
29IJS+URfWKtvJ7L7ahrfxeDZiH4nLAujkKSKSgvEzFAhIpOVOVNKZ/utmoaTjMGa4MU47UQJe+m
gpqTO3dF81uYltggWKWP6QnFheSQHIKtCALFidVqtqwxQcrlFLyePXWQnwhnwXyR/fFwbfxpwpYU
PdWcgFhyAE32jOjm1dy0GCfXDkt0tZKR66/Xb6tGXfmIGjuLPu0Pf/RuoJkk8bwwWcUcoz1pF7MP
CjnQDHYS3KnAvQrOay67qD9pl/ADf+PuX1T4lENyXH08pIsW2n/cinqe3TaQTHIRe+dgPgK8VkQr
S1cuq3WaJhS4FkCNt+p+kX9B36v0qanRlOy4gcYSONFjHe+Oj7YcCEdhu+8slQAe19SVEmNlR9uW
biYPehWb1Os2/neATUGZ2+cXeVWFAeuA0Im3lF3dFcKVH2DF69G/VhQULRiUcKpUAexD0QoP9AWN
2hxWTpwBTIUd0+NLZJsIktbdfoerChynKOupIwFFWn9I8B4KetKlpa/zldPPU+gmmHchmUPaUqvy
btJemy7btM0HGs/BzAw7ulNm2TZCNfU1h+g9sF24ktd5HkpZdnbdfKYSfrQtN/Qa+TY1yhkFAv9v
DbAOYByRq8ebaO4Lg2lkWnNC+h/3MdZiUYPuCxdG/OisNWAnRdgqJ6NvufNmyuUY29n2H0woQJNH
SEq2SwfL0Ld4LcoCOsO726Y4nCYFuuQSEHcqmNEeEo3Ua0prgtRxwEkXfJD7YhAbD14DnY7yAftY
mNsw5I77Wox47dRM5fufis755icRJW6+zH0RtQYnANGsSUSFnEybkMfpiXx6+SrO8WAqbvn768ao
YUf9mJBjChAxFEYFtNH2xC69cu4txit9udmQmSyp8Inj45nJbHCRDuk1wbAw2sugsTmieMa4mphY
XoWf29dppFkiDOAHVv7vCIVno8aWrOX69Yh0TaFfGsCKEXWYz/GCfZ2xrg0DgFJKR927E7xHCZyX
XzDdAJWMLIqdJNPX8MGYpLXRs76NexJxRO4UyNF70/pIS99vSUeozkJNczS76EZZ3TimZ4rV8Gic
gu+/WK1AKVUqiZIUvKcTXXrPWq9xfnNeVs0R/Pl/U7zQCVUlqNkmZpMmVZGBN09347R7Uwlb5AlW
FIPkwo/502s0Dq97p4MT0NZwCTrkKd+ZY5Jmt7gNHHiHDjIbc4glY6r5Kc3HY3xYaCJ+PxzJdnBw
0dY5Z+xGqONHbPDFTCviaWHeMaKKh0tXOJSw8vcc2lVX6rrTNSSWkw9PpM2c66ld8n7Tk6/bURXY
I8TixQccjghtWAfEkWo9gwvEthw+M/TX9HehvTJL+Q6VTzjH0JxCQj200NuSQq51Jg1QvHLcBXRm
zT6rL7T6YfZwkCCHmGhT/nDhClgaXKn4aweaMFUo0+LEdd3gqqzK9QGRyS2bPeZxFbZomWNMVvdt
ERLR1HwJ7uTLXAhmDCgQExg2VL+NkOxTRrlXzCOymSispgLPbaemDYxuAmf2w9PBT8MmWbPVCh/b
8Nwdr6pArqVOS3Ar4FfNXjzqiaMi/0+hFb/KQgJZgeaoczGAj7pzwTBvpNH1HdvloVNrSi4xErMz
76jB/VwzAczey0jUoediVsbz+F9GBEE5So16yHTjWeTa++TR9DSIThBKr+1EakkEnUEIJaNhBiBo
DcEWh4TAsGS0sdFibPJ21KI+uyQZjc8eFxS7vOEVTqkQUKC6Kp94wGTWbvfX5qUuvpnLdbCEPnbP
EL3YeU3jw+SuKkirGqtz7WGDAYl+2eIHP8UfE4ucoSc6S32RZI+o6k4Ehm5v2zYLGguMs1c3iMYp
zAcGHTUg25H28MTrN72gvMPwF9QYPYxg+UkaemHWYEZ4ti498deGKjS9iEIlBa0ILYG7J1+NPj6y
Qf6MzwKEyH1BBm6JiQXeWWeDJxqXiXnAhkyjcoy895NISf0VMIIy3ogMWyXVuWTQdi09W41zvYQ6
LnKUXsVROSwE6Q1SuboLeo/oBie3gEuCqmziWsI8syehD33fMNAI/gNXwu39qDy3BQ8lNqG1zv4x
4xmZsvK0CTAEe+e0pRFnpC2NI4/H5LHIYf91DFVstCKCipGTgcGTSC3EWUflrjaQb9QHuekNctyk
7rnZNaRtCFGwtEgw2SUl3A1rdWoBBjFRRDMmd8Cwp5j6U0+3J8xl9q9LR3X2dNNLs63H6J5/jzH9
8WnHpbFCCEkLKMtliDefTQO1QfjHSk5/idaNH0yD+xRdddIUjXkuXOslWNHIOKkTmOwt65kekkW6
04CncL13Uu7nEOXIhOcJTArI3OXzZYH0/5R/oPCdJio5GSjSQ/MLTtov4FkbbmYDr57aSDB+59wm
BvkiteXoc3+d+6o1jT6l1u/VWCEWMxEDFDJNESjv04rf2V+XXH9A/Lu/9PRsxvc8+hWYKZgn6MJc
VUiRpfwdH6CS7Xl/hldPY1UcpqjjWuu0SAEar266Yhm4Utfn+fmQp1f6TStK7O3mUOtF0nsyNHFw
DyvuMQuweC6pGgEdZzuGEUhoAiDqF4MKDUrT15GcaoRy3SFHZB8eQ/0jgItXZk5uMmdGw0rpQNh4
Y9bLqDWOj9vR8I7TQt9AKZXw/T6B+TwRir71d3co6LNjvol3275jJYLyI/WMjqceJQkNO0TZdvAs
8HLiu/PU6q3LnGhuG+WfkttriVCa4bRSxHWhdCOGzQLr/6eSrPJHGWgzAfIUjLG/LnKNkhmd149N
pGi2xg+0n88HviZ0udAFMh8Sg8XWfDPLvftQKATe1bkRpFZxsYP3PPIxBbfvUZmXidKjgJrexDAL
pWmJwU6/cqJaeh4v4iN5WrD/FhKkwHNSi8KdWTXBMm/W2udcavfplNqlsiQ/p9A4awjGsiR7nDAT
jppO4FU5O6uqE+gV33EMf8TbKNF5gYb6UpPZlZrEQn39tZeNOP6fppyYbvyG7MgfguScb5RjIgfr
v4OjMnkoBTrRAj4T0eT/wapPJYpo3fZwcUIUXIW59jK5UnCSytN6t5LP0wQEJeU/9Q19N/YNdiVX
mCJfcZUuUrGx/7vTkHwBhmrjaYZfGT1TChAxpXd0wWcvF8WIsOmsl27pMC0O3+LrQZ/Ju797rFgw
HntgOfDX0jvm2VCbGR6OHSX1hjX7Y8rHcikNfXY0RL3idRC0zlPWoiGfYjWSoDbgG/La6kObzAtR
qCQ2V8e0YMRHCX4W7VxHxuohn9UufG+et9UOrpj0gbZhCovA25OdEYuVTkwslQ1Jel08KzbZgeii
Beg6XD0d2vkBBxLb3gyLTYQY26bhL/CxA8zgvFAw9rxB53qYSOM91t6pN978oIL9AJTN2/B+VyTg
zJtywwUCN5wy7VxJmmt+QCRW5J1A85Hv2XSKGhdKpccJSNOuXWK/M4fjlVz72TOHklkGiFXnr+zD
SifenTRSPWimfrjdvtNG9SMg7LroZZVhAKO9NPngTVDrj6JyZIEunlOsL8TuPSahrzR69IFmCKGa
QlCfJl9AmMfSarOeEilDTUuIv1P7weVUfKN5fQrbDyrUDDawsywduDRhKYxv8HAhQYmZAUMASDKe
lA4LCeE7NQEoqUeabULd7XUBCMreRCiM8bPdK7f+asRqiakELW0GtPSHKuYqIZJMbhE6luKKUF5n
4PDWQnYm+rM1ZP7zmcJgp1hZu6E25s8ib1MThMfa4QU0f8RC8w2+P9IYakDJHWya9GA05qp8aWHp
ybTB0CKakMy0///mxeeoaprJBwZGte6nYSYbLphkq1woJi+nHci/xtEWtnXs4lxjPpoNA5pzkdro
mq1Yt/aDT8P9ihBpsq+jORGT7QLk4SrccPNX43/kp53yJ6krf6BOx7oqZac2OlEHRcg9H5Nxobl7
oUT4/1jBHFCLQz1Dn2LRVTZUl0gJFmUJyOa/Eu3rnLIHJ7M3AczKb8RRG2nuqSaT2ED7cqs5oAGi
46rKfEpzhUqKUZgHOd9mcw27y5y+l1kvAb7ZIbfeJzlAckklxHGo5aq7QRwqPt5gQt/uESvQpoxP
OSdifVI7K5on7JMZ+83KVQW1+LtIJVurjTpsOHc7CCSJ852ITST758YRkzjqOxIXNyeKKhT27OMs
ayzYkFdp7fEZOp/T9cjydelT6nh8go3NsWv4B4bobmhrYHQa9OXMsZuDvQA/IRzohaqdXcSj4pDI
ASVBd1MBY5zpcS0jUtCdgC/RTpDpx631fFQXk32v1eqLi9XrdgEOb7gHcn6+KNr3mnTFjVZ6H2Kg
ZRQ7bKaw0F6lpYzgQAsjQ6VNuT8ghuO0nBXr5uMZ5GvWVRtpZTHzMs8sdxMPBb1nHmzdWby3TDOo
RUkBgSBW4DbBMStt3UjsknhXhVkYmjYGpIydPW5G7VXKq5EaG3jepIVI9NMTHeTOKiK8jft88+IG
rYHzGe51iqV19+7tMsZgHHHDd3tmIyHCZpgBIvyBg9MkzvNrMPJn3oQ360ubiCLyFNHBYaWpGbJR
YKEqVhRflySocF9Y1L/da/gnzLnonwdEdf6XK/nu90MCY7NwB907ZT0NNj/pmnl3tsMWG2OtHBt7
HLN53pdjwmaCrY/znR8iWzOoOrb/RIsmRntvRwz75IhKnQZ7aO9hPijPn3AxS+qcpxyAsn3SfOOs
glfc4S8pXL/gA8Gu1tJq1xdD7k7vClZrwaVde3YdjnSwpCn6AVympEyB/ackKSqGe6l2nBDETVlk
oYPsjxi1YmkS8wv19AXRNfUJNs9GZGqaBQ/PWXUYsPizAgPwQ8ATwRVz7dgnuJ1QqzBBBwzl3Nwe
N1MRa4LL605m7+GSsioMwQ48h/iGMQ23WgVoRMIJ5nsiklhJKG2N2zbn+BxO7a2O6DjDB+R1Zr1h
hapr5z8tHwKgCbVocbTR1kpoeRU/fvoxgWMN//JGIKkEFa7gQOfkfkU2eY9O2pF1LT9hfqx3e4xq
c+9ohB6NbDMVGNmT1lhiTtmR9UZDZMAhwddoD2fEz0e0n6d8SC8XaZoJUNQAbu6TGQz59VHmcFc2
Lx5jAgiSa97GQqZnS13tF9PWDrIctZ+7MADj3IyuE99UhVQO0IBTra/FRtLNEDnr2xndPE247iYw
03BFoTRJoazk8tvBeKk3ZJiwMYPOn6cBEd656RuxFkE5AmSW08SfC6pKsLXc9kMAnxzTCNSMzPFC
XEjZT3lEBfK84zQH75JLVNqfzgArUUeFhN0AgDQgObgQqRLdh7GOA+XYjdnTy0PV+Zw8v55+WqtP
x4egXJIjw0NieJoJEARgu5XJs7dLKrYF/RjJMbKEwDAiPDIfNutsFhJ1OT6BXJsruhDxFkVxVpZH
vEvXyVATRnFONKOQDqPSVf/11NAy+qAQmaFP6jTBgDD4QCd3fhhYCYBRK4IGQRemF33wZw7jppqU
o2l5yOTvAz/O5fYlLvj/myEmIWSeEdX+EZPdFUN07goS5wHk4XyjAbSPrnNU5TikbGChmM4wguJj
zcust8wDNP0K+1qLuZhbLOG2ZXEMyru1bucLM8G6e8Cu+HhX/7zI/1ejr7eJSD13f5N2UcvJGs81
fTS4x2Dyc3gKqd0xvWhr9Os4Ipj1Ue4R45Zr2j1PoJtfyJUm+r9V00F8LkDH8vP7pkPEjgSvm/5L
EkltWY1+Gq0VWxWwHtH37YKX3Y+Lvarx/Y4xDvOdM21fM+NfzYzz7ldlWKosudd4XAjVcglLGSz4
RJ6P2HB3zAIM/soyJ1ebKkpM4Hf9kl0LHW49FGL/iJ2LQQ9a+49mmzTOYy6xwvY3poWadoFiSUNJ
uLGdv8xE8rJXFgNkTn2Au2TR7OaowcftLWmYnAlpUPm/xzZB5uuXVnhYFUjI5xACt2ymKPVz8Ynv
yQfWCzYg6OiovzYDKW6O3s+bERBqMV7NKAIeGxMJDeUpoi/FPO5pef4JTUZFYjFrckXE/OJShoHx
Rv2gUQgH8p+sb0rowP84Ye0tBElZwmowAbPhlHgF7+d94zTx1wCiaVtxs3k56VDCDeEcTUNckDEe
bxj/XzZAcDK2A+Ng+iwuG/4o05uRY3BonRglXwbIYVK79ATiD1TshPovKsBOZoutdGNMb6vIpa4+
XZZmb/03gXY40Egg4Np1QeQPNPy0bzvEIk5vEz37mTh2A21ev1+oOfbAScqscGoi84ncCH0M/6eN
pECDOEicejYWBZXDRnjz0mIPNHPUIwHXhTRtW8MI9hYhrGgH4CJ9782/4vJ995Y2tx8oeeVgMmDW
xiYcQx6Jcbaba7jMcNnhCAXH+TF609FnmBKEA6rGab5cciOlTqqliOznfKFC09Br5LB/URyUay3e
JWKYhl0A0lCZC8lEQnm8W/mfGe7kVuzqbARfsM+aYzOc4UqHNg1TsrBmrPAildSjqKge9WArWXOd
+I4tuWbW0XGWzsnpg3dbox4JyKN6iOTpGS5pxDokdUYJXDevgij+diSai0wulDnDmQkrUdHTgeTt
pXa9Y0StSDeEXj8yg3aGLZUA0iGdum2DRop3LXaHLs77JUymQ9zYsuvq35oCMJDt2po5zTCS5YTW
LhWWswkWQQSkVoP5gfsev2MP+B39xGKrkH2wejx6C0Q2WBo6rXUrNkt+JgeiG6L60BYBea2S94j5
J6C+ihjGcbOblrHqh9alsUJIjOCY5ngJTMXbrLgtpbrBUjqsCDzv1b1vmWBk1o/DsOaQiSe3uXTi
cdmGF0hmPrgDaLCb3Bb+Biet0y+jgH3y2BtLk6iegsXMMBOYWXUmX4iRBSXzWA617PVF4PAZqMgr
1AlokcXB2y0RlHhJn+uhp/omQQlFQbP2zKBv7+FmcZm/VzTfMBn31Ltie5pJJC0WYAyd/YFFdtZW
EU5NL7g08pGIieRYbR8pLWP0BmvAsaZmkNYaFnSYqL4XkJKkGWgIKgEJsYQewYlyZsMe9iI5cpGt
XZ8Dr1up8/58Oa9Jc8utV55NcJG8bF4fWtMzg0qu0k1uP00uvsZ7DHnhWKm73GfbJQGyJoJLUl1R
37AwZQd3pOmNcAbirXrK4XBEr8DpSk60V7dZcJLA1La2tHeBNpgc3qTBHMV9kW2n4FmqO/2hXp7F
n97bBQ53f72WpxBCHreTYSRK6CVtOFG5sFJBZq7tAXCmv2Q3JnwcQgGN2NZ1t0b8mRTMoBLnN64s
WXw9jqbmzdrfLj8Qy+MW9vuvZvpuMGyfo7xl9cMXDZcfHHdBzRgsgpg//KZFyT9HyC7uPshRakqd
kh8vgBl/NT4qYz6Pg79T0FtlSpnhNf9T0HUPyJkvbrrJ5KvcC0SMRhngY0MLqew1gG5bjH2kFFIB
BvS8pWMLRsU8AWCdVdsqknm1BJhRKkkysQJZ0zCR97m4P2rLX8Q6air3A9Dc5EL7LcXU9WDtaBFV
e+ry7LE5gQzK5nRi9Tu0bEa1l9BT+4FjOBG2NpmKxIzLrQrrAE+b972O4bAoLQlj+n7cSVe8r/BD
lYBcW24HjWAgaYZvynIGIgIvMVXDeavZgcLjFeUyKuPUrghV/3P8EZz8bYuKMY0m7SZts9LlwA0e
SlDwHsp9QhAIUMRFuwcJ+ktALBlqwanKi/hToovez+xXBiLJT7ExpMG0IhUOh/Ws0I2qDY8jXZlc
RBde6bl2Zl+lQva62LbqzXpOXIzAvw31rW6a4NgLEDZ6mUcNB5p04r7a1Lj87RwJtq4QvM31tnyA
eJMY+BgVMXCFoz/YW73ZIkQhoy4B2di+qgQHz5zrPTgcwXzgDUv+qm1w9KkX1BSNETe46fL1idOd
YpwFNaW93p5HOQU1XRVggTc9sIUH7gcV+wOJ28f9W3vB0tCzIkwqzMLMgmg6ysuQRq5wIl3Nbczy
0LE9ApguF59sdce3MsKvY5g8g2uhdOw4iOMER+CTk63IjNProMiVsGV7L8wgsaLPbQyR6+s9E6Oa
+jutCV13hZ5+FJ6agOX4w0dZ1Cg1ZHdMgBCfjNO2+ieVbOSNqKsgQCHBwOgO85sm1hXJ56fYJS2I
iuMxzZOl/qlfNZZbKU3hmTDnpjV6fwdsjVO7NPgLP2+67L8LSkdgW1OoiPny1gsBNhF9dCPIZ+L6
V3yPTtT2EDE3jxy59zuerj7Yzi/42z6QS/S9AUPcgBoxWrtgHLTzDA4zNx84/6mGau2xPphQvQBz
0kRoUSXjVzA1kZc+TLLzOXdH4qrE+xOeCsJw70smvSX83FL2a8uMw9v+5ff2zmppOwcPJ/doqbgW
bAGCClVqVMvBbQscqWz4CyQX9IzBQop+Oynf6W80j1hkbqRwEOdaRIRI5oCe5kg0IaUWY2lTfFUE
+jO1gY+jD00k3rEmFqcy0v+V2VTxF6tOU9ERamkLv+fTfgzUEsZkkdB4GZaYkfkTo6cyrHT7Bu1c
KKvefBTX9PaCha4lK9Anmv7cW9VBzDiGx/vM/5DXlelh1Iu8FXCOyH/ZseC6MWSiheU6k9X/a+AA
NcZ9QFwbpifu2TNSWyyKuT9lAIWgrEiwWXolcMJ3MzPgBh0J9hD++aj0Z/2SWyHES4MHFGZNXaeq
Dp4wqfZjiSPH+kxieXgJaECkR43t27IOJd966bLpZXCLO55j2XKD1CbTXVYeaG2ssBtjKWYt9gkJ
lDeG72mpJmG2wsrFvxkQ87DcB4Hvb5Dx1FDmhcEtA5Vcka3TDP3THDh/6Xzo3zfq4uaUmQS2K045
11BpFWfBTo106asPWgskd9WrVekSilZk7tNtxoVR5l+ZHTfT1JSOYmbABLOmpe8iJ/22s6DjUQhR
hLjFcwKbMzLq7BbsjgcK5vfB4/vm6S+UmVjiZFsrQUFkYgZwbP/+eDtb/5XYZ5qhBhmTjiwRXhsM
818p3rHzw/b0XwQrQLJK/G1MYt1MHUfd7dh6QAZxwfQnlX4uqdIpbN+UzgmFQCwfwEcvkH5YPAQ0
LvJ+5oWhQK6C5b07GH/+rFqXpxUOhgivi/11/iank1YLHN5pWARljkwMvObluoNNXo3nWQOZbON2
5uxOOO4ONN/vS+4q6Hak4Q+2rpIowR+u1QSwL3Dm8iyQviNem9a8VzmycbHpL+DeCx0HeumM0GsQ
0iwnECcgVTk3O01N69P2v5npkRTQ3OT1ayqtfZ268RVqMB05Hqy8otSkHpokjBjBUmMb7kRiI0ZA
IRIMKJKevwNBHzdTpsjtHPfutDwHBXfXV+QpHRdm0LvNA/tD0pWuVmUHpULX6vticbZtv1XP+CpX
nh8wEYgzJZtCMSIRyDQSf0UQwkt5lPIYMfudf1rf5/uRWLBsyRhYNSoy685LHY7TLysD9sb3iujo
vKF4tX6VEi9E+5k0MQ2QRkA7zyphEzjf19mrHcMd/ITZ6BJiv5NDif+wEtRWiG+Bx9fYtEwPtvl6
8XWBQITQun0BcMn/g2Kz9aFQVDWhI9FHAKPDG1GmjDLna9lUIQA92hXST9l44d4dZNWIrd7QamOr
dBjtdSgGiteJ7ZBB3/vVQcZ/FITFvhziLnkKAxQR5BaytweskS5uWVjYOGAD/bpAHvW2egb1gOGS
p9AXd1GoQ797Ir+dU2IoHReZ/prdLWCis6bzKFX06mU2SiF17IEgEDr7u0XQbac9t2iovGwlW0sR
D3zkWpgST/rCpETvWxXM2LgoyQr+e1Arwj4H9cIOwbX9j6DK4ZI1bzxxyCxA1rUqHN/SO6ExEz6C
opNpo6L6c+/3MQVQDLOugkQHg4/uFtIIHEBP/5McMqBc1Iq3dHzEXJhRX5Kdfl6+vqgjipZFfBqs
VpL8ZtY/C4zEfcgceNVKK+AUBnL1NcWVbL5Gb5UW90Wqsnkq1Og1Uk1UtsS0j29joKLtQXYQ82QY
8MhX0lMszYrVAzCdT2GVh8h7/ya1PA+TsBtyWVZ/go4vRb0UIrJAE5Qs1BmlHj73QbUdEbZwPex7
fCBv1mcTA4tHcYkimqgfbb/g+EH+wGyNHum7i+fTDVv7gFWkrBQS/YNzn8bKY3NkkkgGOgBWomOI
yi6Tj/+zOr376eDlMOLai0terxf4vGnbNKcQPw7+KZ+dUg+QTre5I+dfwe/zC3sA6JFy2tRv0nv1
MBkuixmJD7oCgwIxv7xxNDpA2KLi5F1yS3XONzBUf/hsuUCvu/whfph1uRBYJocFfJ6kSJ/Jp0oh
rTgJJKASCaz34DdDOBx1Nsv4ZjH4bjhGMKdVFeVfBFdN8Hsi85BarIp60YYPnlW8Drp8gjqrGw8U
mH7YRv3H6rF59vtpCWyR1O6vLUu8SragU1m5KEhk0q10SL+ySUq34FBEU43rPUa53NYEbLtwvNgi
UskU//F57Aw4uTtPTecEimg7MmEd1oQxVYC+DphqYxmWKo8rFuNg/DguPN1oYsP5vNDJMdv19DWS
JR43mverzB0gaM64SdAJaE+VhhjPQ8GRLf/hkgyJ920M6A82lNNT7e5X0y4iexa6H4Zpa26YFbq3
Ve+gAZQYHCZN+dgB4lBRdlCW4dKeNp2YATXDUUexSN3eCQqIu/x2SpU58+RZttfRgUjb0Fjoac8W
XUxcSc546UjfcqbZjWr7H4EpW4TQFXiWRtb5R9Z47eYZnEpWlKgSzXEjfJrvwUSzJoxvgh+sPGmV
fgbskpZo706DzOUTUf2C93R+LQ4KEwnPDSoODEmeydVTZpo6seULycBX0UHTEmtihfec+bShSLdM
pIRJTx+JQML3R80Mx0Qkt5c/No+mHwM4ENlap8ezJek6YHWlURgs+EGD8FEhN2/5y0wCG/Lcn4HK
52IYug0bWYpv8HwVtTGxfZU52VBhaFaPmeQFO9CwwxyhmKOVCNFewNeO7y3AgXOJZtCbkW+CrN9X
mi5K3HCVUC1aJsDmfS5Lb4sCKGLkctdN01rIv/sPWG+gu1YLt1k+Z7F2bXOEW8bpJEOJ9EQB4frT
HStF4wTfdDiHfiIS25qmCT+ifwreb9uqpQ4oqXgmUf7fPp/jg0L5IpMRV5EzbnXPNKd12Qr34S6F
nkzvhYw1I4D/0UBaVAyBapy5dA/CJ+TjmpZSKq/CvgZFZn0MBIf4xnP9ZHlKIE519I7X+kGFRCJ2
Yjso0PucwABF9Zy5F+YJeFLugHgZY4xR3NquRVb7OsUROdcqfevvnBtRHOK19fmMmsUAFOlcu0Ed
oL5LfLYy5S7kWzM1Q2D7KfUPWPpwEZXDdJ/TAecq9VpEGbNNRy5LQvMVBJq2t1ZxDr9x2oqsNqvx
OKL07B0hDAqjNI89AVCqGjR+W+BC3UGHNL4yjpvWD2xVQ+WUumJBO2nvvUHSHmFwqSziuuXL0C43
xCgaVZyto9lGtm3qRAoEpFNiISCP88g2ZrTHUEKxU/vAnfIn4yoGcxdawP8maUqAPqyVWnvwAH3n
DMLkZeHRyheuVN2f46aQufmVO1GtquLztjvV6exMJnCfLAyzIvetPr6kIts81/xgar0HijyOin58
O8CfiFNwk2c8G6kewP7PaXsuO3ZmOiXI9GBReSahwghJE8qI9wAT5m3LqZZat37XQjqndCe5GI8H
d1AKoeToei9wHE46piIf5Zi2N1y7e1YDLqxjyXtLm+k9C/Om5DCt7ZjBGcAORPoCWr0t7JRzWYbR
Sv9lAuwGSbzd0Dy93xCIXQEBAyn30K6ygW/Ts6DVJ8wi4WoRgPThE2jNIQyYR0OmaKXxEAA2Sd9m
51EZn13GAAwlj68suQv2f/KRsIgyq0ZEiCwMi9zv483lCCq12vZMreTuXam/sEWdcdb3EA68Crv3
DJST0ttWmrhOwQc3iq8eKPEnEklevdgS2PEccG2IiaKmeVFzV80T/+Oe5tNEaZ/s0iLeMXSm6b18
5HwF4xgRqYvOoCnYzTdqqVy82125x9jBovRUhfKFBBmkkPlxEEtLdjXP/QyHHHWjy2OurzpqeRRC
/UTGUYAJk4XPVt8G/WCGIrWfPxJ0cauUyiMbSLX3qtUx84BSYTC9fUZ2TjclFyimD8qO4neM3QEh
A5REp+2sWltcRgo3+AVjFtQm5hGkVk9MbNE8kRXujV5LNbBIYnKXerbkNTBIjOEXGKx2C0ePpIde
sfVXqgOBd5jVpIr3kpC/zMyRqH/JwqGkuPVyAWpAA6cl1eXeoT61RPB1wuny2Ta4JXC3Qj930/UT
GGomLWocAsrRv0ZiuqAlX6mXyN2QrBOvuWp9y3yN0ixipIxf/HxUSFFIYnqKipCD+jAKIM86OPiL
evZvhhwTm0sbmNc+eo05MfwajAOuV8RbkXuLFcTeM7MSN+lhWkeVvajAQ4Mr7ATCY/L+F6YCiLaF
1t3xsNj5pp95PhBcGELdq+rWTxT+sglw+Zszzv/I0Rn6x1gA0t1eOXL5aDOGrXwkTB+cK5UERLtt
FTaO2BzhWct+jZU9hXtJTtjQtNdnkWvqFDFazb1m9HyuDQYaOtqdfeO9wm7dreK2uYnpF+uuLMW8
tUSr/kFNgcuBTGefjG+v3wA5Ff+24C8HUk2rEUs0wdnlzQ6L25kE19l/Sm7whsxgUKuLkbB+1Y1U
gdi5/h20E5uTqmvcstko1S+KX9NT7lES9XkA6bMpbcfRCvkrskI81VSrSOxOWnf4dCzV/ba+lANM
/j6MxIr5lc8Nps64pJ6IS/05XICJw2yBJJkjzCQE2OHC3TKxNJj9cMA2+ZoyNy2wc1gKbfHRBY3M
pLFACwdhstzf/dvMzUP4S4slg3IJ9MurkmK7yIu7Sn3/F8RZm1Jts1cw+gbYu1i/lZfIOp3JjkAJ
kqJpeo4NIvkcxy0gf7vi/D/wuDClvfp6Ro7NIZImr1xOD3Ubpj69u9xWJCi3bjUEBRAVSkZ5BTVY
YwilgQf9CZaBDSR3tHSKW0ztI57/DmC2arLg93ykql9LXR32l5EnTe4DZP9Po0QwHddN2nV4hmhF
zBWbTSu/XMTDIBXWCuFF5QAn5UKCn466ADezSp8VEmkJxlpNal38DaDz5ZjSa4UlxEk9XiLI8TSs
n3KKePBKjIf5zSGnrHhp7WPwNsnC7RuELYOreBp5WWt71Fn+9I92JoIvZjpItDXRIgDJH7WGY4H7
ibPOjv9+xiyzhvKe+BNodxOkHbMlXYfZ5a6/c1seJiwh+B7Rsbu9O1QRpGDD+xYoHK0pBp8iZxOI
gzfTm7IhMtMT/OGX4H+bVxpfnmzx0VtQsj5nRwKeBlHx8l0cOGe0Lkxwv26KlrIbwbkW9uBU91Mz
4TQXKWj39sdmi0X6fOzpC8LYgpr1tK6BVoMWbMVSPYu7ku/278ImZVUPWe/9glbuOKB5I+dW7V2B
FAyTVg8K20MKqZcwcWzOhmGmn9YjoASxWXj1GtlpPbs6zjtFpCh+mflTDZsat2s2RiaQ6FgWVk1t
dokCfhz1izTXc3J8p95QkQhIcqaHUrbmmOPMVb0ND9Wlzwg5znI4EqmFiq3R6ox1lFgGjtv2Km9T
292oGJV0ceJxqjaHEFaIZkdG7uzON60FBHJ2VG8ngxl7h2x9KMn0n1gRin0BJVIM6xzlPUd6IGYE
GBpR3bmVu8fxSbl9wSKk2Su7rALU7BNP7NhZkEaMv1UY93V3OoJ0Vr1qQRYTwYogOauUFi5ItPEU
tWNgTKBYmK5nvHYgzLCB/iM2TnsT0rL3iGk6IsHgEmUGlm2Tkgytmizo/GXJjrUshBklwG6CItpl
7+qYtdC9iNAQATxskAEdpUhTLPzZFQCsArZ1A/ybmNiltNt8mAwfsTh43Wmggsj9243+z6WhcBQO
fsnue9a2EHRGoN6vcUnobxRaA2kzYWiPXnUt31oDpmaMHypkfNblGAv3DJcu04E1duJVNxiwEGaV
qafrd2SVMG1NLLqiKddcvWCRNfk5FAtNF+fMRWDUaIcSmbhts9UgJmahS89/df+aiw9gnib3Cpn1
mrw5m48UF1yMwdRjONPGMLKdC7WLpBZhR6kgoR8GlLbJcpaIV7qM0b52dgNvz2vJ8ZyhI2towzfv
OSA2PUUgWUsvzYB/A2xVwX+65Vd9BrNaIAUmUIf/kgkNztVVAhLyme448GOiAueI4TxzfkKyNZVG
VLc7IMqM09F8m5ZtyOKg7BMK+CaZqFGQw/rzlMb5aZpRWKg16JZfDMsHqKrXTMTzYS3P9w3DSD5q
d3KtbisNPvD2VZPOw0hemGtZm4BFZ59Tg+1OxyZX6rRg0VGXRoHw+myWRLhDjrOxwbqxBb0dxOzJ
/z5lU7qb8UiYS/Ojet5BiLTvocju7HEaGMCpRbW77TvQgle+jQxTQ+6/e2gneIHzCcwuZ7+yl5uM
B9jmw09aRlcI2vQZABuctUy63oRvu3RzwW4EIda0nDaWPo5R0KJOGQP/Kl8NzfWdTBCqr0f5L5Up
4ex2gDdsWiY8/toQBBvRV2DrqE3p40RYyQkxRxtD9vWAl1znID7cY0GY722PKQDzdvMVyOQr68Cv
MlOizLC0DsxzcM9ECH1xfMixBqdjZShQFUZOvrH71LRa6XPCIa+sHQbbDpQTepXM1v+21L5yz3U5
40UgnD2dHDmrDzNf2/Shk6KtnY5kroxEYY8BC1mlHKmz4gkrX5dm2mkppF3TaFqc8ItEUo5iCHeZ
tZgpcagZnDJnVqiCsIymgEH3+1x00Ikul7O7XFcLgIXfRgylMS26f3WllleI5KdvP0XXSNDcnAX4
fdfwIGtbvJmcQKuhYPRxIkZG5RaMMO5lo4tN/tInyalGjo8Dnn52YG+Ij7L0ESZIIfRUzWITNtwX
VL6WWrrE0CPkGYgoP4VN0LkMqB0Q80e5NeY58MvP/rN9fyPqIiPil28dp6KIFjScqMyq9KBq7kiY
Eh4xrA5o9L7hkAfoH4unoLwzskRUxXYnBtA/uomxzw5yRF9cD8Tcqj3jZvTs8M8ORf6XTozRkLXs
EOF31dtjid2yskN8J7IlP+ZAfQsbm0WlxeUqcAN9u3Nl/eeNQRkOK3z8i3VodVsXI0zkuvrMgFdo
+T96e5TJX9cg2WctS9a4sMlRxc8Y+AuKlgyBHAMD8Wgu+RXRmikHua/ewsVBW96yXYajNZVU1Gn7
ENwzg/8U/7W5cUiibu98aB0F4WDdklQEEAKFLGwvNvHTWX+c8HLNejQJ93wKIPVIef63amyLOzJo
QP0ozfdJQKnL64+78qpe5xq/agkYZpbvFwZim5Es8p98hAmW3aeWt7vdfVtMCZZ2LJqNNkoB2ILX
zsYwvYKz5D4NBYTyUmxeyt1IrKObCGKLjadtyEu7XsYZQkgJbFaih+kOqDKcbdeV/vNAPl7iBsmB
tHj+kmiiMNh1KFOCFxvf2zBIin/7R4wf53DAVnnZzDURPylCXR2d8dd1AEFI8oF1pB79uBeynrbj
BeQ6vHMi5YO+lzc/eyzQ8c+3/O7+2ctIRTxfI7po9yMtr7L8te8KfvBh0hFpdZm60rPwCjmoe30r
QLQi5RgNhaSNrm0TU/R20slqcP3H/uy6iJxDkzDFG278sEZcM2ecNF5oB9wWKyyL3Mks/2NfohRy
hKItGHHdBGsbXXbfjJIqpadNui6XoTLQLDoIh42HiluZ8ktHeO2MVLFrk4bhruU1ZYXjj1eYgFZN
R1scEMglWdS109/lW94vqrBAGKl7EmsiWpw5qM1iMWsdXN1QmfQ8YkHR0r06DZ6qeBdg8cDpGC6C
wuyBKA/anMrvFPaGyDh28wBU9k+UBlqqo+qy808zdVdqL960+xGgeMQ8onBxvetWVJA1qQdxcLrC
vYuDgQSCKnzf7WXTopH/oS8oT1rLGE7tf995RQc+uITHM522CLD7Kt/I9ewdbYj8NZ6e15Y4p9GH
NXa6TCKTZqEW4IHf4dzsLa/bu9JkuZv6nbWFeO2bksBeFm7/scz8j5nSrX016wl+8cAOE8f+fZxV
czmcsGYiH9zrvtsppivxVlBrEwTJjRmaPCt5xY3L5KQvAGgBr+B4SM1+cDjbrIAADQuSDXDq/L0d
jC6b8ublbxZAmj5CGgdrw0csmHgBBz+Q0ymwMJFwScGSnijzy1eUWzL0VfeBCapqS8cphx18ktRD
cvTPIY4SsJX1RVGSUgKTX0QUl7Wr7qU5QqZste7h9OzIUD2Iw5tVFg54ETKXFJuEdtJ1wl8XuRQb
FAp6zagdJHQBfQvmK62aj6/1+b66JJ7PTEnA6a7+xbaUNu1DH1LQBpOjtvve8IbaTn3XSFixyfFg
u+FgoWq1s8YOuQOgfdQSUkGPab98DTTmLrB/g23WH/CuW5tt5QAjxzFIpnK6/ZB4tZG7hOuqBIBc
w9JQ9xYy5LBbq61bn4vSzsB6v/UXsIVC0ukurwTnYkHqVT7CQoUhv7RkWwg370phvHepa2e8wxBC
h5NbIW9KpqMNw24nogHLghWRUxECUTIZIqttOLWi294L4gTsll2JZdr/xqwWEPY82nfbTJA0efLi
shKKwK9FtJbUd1iGt8TWfHlvZtaGCflC/3b4ZEd6wUMjcQeLq5Z6pSXMdvVRWvKeHGvt7rKBW0ks
1TEmnkzkST1NSsvSZuEtoCSPIMY2WYrNs9jhOKe1l2L1qTHheJHvgn591GWrXsey1bPPBhuOs8WF
7ZA2+SHMp9pGtxPH4b3nj2dxAZSsDoZ+Lus7tWhr2pLGD7Ja2yUO31HHRkf/oy7x1fSOCDwzE/gI
J/sMhC/SccPN8BqXgMx2WoJtCjfIEyvnWIHalredvS1PKRDaZRJy3pKEtkx8iKlW0v8uY5K023G8
zhjXVr/o/NAMiPEg9xttk6hkeavxy6fEe879ERVcxEe7V4N8Lh8d6OEiOeS0lbkuOGi/KXkWr91H
lsZgR0ICGQdmPg9X6XoQM4KzcVoc3VWtyr/hpG5Cm/215jdLSGlocaW665DAYms9K4GNtGlTgoYX
G9cWY5qix3/+Tdt/fOqj1eZcI9w618BufWu6tJSfDas993C95x9OLcnJfARYFejtnI0cZNxZT9Ov
YCJNc/z88/BKWzCRv3gIgQ2tG0R5F0N6QreDEof9Amo0yG1EwOqEJoovtBXRJwdyjTqYi6tx+zqi
KPhIoQEpthYcy1YRLN0yKuT9OeMUlRxA0UdaJ3L+fNXOZ8s+r19PAe+Mr6WrK3w/2EnwGssypkXP
96OKy/inPbA1CVIHYo5LJr5YrZT0SQQZ2wcUPfA8MuH6ABc0aIjC6Ez3ckk1ImSt5eZ0avmZ5uQO
Y76VytAYfuEAQ3CCTb4hIYS2TDkC+MORqL/EQRwhrLXNq4ccZ7OgBxYfurtL7D5Zeyu5BYRihRWg
mk22q+kJyWuKt9BfUF5QOAnwd6uhKxa9J0DmJoMaAr4/23RHv7ybkBdHzVaXZqjJN8tl+xfSKdbm
+2RQeIg7Luc9TjrdhhXz5Cai5+wjbZwRf/7KancsnbrQOKf4gX3+2TAChZZGkk/LhsyRichtF1W0
KTwjyl9qithQPY/XtRjd7nB4bh/7Ij/7+2jHwUuiW2KdHnyCOAKRwaaeueJEJW0/UvIqqB3ITV+1
vlzsbX6CcVdv72wjUi/91Nnu1/GRkzpmPiV5iaxf0+oSduhEI/MDuOLmNBtgmOz7zDXpmeWQiI+n
Ewk2oHEdur2LgmekgZp0N7g68qRoeAKmRG0cYOy2lwUtK08HNNlFrdQM28lusB9FTRcC3uMRLu0Z
MjYfO+Xgy/RMAch2NxPWad/cSk4Wl82qHzWW7f90d5DUQRriw4xluqf/HNhbl67vcywLyZNEaRCo
jKtEgyby/aNpXbzOb4A3aMqC9SJiZBnuvdBgz53JTexpl7yNJ9v4DHceUQmUjM8EnD/2o7Ql+bMa
jtpngxQyrXJYtHHTceheexUTw1fqvvwdx6d8yH86lrC3qVFjInwx1idKeni9zplK3Kg/hVOdGvGD
znU9ND5umFVfzHJRiwIFhRJa599kypOqI5SmxDPFDL4L0XyvsdZ4cbxTOsqn5PzCmP9P0Fx8zS/7
XPkjNIz2VWUQN0yJ+3c+T6GL/zl2itAjkOFzO6WYTbm2/13tCVvvCSNXAPNQV6Is2PA6P0jcSp2t
qIOlFYPcz4xhxOzBKlRygFNEARPyeQqZg2bnfiUepKIhVnnazjMmtp2mk6lKfqAiCW+WgYgvFC27
CBZp0f3QWut70clcn9P2owf412XswlGuNpNcWNyVytPeActSoHAQJ4s/Gr3CxmNmH2lFkSibr5EP
kWL3Ci8X8R7qu+9Ta3tVD17UVFnmqpYibIugCJjR2SgZIAvNWxfeg6BFhzOsbAh3giy5aHzu+dIT
V0G1N9+Q3FqFqBzuVxIw42y0lPJxKS23L+vZnDMa0bWg68LanWilcpHSQ6AZhT6hAbii7tzuzGpR
p9045admwTmnnXk9fNwSHTScJfNyVw/UTc2VOwO3V5OVJ9JmnPDRvhKe+o/cXls1QbS/GuEXi0j6
0eW3ykVwGVFCxRUWnio/mTbESyUndDTnWerzSR28VjGn9yPFqfOHlaqAAFSjeWkVg2AuHtlHBtGq
zoLO6QLOo3QY8ZOuScGywH2r1zMoOWxFfUk6W8g3SITHBrF6VNlVr1xFckJDiqi4XtE1HeE77Gw4
PzvEZLYzcotFky7Tp6BLlTUlOGNiQwhT8QjFzfBO/7wirTCkllun05oMC82ccpPrly76eqwVjU1q
xQCMQIyxzNXJUFgj9GuzmHICOswRkYlJRWxSOr6+AfqUynm+BURNMRr4KPH/DqebpOkXZnlrqiKZ
Y4Twev4yoxqiBkkJ0+QDoO/APrwJZHRupiY+IBhlmMlYUXiE7/MGBfbniJGGTl9xhWzA540vBQrn
P63+MObYPAwILwDKWLQmuUKVacchCeg6usdbbhDGB6X8oc/iGI8TTHSEvpXk1z2i6+fVW1ks3U46
t0tW8fl3Ur3vDtSvymxcgUY011YxYuH+Tms3U6aq0xC2RLxlxiYjQxlU0TMD/N/co8FTjRi0aGHI
gIao+KJrMmzvWRhCLis9VK27gVzgsnzxv1qrh92pDVY9f1WCmpeLLzVdNIcl09rnvupptFgwxlhO
UGY00Uqz3KI3g+BzcamKTZtAlwiRVBof+dfhK5vzKDCDXvMjE71G0oZ9IDMdXrj2qB1VngWAzW8b
uBK2jJvtxHZg77fPkZ2uf5jQzfnNlVW9XDypH1Vhq9Icc/D86X+Fhopu4uKJJPS2ViCI/MpTxNLO
/aAOh/HDBFRSJPG44h24xgSMVlJ0ZfFk9kUMFlQ0ADYcvSTyA9pkUmBeVWf6CfDZemxmcxfHX15m
dyknbamk0fHzHo2UqhewqFVBeGRmfRhDQkH/iUUPWmPZDhktJ84Mzy9JAUWWvEhfgC5enP4NaG54
cx9cj+lIT75cXl5oTG/1PIkryr5TZqIkLA9WQyxPEqYfwKkJJx8sHz1qP9Yx2Nkw2x0ED0EM5WPT
TwKKsEmx8PvEyL7tfCOFRr6OmbQXlVRUyh19emOSyee5u3NG7LD0noN3k/xLuDa4jlfEhB1nMk4b
ok3Zo36GGFaigk361OeGiw4nTInAbjJeFYCRooBQNbR2SjTPUuyWLxChsOOJ9a6DUB8yDYdY+hqL
mMIx7aipt407wr8QfIAdywizmBLIUxIX2nm49DH2P3tjXljr5mrD6V+ollhljDtVGtDsZaArjGUg
VuvZ0+amo+GLTrZoL1xGdQ3fAGxj+Vn1XxOnK0N5l0qMARExPbVm3sTF9C9Q1TGxNyW+mC/FLoL+
pwJk47xSofM5mi0IbaVD+Apoyrji4CZz8tGKJZrjQPltQvNGPWypzukgrWm/SY8JNGTlSPtp/+U5
4YI7sQKjY1KoxWTPzQ6NFiygVsjKGA6oSKH2IV7QKKfYLU8zNslsWgwH6lR/MuPFk+ObDapbF1Dj
Iebl/8Q2IZsPnnaTKS6/NlL4AOD8Ah1YaOzUZpsjdkcmwzQCuU2MDCe9E3PVq57LWzXCTcSnA3EK
E797RUXozT53jVZwpscpOJS4y+kktB3l5dvHCuz09K7/7T3CAK/BdEh8NsFuMmqkBajvoSczRToD
oXb42ay8euGNfn7QaX8PHbvteAXvFy9OmWqyXs+cQ2KSALdJA41l8yfNwCw/hQJxasiNaJEOOTFj
u2M52JYYnv8kGXvWvQvMOXCiX9/yvGSqvGuimbDeKD0eymap0idQ8jKWOm5FZHeqrdg6DbSg6gur
V9YovSjGqBB4tQkq7ICkDeSPKdL/J34mI9FGqTI1T8v8F6lmjFzXLNv8hbRoRSbBI67O6RixFt02
PipnAZgobTIExJrTwFLJnQ3pNOQaZThi6Orjlbbew8dYfKfjBLRYTmhlMw779u/0DWmPCizJwd+v
b7VH960gyTY59wXmI/4yDTTtP3nVM2Uh+W+a04+zn3D29PeP9obTFDG9bse0hyXOXzdWz+V6ZVhc
gQiLe/8ja3nSxr/vH4xNzVv+AtvAQhAw9CXRzpxzLCV7DNLouejB2TB/bDDD/0v4Xp1hLABsVTte
/bsQ4Qvcsr6jbMMO1BDJntDnxksTFJEQr3q7pW/3Q4SR0OtYKC8mk5aUCaynADmdoOyq08I5Ld8O
Fhp13yue6kD/EP2zYqGqnMwIMHbCc1c+X/7JKgLd2mU661ggRH18z9L8M3q7ogd3TCZi+9qiViu+
I7b0cr5y/q3RvAYPnYxPCiuPBQZpZ6hoxLgUmeDeUF3y5H2r/rnCp6ywpxgAcHC7PfxKwtSWEZOt
3ZoKCv3o72MeIFqOLAdmY8plTOVXU/e6svzI+0gQFCY18+t8+9w6QWx+JInJrBuDSfX8IYQgy9cg
OwdYp9PjrCZ7wDU8wwMoBhMLRdb+ejozd58UXUkcrb6/N5kRhyhZB3/NMyUrwqQuQze5cyCXWaiZ
Zmc/Da6yu+WF1Uu8PQJ1QptvCtm3SE2ZEH5ruv26kdNt+5soPByfiek6iEpp8FTTlSbtel3sHiaI
4/tLOX5iXCiZVqVqZxrT2qc1HBVmlScFh03PoBKJNYj6DiD9NSeHabqLr+WGZ2wNzTIB0ZtIchEU
CDIve/5xO1UOjyQWRgTn4Wby4JtxK/V46WfaT/Td3WFRVJv57wKwzDyYRrzesTfLjeuRv9TDj+2b
hur55SOAuCVUg2W5rQes4Zb8Hm8C/nQT5xjzHcuLTVeNsqJUcGuzxkTO3Fk4Ztwpxhd6QC3KrfK6
UM3fMefRlu8LBue7I7MXv6Nm8DHlU/ILi1+JjG+hFVba69f6J4Jr3RvuA/Xt9daxAaFWGjhpnf1I
kIUKJyAwr7rbtP2znp9hnhx2sgPo5t1zBkQ8IkanJc7N8p/pgdXZ1URexE2liLi1H4M+aXi/sCmP
Pw0VwFSkgj1lK1pPD7gEJEYPMsUkMVKkvxf3jsAFfrCXy4Jz8dJ8msgSBtzLpkbvhN1foQA81pwa
4mXz1Kjue/GeXbOCom5/gp1OEcY6bm2Z98HrM9zOEjKv25HS4OnK9M9/ST5XATwYg6TdHiUxanjB
wbUYSdyx+0SWD6wZFir/L1Ican6z/C1PMzABjc02o8zoD2C7xnZFcm/+t5pTb2rddHDNjLmI7tbH
v61kPXHRAGWm+FC97LdT/GBYqH9KDpjWyDObms63+t8XH9ygMlne6/UDcO4Ju8Une86N1s/53SSO
KWfj/pq5a+4JQpGi3kVTdg6MAvZsGHAa+pgcVqvOLkSqcBFp0ORF8zaty0rB7wAbljwycJxzd0Dw
Rd5QnglahrdXM6jJcS/imhhNRaKVP9MZqhaT524PKuMRkf9tSFoFD5n8+5Vq0iR4Ni0Lu/Vu9Lh9
NIM1eTObt0cHJOp3lLZHDXObP19C38wA6euJPdlj7MxUi638TActW5hUnAIRXPV1sg+WGGp4JsTM
dSV7uriHX7F5RkZ6l+/TgUO2hEr7Wi3FoKlEHz/bpMageTSgfMoshEVOZL/1LcyiNzag2GaEhom/
MS8III8Lbn98cVTiF+zoBJEomSW6qsRtObZ5xMZ2ZNspQ3RAvEaHV6wSdDh9yFqPfahDrn9FmTsZ
neIJ0NBOTob2tOrrOkDprWBReRwmAKFanGIoURIHnC/XswWZijVHT0uIPWddqeqoGXnS5Axboi2k
rtlo7eCdOGSPc3l9KrXh74xM+Y66wvYHJKcobfyffgQxi+r2C/L7dN88JvgXsunTCsW7O0UiJpYB
TkhKb2CPjYuHd9IoskEJU29Tp5Mvs3FD2yzP8JJxmKlD
`protect end_protected

